`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gNjYnuOA9kZ21ZKcKTmdgQx4PVvmLELIL/YInu1OKEATNUsp/+IjpvWZFh22yKXkcOtVS/1PbRvYB7DgUHlGLA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k3DKY2eAqzZhMKixr1blbXCTPXga0x5Me4uD4wee8gZuLdFe0XC932kSUxw3I/oBuTvxJn53iSg/ro78gqdvqEUQAl+5FOvdw1vTpQZxi/bTl+EjkeOJgeqtrFC8ZcJKpOZeaWicTM1co1iIvOJpLYZNqtySNDB3g+8aJ1WwtkU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wCvTJaU+d0n4bw1OSavwvUdrsA/3/A/lI+IyZtPW5eHV+AOFh9eKGoAZLo1bWVg4UdXqCUQ11gqGrBPv92PuvdgMZoWMkEWZypkP8owkDOvkH5d3cdB6QqgFciRG4viH92OXcVj0GoddsXKCA6SV5224jqLXsv+LVcchUdKLsZtbYiS8AjEwY7d8Urs3irR73jqFtQkzD3aykX9C/3PPYblJuwDCM6QBxmB6ur1h/sm89c1XcBOx/WSLQha0vdA4VHA9Nazpv2R2kxUc0BFHPR+/fbYzvE+XuDHO7GkxgYj4EI71Zz4PCstVUIa3u+9Ih56HBjegK+5zCcz+9CsXsg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IAGIMnlYoyObDS8RZP/iGYnA5rCr6ttluXjZY8yQMKAhPF4aYobUzncSeyuD1p2nLZnGMEmI2PzZRvMSt6CVJZ8dYnopOQzfAmzD702VMN/jMBKgrUFuwmoLUljSAzc1kiQCxwTl2AomyPLHIhq3k6s3kfOz1JJZwveAcFcNXpk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nu4BVb/QJbnRHgvN+tq6ACSuunlb0sw2eFtZZBcwJKmwIPCWJfI/LCs0B1alLpchBVanqgo7j1jC20L0lsybuS4HSPyCg6/Fr5ey0oVUWgBnFktiU4Ej0GxErncjM77/qEaWPVuFemru0groN61Y99m/Xbn9DeB6yqZZSv3BT5sqp0P/3gEX9uDOzvyzGB7iWdgjbwExT5bKX8CIPgpYJVJ8kD6+ROYBfClSXekdstnw0iyMHxLjEJJHMAYVbNplwMgyOeXG5htDTO+QSVOqAiL0TCTUolt0hdLz3C/9g7PW4cx+1vTqL3KL+H9lZh9IHyaswNgWvBqeUMHdPRhd8w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 33031)
`protect data_block
CVF7HmyTF6Cr2diDeHuj1EYKKCXQ2epfRmkPrJubo1J+QY2azmCqVoapb60OY0uSOQF3/J2z//Y3
YeYd2RNda7lUFbuRdjWoD8BcONyhZTdjzZMd6Nbd+fXdKND6RwwpzFJo19hUDyP5j8iUu8MB2Qy5
K/V7e1VuC356+naEX1E1ynE5WiAJ1W40HKKZcuQedWUMydfCJH7QtrKeVrOdFUURSrtSY0Igk6EA
ZZSrT3HhmlWMp7eBnyScYqk6qaTnFjquLmHKqln3DTsvVfPUO4Rvz+Gp6sEOvVazy+G0jWjoVgnO
CmE2B/qvSZKss0C7xxwd5uWj/VuTY/Ma1CYy8K9ejDtg1Sntb87tQBx3BC12U1CyAnn5lbuSkwqc
cS8dCvWam0yroLp0ujgW+wE6I7qa1bd11fzPu/cgF8itH4ySmh6FuFNuGmjAyTo0w+HhodnJ2y2S
Huuleg7nIp3MRuS5UFKPqQXcyS4GxE5F1bWHyGyZLqwmyK8ZpJ80+wKCgAqp/KE+O4mYegHE0bw1
n/rJ1rpXK3swrBEsflu5r33xrc1ab6CA+eWxas5lsuykh3VJj+j5JJ2rMhY1/aJuEoDriUPJdSiT
K5Wtt1Q5VYfWlKJw2v/QCcdLkHdvWhyarBpToEkUcYdamTM0aUVsiqVddyR4sPPHlb6mAJvdIYej
jwGeljGL3BkBqCV+VVjJKSH4cxSLY4r0qVGz0BJAcIAK1GmtJyk7mADVousAbr69T9kPQbzTTQvG
05F9015v+tQa7YiE1FJg/jd8mJoMYksYTFJ9UdpiIYZSvN8IksYeJsj4zHwWnVTdtlo/DDTi7QbZ
v7p/+V6eCgj90zsyV1bPu3S/iEoXIKWHYFoqppYib6nrQrM1qt72vluLZQxboVL/k8hQ5AoDrKKO
hnT+ziF/x1b0GIgh27mFT+3gjnmsu2z82GMI0IiY9mZ3Fsm8t/fwwp7CCIbgFm+kReU0hwwRNjD/
Tvk7vt/PXwttJ9XF83DmdWTDeNUDLU/NhYZW4RznnZiBsSAMZXL/TX2wU2Frj6ncMpFp2MzullEe
OrNIiq8znirYSTUhLA17JCo+7rFEnd7z9sTHjKA3kaynxUumqvUqLiuclJPt8Ton4I1iqbHw7pEj
dMtos3oXNXH0WXhl/WmdFBBwtuHt/t0LDAsp+s6ARpMHDqaoYrWb0xbrH5XNnAAxzoNPKQyF4kT/
0cFTt9gjpQNHz0tVDhUiQy6e66spYcFHi/BMuSE6p2UHa9L5TopZISHpnZRsF6sn7ARVIfp0ZUTi
pdM4kzEh3RkoLBixwOXSUVBKc5MDncYJCwG5h4dEX3/L7o3KuQ5QYdjGLKluFIU5VXg5TDnNrHgT
3utU7zCgmxK6box52aOkkuBli9jVsJCt1kKDkFf85Xn1IISTiTW5UyoBzoy2Nj6OL3VO5UPUo3sm
fCAN8rJmeKDjjsMs6F8QP5bMzpNF+HghK6MFKZiM7we//Zqch8ag/b3IxApqH6o1U1x9jcFD4CoG
D1YXXnbcnRdL9et8zvo68eNBfbl83h5M817RAgVmgfXdHwOYgQzH2AoTwwSpjicsNWBMiuluuPzJ
qST1Oegk7/tf1FBcdFmMTwzFJKBwsERHyCuFbmbQu8KlsFvYLQMa10YSiUKddsa1es87orTdKrNt
5SiYnrjp6W54e7NhJ58H5+ddRskPu0PWwuYJoAkWZAI0ep+L68tTtZddPZpSpKR/8S/LpbuKkQBn
bcWWwtifAh27sc6I1GA65UAvoD6X1jWNM+9ehevISLGPbdEfxXCziVSy5cUlFI/NKLhNluDJ7dNd
Bx9ae/1yDu3DMQrcfZ1xGleqZXe/8jq4m47tUR3ODhp6L8jgC1bmUDewjDPxbe9tK2sXeCXiI5j5
RYgKQ+44U/bCkiT9roavrGkmeK0wVkrOh7tpo2I0Sm9SrJ5a6Xh5SW6vvONFsRtpIu7D05wrIoxU
7GeSFyexiffk4ZmlifmPXspWFxxLiwEVvFzwqN56mdPpolgGTVYylDuW43WqsJOZJ/wTd9y+XTsZ
B2jM7gOdP9Oy4nzpih5PGS7MFzhiKg+R8QSjlkYLJnpmPt8/KWNfYYVYNQaDDRpJIqANdjEBixHA
Fh1FiPE30+3rSJLYfIOOOA/Uu0D00lDSUyea0jSR3JNhGUySsdXdOY4L3VonCVsBf59u87aNZqb7
SIrUhS03ZXywq4Zes88dHNUWGWZ7ZL3k93fD60sc2xhvM+eTqI4o+bWy0w4VZEbKd81jPYkAdvRL
nH2aeNmRVX+ghE3pk9+II1bN0jWM0XfiyuA6Q7PrB+4XmQwJZrNHOFoiyejnpp1V/xoSvWzjLPmr
ZYQMuFmbOlP+aYDW+gmnUJSqddwDEgxFcomMncB8dJzgA+HwevsW/lieqFSss3KlHOA1I5idOlw7
kjmVmeZSoBqrcb0Aj4hQMwvHYojPSRHyh8dr/GUqvTyQ/XP6OBeBZcFYtyG92qRhfn5xX71L/ht1
EogaMvRqf2qcIcWZXbSIJbiENuVy/nyEgCSTiLjRXlmXMdRtaEnsoIFU2a2PqvfCOcYBJTWrkw7e
ccAlbpVmGHL7A/0nr0HI5n6XHGDPzZ8hPKuyymWqfmSY5vlSdVDBQQsONGG9E1VOt04OqaafmxW7
MTOzVgwHnOszrJ3TQcVnmpN2WmB/xkPVCjkRx+5ox7ehgj1Ny2aFXCl9LgH71D6fBWRrcNndAE7S
harccYFGQv+xUW6zvUy3acf97WCU8J6R5hWqKY6g5yle8DN11drrISN7kROzhF35kW4OKnikw9ui
RaqN3mySzgLdYke2e5eqFdTkOB0xiPorU/2K7BlrLt7QSi7uzjUvi2ZN3Sl++FelxG0sZgnlo8zr
iM47NVmtakb/sjNVzx8vcJEY+ayMnW1UQErAurr5AQVQ3oK3Kdwye87oXrxI3/uLRCgIerFIgJvV
dxPkjekZc7BWdRJiYCOlb/Cww6Lboqu/JDbLpWDT8fhVhm7WQ+560pep2rHLqtYN0/saLNlvDA2E
bLZH0eo2xHYcNUxfWeF+L+wOrGmJVFRlpIRZaviIlcdyOO4KMZBKc47INSYtQL1bOIXt+RHccKTp
AboC9C7sDTJC61ThrXshw8Z/09Jmj8qPluRruBTuE7JzZMgDxXZv7Xr/gWdTs/Xa7jtWuvSZryqr
guMPqjncHaDC7S4CedxMwUHD0wtkxEGOl6K7Hv7jvM1ZMllsbSwq8SNBI1qU2LAMVsDqvGYXya5p
SHNbsvncpAg2/FLA1yr937WscUl2l8iv19+DCfkFs/481mKuLNU5rfUxLisserA4FJlsIT4k/ju2
hSFxlCvINaIePfqFl0IIFQnl/DtGr5a0bzYOGuMWE4tIwDL2uxOU2X9Tlhyd/W/7fNAmL1iVcY3U
qGXRwvIBQzd4oGIF6dZniBK0/PuxisuMmbyjLd4wP+1aC7lNLvHoHPlk1OyvpIFlhwOWgdEK7XmP
6NZ4slG4nTWaYSC9fCAfObKtPeNynCYz3xRi3GEQ/fZqY/5rGYIXKhfMZHW++I/5SRXdUTuKWxLg
9/5MdaeXPNCQdzP4Zwl21O/pWccAm747ZUeZlK41PIphluPT5oFuJqsyfuyCjmcWkL/Yof2wB+7U
ybFORdXURgr6k7zsDB2a25o9WPPtk35Fs7TvJJFvFlSYsKJiKyryyU7XaSKHwMQ8Etk3Fp7vN2Xc
l+sZ1no4StRc3yrViNTjg9IJsi7MZ5P094hQQaTV66Igc/ATRIcBkWa9Mes7YRrFzu9pNP1mk22V
V4HkBGYvI8Gfo0Km470AaGpD7BxtryVgKyu7JYjX0YxnePDnk/WFRpGgzgRpRTXCUZtoxGHftpbm
HSi50fylhkT9nKYRSRaMUjhgdoivNy9zeHX4b415mEKaL3gm+tdxfn/F9vCa+rNxCUR4jALv2jA5
IKp+sHNGF04k7rC5Welv+C5Gs3RkrWRQpshWUoA7GFoIhW5L/ZWSs8Ik+UqFaosajL5XRM4J2y15
gZVeaEeJYSoLV6rwP0Y/TEJFLLMEWeb8zfm/Xo40GiBwKjaqkS6B3QzpJ2yDkerGbCLgitnxmqkQ
le/w3ydE5wyQbXt5sX0eA6NV0p60DBMaj9A6kgeMUy+9UbIIiGz73OKJZCg+5bflXEMHMDcHcUmB
vVCppwy+8Vy4MOotD3fuOAF8CeRn/kIxB2KGr5Q8aWAJUhAh1COuXgvkHGUbEYoCrJHLNS7Cl/Hb
TuNSjI7eicKFgkw50h2WWOxhGQoV2UAKTlWtrT/rMzKUH1KbQjirDBYqcVpJwewhjLwToWtqk4Vn
SF6yAnw3yIu1h59ax9sP6Lwax96XoWF1/1t8WMVSZ9YiunG/eIaKiGnUq1N7Nc4DsagMV/Rdny7j
UXlLOmQX5JSAbs/cytfelOLIHwwYH6zLePS1xzBxQQig50QbgI1MTsFL2QwctdhuV6fkL8lLFire
eudtkind8y36/pdMA8HN0XQOTNLsfsMK2eg8Xnt4rwNZw4zUvTR48S2dKQKMz7d8db0ZqmpgRkS2
b1yxZOgdcNBBQzjQamTwX62QBqj9UZTRz4lZheQW+LJbmFVMTWw9hdVnvQCqfyXkCGccr591r4EH
hhMT3afuc01ZeYSVhEkzfViMa/YLZcl2l9oY59AzWv7TbiS9py/1hQuBNkf61rEpixJNXyON9y0A
Fwc8gDPbrEWaEPQ5D2HRC4k0XEnKUamQQvsA3wFapmCHzXiaROWGC7EMhbgAYfwUyg0SK9tpe4Ob
dV2T+zXYbQodceXFUVClKOU+wZS8G1Sk+8w1saem+7VrCr33ixmhspE/ehenDAZJ/7nT/JHEsm1f
keBHN2PUNanX+x2gxmWtoxBH8o63pmc0zGCtBIJIMchGsVvJWH2eog8VsSksX33jy4POJwPPVtg5
q5cECU0BKkXEqv6KZyh0/4MSSNmrKg/fH5FcJuFm4p7vCBPy/o0l30GmyflcRw9zMsGYnjPumJe3
5UuHSR7bmJCAV3fkBSAgB2uIOFYu9W6rqh7oS7kUq419eiQTPak99QFyctnyEOATVMw/14wcUnqX
DNo2a9ifruE60V7RMV9kBylauLWYujzxWxpaQPbiRpABio3zcI1JCQ8fq/gwByBDjSnoMg2fmCRL
tnaDjJQSEGxV2H5wnD7/dw4y9O40/B8x0t5GWQEmApYQI0Thor4KkzLAb+bIenEAgNBCSPUHVSXZ
Bgxg7+m0MwMO1O6nzOEx2Ad0vL4pK+kSoXbWkjTAPSXTLbd8HNSyozzwF/ldYr4w/cUCoaxjyohY
Vug9Y03fyAYL7dAdoOpDnbX42eBrrYyFrkajGbwF7kqw13vdCoLkjribZJra8IOqMUSYjdhsTJIa
yG29joQR68eyvNNcCnX4uy7n08lqz56dJr+3wbZ6viKw9+QbTOSIhyiAbzdiXW6E3uKNlGa54qCv
iPKK30Gumt6EuQXyhdQKr4e/DnwUmT7/eJ5qMoB0zkXG3BpCjWoGC7wwDAhy2S4R5JqPrVlcx7ff
ProryS40sEA0MOFaiIg4aB1+2CAYNjFlfFB1FOSGu8ahKw0bTB5CusGsiy+5CZX9VOKOsa8HAUxB
IqYcA1fGP3kr6PSVYw3zq/ltLdgj5QbWJepZYOULRcIgx7dxPqL1u7yQGkDwVPk47t/bpwg0JLBV
tw5w/vDIGK2xOanEfGcG82KgVm5xOTA29UxzmB7sB5Hm9W1GY+SO6FtGrYsFUEiUm31V5qKNNt7A
FfL7Fg75WAm5IPReZhN6kZPRnL05TtpSoCnip/wUQ/+ir+6nRxWMe7h7870vbTHdAHFvOHzQ78PS
vD0sLtsnFbU8G7PKwip8XpCJPfERU/UoXu1uGfw0vV8RnVE5Lqyro9MOY4zWObv+TcsjgXDgYqZY
qydp7W6CMcoGSvFP01tCs1cohhpFX0t3+EJWziAPSdPqExbYfxXOuStdXb205YTRYEUCb5a9gkib
7jRRqC99PMLaeSPCVYkm0eUd1TcdkIljPDAzSyhERDwk/NgOjTavu2Yk57tq/g1dift0iMPWk1Oq
XLxrrr5lF7FAGRM7FKV1BeGOJPuIJBHAIS671l3McpOkDycVDEs5WTqSFtQq86FGFSLTYlHEcDCW
wskPH8HYJELe/zKw+dqacdnYhHdxAc586qEoeyazKQeF+dJD819Kgwm1mPSgwfz0rsfvXZT4jnS3
BJT815GyBxSj09SOrNj68F57lXgr2bKyW1UyIZGXW1/ZMPJnF3PSJ0qweRN49nYCMy7QKCwoTN13
EoLBTrk0ozUiHY9xQt5Ss13Mr4F32S+Vt4UGLnErZOzLuOpXF+CmcaSDNNDFGL+EqH6Bue1/S7rD
fzcVktVv2p1NqZ4ORPV9if6wZls9FpB1ZPqhvap5gMtHDIFyQ6e4b3Z1EYXiHddnRHrOyfv829vT
5rkqPaov20Iph/U7kbKC34iWluTDIIdgFRWXPyj+NB2CN8Epvh/j5rmtetnwiLABqGAa0sB9434z
HZzN2Z7+qN/yG3dl7d/7xnBX0+yUdhXeiTBcsjNwu8wkB9a1RCpjaoSyborYcPcOq/SCPlR5gJaK
9WKSiNfRj8pICHRJrSXqanRCFMo6bK8Zs6H5fhIV7X+qSEi7pMjQ/rjLSNqtTEUR0tBat5zPUy9I
avNsPGbn6Nvtp5FajC2CAThEaf+ovexM90tK0mRg7+KA+06N7iwnsrU+8b5tLZe8jHnOpMDevu1A
MHjB45HgD+MWs2oXPJX/kVhLAu+mhelr6B6sHldUXHP1DwblNerlyh5R841rbK8cEorUf48tFXcr
SPTFlYgsOcrgtBAfgsJErTZV8tIjfK5Ick+P7nqv1RCjwC7kVXHqSyfro3vLtuoCyOFBdFbkb0Wu
i3sbNDEQLv0fU4xe1D3Q0Zu9lfaB6xcd2LHbL2di6T79M02A/GDHhf70OrhVR6WJ8k/8LNnms03Z
J4ahLFEVamrwiF+w5tuxxCQOu/9sZjwdHDF7WkcYTcNyTkiOcmx1K9PfRCGLZ343jJ0FEfroST+M
eldMYiS5Cw0xiRRLtYvDEWJfNAw67x/O0fa5Pz4fhQal9iKIKh+YOlTUXZxYvjpc1R5U6IwMKbX6
cLqj1EVDgldAQhcxqaL0cl94115JDHk8W4F76F2qswaoq4CYL0OBzfOoYyo1Pl9u9UdOfCz7mybD
KRZ+tfyI8NI4JA4OMwu9/9uaS6Eno4RzdGvNbtz8Y309h5lclRVtBUvj3NGdS99ETXPnS4dUP657
bo/g8IVZur9ah24SzcV+a7YMlQ7280GU8uQVNI4oNmPTeSbWvQFLttaPRg1oyyhCkoezn2n15moC
v1TUrBGJ5vc0kNPpi1zJ+47uGUqk6KGKEEySl/TWVFTrA02Jw2iPxu2XvMGrTAYbZG61CwIgVMIh
OYwh9BbKWm8l62O0m/l9kPzSQS3fKkYXZRFJPPajLAkrSeNk5U5GlRrp1YjrhfwA4+8abJTFmeUD
sZbwWc2/IF1/Y5+o4W6eBGXqbsyoNx3jPaELLzHCRWw6RHLXJw2UdTfy/ZQvOSFnWfZcYFds3hdw
F3/mh/X/yUH4LH7h3gRHbZMNNMZf3F5OzIu8DoS5NeuVJeK16gfjb5MyLVAeaOLcss8nZXopo9aO
foH0a4t6qmJegikkIutAOVCLDGfXRqrWdZYDOebmOk+XtHGLrLbKONOatXlzWNwWPj9ENSy074gw
awuU0LiJhAphNlK7dUSDF22CRGLdup9PifEbp0OpAi56klo9ZxHpyTXk1uFYUyklfWsDfm+LTWXX
eJYp7eWx+25uOUfT7aVUrHjjTdt6xrWSCcTDws20sRVifpAHhniQTH/9ghF1uf0aOJHmX7cALkZb
hOOeET3iCoYoorg76HoXYe1fjB98rxbY2lPAhW5LpeWOpw84YWY1z34K9R29Siine7CfXKIEwfzu
FZrLHxPKLpuN3YvUFMsjp419H/oWwTu0u5JLtXRQtwy0juEMTCHVOzPXYbdHwp3UfLBay1r0gIYh
ytcCHe1W0GnZQEkuv0foMxCU9Hwl7nxbo9S2/NiYEAoPkYmEGxQpbqCs+gSRe1WtfdC1iqy75nWY
I/F+WuV/kYjCUbRI8VF89UrbxNJ+7YmIbCYUXoC7g/gMDkN03yC7yeGSdxyxb7yDO7oN/AWa5w+O
tA9RljuRMPhOrelvNevHobp7tZ1qNuLalwrXdlvt7jbZz/O9yZhAAPbXX7LbHj36HMlBQggOf1cw
YvoRGlLrgO4ZYv2pU0T6/0Nvvi12TFjR7bAS/YYhlYdAm1fAER+1PZk1zWz6Q2X1iPTYZKSO2fgL
X2UU1EoJbNXGtnJN1e0p69B5DCpsmwAZ+JLy6xKaj5htK5JEioP3+KxfsPXBc8/X0I6wS2FnVvfK
lX/vIierPyroMwEeyFWrsm1BXLHZ94a3NkwwQFn8BzoFDFgB0KrKcoqDtBFgLjIpS5Lih001vZzo
PvMraVITlMmTOyz7geHyiPpWWSZTc9nIWX9gAvUsoakQ7/MG0QUcSweeT5Mk0sy/IHEV6CIHuPSu
wpxNglGy6W0hndWB/nsJww9aoaPKuCXyq44m7aIoqeGn5vBFJ2o8qh3AWqIpGVYcMHgGHiPfj+9o
fxihYtOdMG/tI533qBYIFR2LwhYQf3DOp1CPrqPobTa9Q2173YJnv9mtQ0Bb4KXZZTPAirTo7RDa
d9+Cep8wtV5bspnSCxG10UxjiIPi6Rq5s8GeucJqtjClrI8ygYbRVPzc0Yvh6e20qynOmfG9CbGE
fzdRfPZWOTon3r0j+wBWW6xgN/OVE/lnx403IgsSk60BsvsZmrg2aeuE43cUcowaC+XLh7lBHUJB
67BDVZR0DDLSuOnUM2R/J8g+7bTLOIxOV6Kd8L3nIzSxj8Rv2VphZ80K52D/1agARiwVlK+hbuvt
cPbA34UdluWj3YRHvYJj8pbdl7uLggdFPEg8wMvRKZZKR/alYiIiJGcgqI85sXaAIy/PKwCvbh7I
neaw6kBwONWAP3sMSpSIjGk9B/vvPBdoAceYudp8Dxe1zlmjTLVT5A2S0leoExLJYEGK8JFFxFqP
m3ONxiPhoY8hQvfJCby3WM8izUEFgSkHIXa4lOltG1ppBEx1J/0TWo3nRQm28lSALNlsA/XE8n8I
fFdMlGOUUSKhsBLVAvoq2COS/PpxP93/qm0Fgoqm+Rm6Q6YMmLP6buThe/3T8CopI3+ZWfNRxlcD
Jlmr+AyGFV6MZxvT1YedqXqjZZiZfEU0dmUMTsUukddYMC9QEFtAJGUA25kIHmRz40uLlbZ8IwEu
5YQ2VvsipeFkJCjItMlZ5iG8aYDSsnxGtEFh25BRy2uiqeJpYsRHOqXuvOjLr/o0Uz41bU5JzBQY
BfrcxbjqJtDvwNMltp5fAmPcsNBMQl2Y6poEYXyi4+j/yeYbDNjdXDRGqtqejhhRFqm3GQitJNfS
zcdPSKMTzgsOhXpEnnnaADOgQ/wInzTgihmNtUFVp0wGsOqJ0jygdcwd2jtg9y9pn9+iCUcg4Mpa
fxemYnPvfUulJF+crgWenueGjJb7LkzjviL2PB4uniwWBxHtxWxeZZGl+L/Rkv6Qni9ai1WzfnOY
UbiZVo3O8n/e7rwgErplwI7fbugeVTvghmfdtmw8h4mo8c3eBHcx4GQQPIGORKNXoi/8L9+4DuOi
7xT5ZGzB2TddjTgtf6DeF3N3E9n5lDhmaBrfSllFbUIiFovKNPr4Bnm8OStTBTrlSq4pRsrd7Ozi
R7OAUMb3n3Qb4wnXRXaYEkb+pSWy6aGlzooCaqmZszDhgD5YvhpqtNH0iCrZ49zuwNvUHA6R0g1a
nJBD5o0OdWjw3LGJ4MamsirAaocGP7sO44twFbqSn6xuEcnTub1KFUE8OPodD9qVIgjkOyBGFlEy
AJryFVNSrdhvWz/cXrrwQ3EXQfe1Ah6S5KFX32RvHTtJapMZF5FdtknqgIVcA7t0s0W+OJBE2qS4
xbJVzn3pYtbC4gkC0Eml8MOmEzmChd5YA4fppwir8skz9EjOPqUDJjgPBvt1mWg4Ptx7ZYPQSIgb
WpRUNjadSoJ7o5dNpiRCw4VMkqO9Yfhf25fHoQej5UWw4C73IUA933LeczsJIuvFjXSAO/kpAYFB
HdHmntnogH22R4FlGhyQ4wD76+OSaVuDL0y2tgDVjJETxkV8H1HTfoS0t8tiLsChnVvswEa3/vIi
aOaI6VqlQEKQXWzLziz6n3Cbte2Hav8VddT+e4ybV70BPzEsD9iXtjc/DA+uC3iN6NJLBVEDlbIO
P7nsRoX8ne2C489RXSNh9RRzSkbjA6vVQrf2/7YQqhHzJS62GmjzR157yaS0I5o8q79aPVSxFIAc
b1DXlNkrwucBjsqD8jue0iD84duM//LMAvT1hCMTOpJ3Ir55jOqAn1a2vfwlk/iK2hPFzUs4S5sc
e1UirqElehq2qykniQZzozcFyqwm5QwuUvuxKDKx4rrw7DxIKvQFXRRQ8OO+dIXiaOwvRDHu9YzB
y6Yr0P8eqMItSuC1UWsjD9MYFKzPIFI5HFeFYj6j555L0MlfywjKx7ZDUpjldV8lHcCwx+UPFLcQ
sHnW3x6+kSdMXCajD4LjoRhRuPiFgD1kD2K6ZZGmQMi3Nzaa1Lp/dxBRTs5gKq6UankEkwnKHC9k
BC6gT8wZ32BW+7T1oo1j/i767rwRJmNWgPWmaO37hTY06xkMOpBKnuqqtfH+/zpzdLShawQIVipE
JXW3dweez3VAOe0rhLSGyYewILa2kRqWDsnF6GYyLJ4eNGwa0JFDtQOFBqqEFLxj5Z+5LCfW8U7W
6SoikrH5ZIY4EinjOkO3v5aPdnJU82efjwyKWK5Eu7N3qUkFgG3qBLjAWPcFQ/gvnTqKiMbwsBfJ
KUIzf7Sxb3su24A1y4V69LDSGZscNpj6pcmiBz6pgI8gcMvMSd6Nr+Jlf5WX2hvKPy6MFAikjH0W
bNk4PLbWVDmWpZhR3mhwHkLZVR/XqQPqOxyyk485TpYrjToAOfQ/iw2nKdpQWngrTZIsGduZTg8i
IbPYI09wiH5PowAyQZuE7/pGjRonpBPYFYAJDbTZTRF7KpKjmFS37Rgn2sP2uERD3Q0IBwoXjxHf
FDUHDKbxbr6WLE8/R4WiO0Etp1jKgyd+i9Xi4cCLvU0zoUY6337CDn2ru+/yAJY8lGn5dnTIjqKM
o0Mh+jqoLAqrMSuX3hiP2+c2oy8lo1ctdrR6aFSEhAhAVljJyn2/jG6Y6fUl84g17zfJWsCEV13E
uRIT9Zdt2WwQdtiuC6CTOAElfKJLpGhrG6lZw+7uvNiknoRo5t6wGmD3L7iz3Akenqvjq7Xh0FlC
fAi6Ssp4LMJsB4S5/1Yb7DrMOwFqdfI76AhVXTG26g/OCFbTUJDRl1BiRnsqFHcWWFqStxpzK9dO
9btNddoccgbbrXbm4tZL/KmMKhjBMlMX5y23C27yH39y3wIzElOjoG5iXo3mfX85E/CfH3lfG3iL
1ya9pJgNRcs7qVFfB+ngev7FfrtAneyLbq4dqHKUsZDClOtFUFma5YLUUvz/OqzUBHDHrmNZKve/
A5HDFAQDfHk/a6Al6zHUSoHQM0/yIqPzTI0hK3UWedWd2tPTx2yZF6mOXhdeZbul3qheQJqtVHIG
54FdeOqDpbBDd3IeR6H86mcbba8ePIncSvyTIFnBWr7f8Q54+pTsO6wRTUIZT/4UTl4PK/1NKovZ
wBXjLLUb6PiGFZiRLGuh4y29xFKvV2Enhg76qxiqUlee0XnPLLhI7i6RovbxQmYASh2zEn5Dnbdf
coOK+dgufn8oVZJ5MtqJ7hKmCWX9YgRvv7Bgd2G8jw6gpKfc3ETpvEwkMZKsSoH7M7vZ/icc+syN
ArjLaXxZr0kqGt0ehl+fsEbK+edjhVfiJMvBnhi707VirNQDt5R6Nubo+QOshto71eHJM7QqsMTz
TXdIX0AiL5hGV9QNO2lNdP3W/t1yWVUOXaGDptQ+PCrOi1Wn+kl2LnQar9f/TWwo2UcK3VhIbwc/
hY6HoZipxxwrBtBt2OruXnRwdZnhP4rLb+M0jkOab+gIys5b2j3ei5Gd3JnUknBtIOh6RgSe/pjY
U9Ak7SIypCp8M24P4XHtpX9zs4XqVs6n/2E1VHWEvBb+Foi4Q83KSJHRxlCtZEB9dQVMU+lzAZTv
A/S0xrsfZN9MPaiN9szMeESdCq0GC/6T0kzT5s+BsyIZhRs5Z3aUZELUvs/u1pZpKyGm5rh5okYI
QO4Aa/M2CiE1n6KrjGAU05l53nVnGZEZIorhcP/EDqW8RKRoEpttTIdSCKc6cZlt99NCeMSt/HWa
jJEd0ar21+Dnc5j6UTTUmgUOOKKh6b/TNJPJKD9bqwO1+izrli/SJjikA9Y7MyfVjs484mPaXAAT
k0n40JFzaIeO/d0RD7RwQk7O1PaRyT6/kgCz12xjdz3i57yscn6NfGSr80ByZW+qTntX0XPnc1U9
Vwg24Mz7X/ntGtGfF4OuVUAZLHy8zrtyFZ7JRtHup4hsbFtKvj5qLUSopOdNFfJ0Z/KZzuCYxsBB
SY2AccTDdju3NhwfgS6P41ZmInwRjafSOe5GW3qhDI8oc+nahjrdAo83rgoiBBRWpZVsaLNioqcD
U74vuUaN5T8B5j4oepJQohkEQC1h2rOiYjjd2zt9t9wEod4bk/VTHPoeeGJIzJPYQVRsjmUK1sNu
kyhoXbhCew514GioietMcaVgUXQZJBgAWhw8IsH38jBIj/LQ4+qFTUEasrPBW+fRR/VuAjoc/T1K
j1cnZJ7lrhKml0XHS0gXlQUvz4DbUnvloPkWvR5dWXdHjJkg5YtTmyJGfsx+saZ6DLOZTLj47TSQ
i14/QL19ajC23L7MClhpHOmuAvm2ReFLOdg1VlJtvP0r6AY28mZp8sL0kIE7SrJwdnsvNOV1RT+u
UZNhlTpBRs4IDDEtyIW164rLpBLfDIGCaL2uct/nlwFafhT85i3EwehAMQGhIG3N8gmFsH5/jrV/
wTKHAIVpItf7fUkB7+kKbfJPEtaWWmuKMvSDLhuUREstNqRjYpIPo57Wd0LqiOEOoYQJ6zLq0t4I
F3t3IPJTcB+4pP987oPbmG2ByMeI8l19pAijIYTdXmN4KwIrJk/BkXSxdF7MQkwixjCdQHtsXd3h
ZREs30na8JOE5wk3p0bw5nwtwvXPOcMVp5nO6yRz6wV3oIpsDnDoO5WVOmZFMDaA6KyCc2/N1vNR
Nti5EGrReau4SY9klyE3xvW0nw7Co561qTrTRyl1ux07mkyfJyD9JVGC8RstsRVamqyMTQM4Z/aA
xvpceGsNZ+sumIRwj3qjLJ1FdrjJpbZ4eA8cwpshirZhPAuv0e3ZvafvdBLFLs35mz1N9ULXFJmE
fR3GKjofdzb6RrDvOLr0mvk2SGy+MZpIc/c9ui/7DmQaE8eydsUMEjIhC4Nv3Nau8VsUL28TR6eT
rCqFnpJUFtTR2+qGSDLgRVuy711N/gype/K7UjqfUX/JnFE8FJ4w2vZH88Src4ABBBr8kXt2Aq5J
oXRL9iG64Zizbpd/7sHRMDpTEi7LK/N7IInEkZAX3vRilFeYTa0LYfC8Pg3m4LkF9ajrQlMOq3Hk
N0BL8UaOucKWKIsDVa9BDnJgNFe7LmGleRIxhKxEire3/ixN/73ht2NuoBUl/3w60fCIBp0jJaae
2XT4a3URKF00mVDKP+q+n3bVbYX2FDcISAL6+95V6u64zUclO6zBhKYYFqXhNjvBvamlCd+ibaAn
YbkFWppalqrIJWle2k2n4UhSiwyZdduAFSCoaXMF51zYz5MSG8lxcBRhtQEouVPTxDrOtiZIVFUL
Bl0fLD5uI7/Hb857ldPKLr5Us13peJ4TPNPYbsfzUymSQUJbXEC1cmy+2yOcDOAgd8aRJcINfmht
fiDpjAOSWr4dMhqc4CKEcj64LpMtLlJ9fRL8hXC+RJ+K9B2sN9hxP1pkFwb6Us6G/8EGpftiZoT5
T9l3EuvimhMY4HZt6ANFS3fNyApMWP9M2aHYuFnNUUVC1sBvzk1SO8YYiJ0Uv2uNosOXSNjfmp5X
7LKBDvQLqhGhlmXlERbv/8j6gqSw5UDP1JL/qQS9y3teEBZWnyrb8N/QbE+nLvN5Q/lOrzqlUk5X
QA6dKIku4KHt4z1w1Qsl16w3QQp3A2eymNIzTltC3DtW0LM9DCwiXTJDm5Ixe8ls4v9ODZ+id+iT
Ci1dOW+S/Z8/IFY5r/VH6JIExpepwRlUfA0PksuUt60hm458PN2FyD/oGwCietDIkH3+93/PYdFi
gdq9MlLyJNsHMIhNM6+cKGq2L3KWUYn9SegAZTC/hkNhaNY6EixyzZGuuaucVoAzpJ4GX5Ynfxvc
i4tPp56mOADURi0sm3yEbM35JyaTihkDh/JrDI5/vMv1Q367fLjhHvpsgZdTt1WG497JnRkEs+uR
CuO4loN3i1X3O6Irrr4RPGGD0hn2B/Nm8I3iu2mwdMpveLRoSDi3Mwm2k2aInNQ0vws3Mrf/UAAc
TWDLArQcGVoVKCeKF833usTwGi/2AYpJUlC3ZNZzajv63Ms02NZ0vjZs5fYyigxHo3sHmK4cGGpa
Zn6Jz5R5IpVN8co5ln0gyCCPMdDbI/NBvB6CqpO7a9WKlEugELIozfgXXr/sPqdUVfdlAc/H/l/R
8DSNLOFYuTguooqHW1i5fKxj6LFnZpN/zJBTI7PnVlHYgj1u1pVL3ZXyuCDPELiMYxZFVUCnH5MQ
N8xnzwEpZ0KbBS9PiNc1xpBp/HsBQfd47wFSN3yCYzVSKsNEdQKxGCaj2RxJxUp+LQ8Mr8y0bcHw
vyd785+Y9MUK81SG0tyT3WGkg+gJ3CoKB6l21/Zy3KuquWbmKn32UMace6PEk1bSbaDIunxL98B7
ZNmDLhriDbwhhJp4LispRgO+XMUwgcHcMNbyEYNBxrkKEDOBKcl+sEZO/OsTJJAe6KwWQU3rOI8B
8QUaTy6E8XNNna63AecZhDG1S6kD6Ojv3AIXYD2inrvfnvF4F+BhDmSTEDWK99t+WRFOsLHaBVf8
VXyKKR2PhJSSvPaMyrXV6f0SnXjLqVjo9uRiIRpsWPFrK6J8KeW/ceh8pNanWiXwRd2wTfIytqOr
yXbXxjmayis6GHVUJfi4D0Ypk/bIiFL+X9/aLQYxsFVj3zl40PDkmy4BsdnIFYGoJsZYcF/kgUUX
XxJO6xXWD9810rmRyL3L8TivJDslPLySzKf1RVw1F4AC25V5BVEwaia7WvL7+H0sxNHYL5wdDEXT
U3+aTjoD5Kyb6zMa/VJl+qsJBlSmUfbKrRdbzdJc35fqt0F4G2mAQCpqoSfCyA//EM3rG6qcIX5Z
rzG6+e35DJjxz7P9ETtbMknqGw49Yk4BQRMECw5uFAS/scPJEOROHp1F7nLU5Zb+aykkGzH7DAuK
YSvSul83gD+5jjjynpaVtz/NRUZwB662DmLgY1Qd21Acmqn/k8coeyOy9cYJf/iez4SzUNAtbuuD
3RjGVP74L10xYc/KQ5mdbWSn+5D3cHm2ZmUcY/DIRtdxM3XlHiBg7uHx/+Q8l9M4tsgwGSJOxv3X
Wnz6pqjtpVyp+zJbcVQYma6Zr2d1xgD2XPK14DlfdEZuYUguJczQmph4o9TYqo1TkyTlJRwfAuT8
MX2DgUxpGc3XicG4UppmWS3UqxszY/4vXuzILxK17FnpGikMQ9vptfc4CWFUhXMvoLUAkP6XZLzQ
CHhFQ7f+YIC2uNYm4K6UhqwTFLvedDXZ8qotMxTyFxekcHS82MxxBqk4918Vcx2Z2u3LZO8HMeLE
rId5SSxIjmmPro8K77skJ4XtutfM1pHpFVLfZs67C87B7iBEX5lTLfQgR03QT3vrH8M1K2uFys13
idAZ+7aUTBTNdgpHkWy42ARROEEVC/dGfv/edefhcr8ayWR1CHZA2G1drmXxNAX6pmc907UpZb49
Wq4LoLzTDzs7IOYlOwll61VB0fnmVGtsZxUuJmH6eakQEnuS4Boh9sjop0t96cO+1K3+sWw+ioke
btLXjUROZdF8GnqFB9BB51ZM284/aVRHlAHTJHxDnrQIM0Pq1zVSMxjjemHofEt8nX4bOCOfOOgp
9LzYfxrgLcOWcCBVaBY20o1aHgUw/ANxc492KWhynzSt1+Uj+468dXN2NPSKDAWgNjPqMtdfSUMq
qgYlbDLqdIBweO7iG8mU+EXNm0Mlq2dzeDqbd+dz6eAhT2xSkDhAsjX842zMAPymhivltne7Xpm7
nBdhFpGJbM6xZUO8jIyfc9GZIJ2Llug0hIl19fvj/GORYpPL5b8AoOoTpyvNOopyHeDi7dOhZ8Pe
cxTFGLrmPMcX1Ot8K7xfbu1Ne76x8iJ0/IYeFEoWLE5YMvO19yccS+6i8Fgvx3muoJv6JsxBHWbv
oZB22dTi+BHjHX7Z3x9RN7q5+9pSz9UA4TVpAXypVoIJmVROe01HCZFKcXWLOmgukGPYa7vG4U/L
APSrvr4LboBDsNBetXCiktnXZIyTdkOOzgvTvnD+2PFZ8ZbbO8m+t+mL+KM/Fv3JemojFqVpTAQu
khS+zgle3GvppnVH66HRbkdaxn4zjKRzWYTUiZ23yXhMNbWVBZ92mqka10Y9k/YIaHKaFlFR8/8N
omLtwEqgTTIKqugpv7PK3IfLVZ3p4H/fzSXHCYzPNbR2hZMHDAsCcYXHvvbsjugqIh4umC+vrOo9
qVIoC9jUz2Z0Gxa88M0u7gZXkOT5pvdknSzLMttCMNcXw0wNJEcdUJ1f/RkPEGc2/YwOwHoNONDI
GZ+jQdsaigUfy/EFHQ58gTPCr3dyCJ1xgaxGX0pQf2ayL9QDHxoEw+eNhMsda6gcxno1Pnxx5RVt
StAINZiQJFdiy2JIsGUZVZvhnejxxchMvnkbL6NzWkIpjsFIIYlK7NXBAdeZMLLBG+iy/QWN2QiH
HRQ8/cB0QzZj688jjg7BY0pCRaXxxIQU5MfEfvzj1owlmgbQSFAFjAxFp6rmbvRifkNrSvDpt2W/
M/DqFkQMCZYtrr/Qb5YLVnkHtr91lnld5FUR13xsUYsOfZdKy+IdSALvrr6EswCyEgSglScuDNKY
NfNcSEovw9YRfw/q7uVWDJ5AfNUFUXO7ixi+Qjj7Tux5LW7dykdcZg+9yTfzwNz0eLyUJrK43ZGR
hGjGwsz21x/Uf3ePb9YkWn785qtCdBG8qQvqKm7nSxBMMFpH8HtscMnWKeH2l7/gLyT11IDXh0WY
2KJUhDHmGvqV+0wZ0zar+YeQ5cp8RCrF8TH8nCvV/QAicA7guIm59ZivoVG+FhkV27N/sGts3eOR
4OWAwosBczpv3HHho2qJkg9S8m0qK+UiXlczhVM3G055+MPqqFADmF7AzWwlegjv63xwOLQiFYqU
sfctugt6l9Ohtv8n6RmoYbfKaApxU2BVy/3e7MY3tsbGqHZA2IUp/d2dVFmXblVjy0IxUwogPtrH
Yp5lydeRrOAdaU7484j3E0uIaZQlHzsp52OAmKE5bdLPSvun/xKQOZ1Eoh91ebOGF9AYODHJu+Ip
GoJ7sUoNL/s/fTSR5+ZnsJaCZnSLq9NRffZ3JvjNY6ClAR8gUAIAvzeCnZITszFfZ/IrmwFsvJxR
0hbVWjUSmoPR+OzQi7MA3+RJgLVRfTGbRbHeOJqUN+QujUXr4RZpms/wLQGaseCjKpKeJnx/Sghp
RDgS23EGmxV12hyaQBun5Duv+ozDuGY0/a54uNW7Nm95YZUmuHOY5IUCUDn8dcdmyiTLAf0e/sfk
ssEwgu3JjGm2zCcE2lYsyv7M+XQy6r/y8Qsti7PXo8L1PlhyEskZz46vG4sHCo6XYna/Y821P+a7
F2+Dhl6dWG5x3ZIJzMdcxTczjEvlhDkFFNS5Z2AjKegacmZkoq/TLe0/P/18d7aBDB6PNV33ERfv
KTxxqxtiwIiAavASwd1k+vM0uaqYvY+LyRs/6tdkOQVZ9b/3RNYC6i1YvoQssRTPO2N6rl5SXA0v
7ypp7CqxXYDy4WC/lRkhGIrpAqHDXjqkkOYRXB+JeFPZP2CZq1C4EWibPbPDNvF2taI7E4zto8Eo
S46rd/e5LY3SSmnsJRdiN9o3Wj+P1ZsjFyrN+EWjp4vTjYHuejkvWtYD4FjSC01XsLviZyu06kZm
vt6PkfNKZX/7+IOT8A3sVH850RDC/q7L2wSJawqcPXVYPZN5wTeATR/JdnYIw6u0qa/2cp3WJoKS
EsFKcYHhHnLeMzqlT43Fvlb7fs9fy66UzfHd1l02CVQtJ4exNdjNCE0Av23MBwjqko0eYqREwitB
jYY4XpKRwMHoz6oPfXbQs40kZx7DbYFgedbEZUKlr1WZWanfp+u23TdxarfbUiMhD5ExpCUIrQBf
v0Z2C9CIWAehmTSH+gS2b9x2kPQysh4XIhFbBHv8X2RmyZ3RUvSBEQ3/o+wP69OwfQMxnVbZOP0I
mhMsnhrvI4085Gj8EZvoLgN8DfyMHPu2hyHtZ6GjEobfbAnEVhRVXhV+3Bw34/VbBV/Y7ajdw9dx
znqd8mBoDjUY+byg47tbp3AqsZopmaPi8q4a5ujZkAG9aKf1zjKW/O+Ih9JYapEpEda4n9hrAGir
A5xUAbO6M8kPvSUiO8vTXXrSFKL392AT2SNRUp6qTq7tHaSj/L+s6G+t8P/k5shCkzhBdHu1cLjf
F5Fa2Zw1GZIpy5PRGmWwCnBjVXPpFS8p6XXmKk4Png7X1nBuNwy1MVkTHX8uKEyfJENR7CSerT+Y
CUJqN9DBh6KDgWGR1kPqENVS0dij/qceK5Za91thttj6bccgWuB8ydA0qvfR6DKRcrBG+OnVaDSe
MkK6MV4FkzLt5p/oY8y1MzIX27cIVhDQGXqPe8/t2FsYHFu9235Cwq7oM81HNiItRbI7+aXkEDIH
qhZLjNgisi8SJ+L7F32BNPc3wsX6saO9sL71VZLoqc6AcjRvciex7NZM+BZH8+rXVpIh7fJSoqk7
LLCezNoDLfxdWX6GOWdzgyzQsgzL2hHqxXPutP015+uu7hgOzZCHYZz0Y4U99jXyHOBZ5CVCuSiw
XFJQxKzXYj+vwmVOJVriYUAV13wbfROQs0mwFiRfhIlX73WsJO3Xw+vBKEcbVkHF1gnxx6S9V1lc
GUKsaf+3NTnTkV9ZvoZc7dba0q3mRYxMpb52KuLexf3XPo3vc7V2m+BRFwDDHCd9J39FSevtM8vs
iPmFMUdd7leax8tXennnI0TH1j4iZqvnAwWq43zFSlDOewxR3l50Wy0jLSqwQ+ZxwhXQ9+0Wx/Gb
tNqSNCIzF/3x/99pi7w2IgZ1Em5NcAJh0trSheXVGPMDxCFv3scMx9joQNiQPzMkGhH9gFc7dEM8
A3FwxmcRwG8efIe939PkxpD9JbVOYyH6wUVz/wzhzVe08G2hmAMUTlbHJyyLK/S4WTJtYbzyPoLL
YrfdRBJ2Nmyyk9Ugy6nRcd7VHmnUXuBnAS90ePWMecNYae3BBzhbNu/CHK8DAzcJcTpVCSqo2zbA
9UddIl30tccwKsHMJTkS2q1m0GuMBgicYQmLUcJ2cFLXVseHf6nolVxBmhNMYXxCb02ovxb+vPmb
Y36h7CaG78DcIeUOdJ18C8hINsahMVa8u38kE2ed679dseFpC6aE53s2EZJOVNovi+dI1E7MLNXd
lhHfYoWcqakXHFpVGLOVE6h7fryrab/UUPQNnxpGPf/sx8iwbaS4CI8hRLu3cSYa/OUUyCW4EBCh
ECofDvO6Qc53s5KN6lUFwtWEn+uQ6LktFm5u72R2JYF06YZ3A0xHxYlvB2TdatuFbhptpFCWOKCq
Gd/VT9LhlIudgd6zjt8WKjEHPsNvsVUy1zugU9VatSZrj6VwcFpX2XVt1xzj6sLgFSCJFLM051bb
j/md0Tpdjkm1ElLWPPAll5KSt7eWJnJ9vj3CDptDGDi5WtPATjfeItqHxL5OWaQxFsjpGz5HDqmw
9TUg3n6rxLUB+KguBQkWPKIjjX1JQAbZv+3v2UPchBwZc30J7eearXwuYC7TomnQmy+LrFebhMcK
uP2obw6493siNPflBMo4Gpv8aLS4aU2j/jD+Gu+H3D5UvdB0mRgVS/dqzv6IGU9nXLQS/6osBm4V
PirFSf2Bdh1IBv7OGiwUUPlmxiR0UJCAOuG+i23viO4BS5/G4rK81us5SS1HlXTvvzhMbVwnjAIf
nQifzbgGNTD5T9SZ4FNcUsQo43iJYrVP0EYyoHghlUipbM65GyorBZdGXtyMDlqz2prV+7VCfSdn
kSNzPMTccaef1fHzHKnZvlpB97k0kUXIbPWWledYOqIn1sK5503ieJzyphH+wHUZbwHshuEJVkxk
XJWknaU5NX7BZCs088db+uKnjLASVa7ImUbIi4fHUGJl268kbGx3cw81+tO2nV+2BmwyGlb2T/CK
7Cn49aFiRykNT0Wv6vgBV2bxcPxes7Lq2PgQEStjbCjKnAmvBl5m2bPzJSanjfjLlFS2l0ivkrMR
U+TwhYai4c+7QP05B4fYgQJUhGgp90u9u8d+N2FLMSiPCsJmmCosD6sKQyhamqNUUHl4XWSr9b99
COSaVb63pC6L+iT5NTXP9n1kzmalQQvtGrA5jQ3x5TsXAWfXfkX2wOY4aJt0fHT1sGqYWINKWEjn
EwdDXoblHUXQih6QZMUkc7/U5UYvVp3+ZAyNb6hcBfXmCbZTWRRR1//iZM2lu+D8c9Za6GjRUOk6
tMq1QB+jtBuU29KFnHVytohq93b5lb7P+HjWkycqiJfyVC26oF9y+lJIN6pvyH9m0SaCMZ587YoI
pcvdDxMQyrnpwwB/XUBZGI2JK7BtiKeV8nwkRSZfBuJLwVMTiunyDHNtClQcrWQTgI+JucVzFDSW
4EhW4dngp1yotxkXH8VKpTmvkuNdF36GE3s8vkGLTobAz5DKHJVur6ub9FV+GVr2b6KZsNlQAYFr
b180aAg+OBRiK5IY4sbdicggAljtLhfuCv2uKTCEdCckK2NIlZdXnIp1BWcNIg8LO2gn8iQHhaPu
piTvsZpV8l0aJ6mZa8c7UPtiMS8iVN897iT7W19M6hOFcMGiRKtIW0QSfsuEnmgdYt7krW67Iy4N
HBx8tJ3qy0LYxWDfO148UnbWa9wBAvB46tvVA2Eju1ldaAEgQWqocHlu2BqBLPvJTBqvPMJ7flKb
uN2EnNvYpJdSQp3HY+8w0auoR6hSH8rOEYasWv1nM6egLOGo7SHD6qoCfqJwm6u2evByCtH8m5FA
jMxfcfMrr0NWJwI5WGldkG9BMy9hVhkS5kmfpwZglFYSIVdiYV/Yw0Dqy8UWtkinCDNo1AFj1gDW
rmn6LgbcBl4nmxEcvzl9OEgwUR5K9wqqCHzJjuWkeq73Tw1Nf37p2qqYWVkNXNUXsYqMtDZWgZbA
LYZXLgunlNCDNttYnm9xbafMikIwpN33Earao+D3ZSBhRKbhCzT98sH1a+yOJPxV8JvoiAgQCg9s
osXp57SvskQGtozXpYNpAZzK5qBrpS4jrytLGpcjZodH6QTKIh0v6LN5LaxiBVMd+so+mZz7FZ3U
s+0LLBUzAGkaXUK7MpQWK0fVcdpRWRObh2sTtUsvBtGwZvRMGAbmiQ/R2gGMMSTOLu8XeVaDig2d
pNQET1a4ZWSh2EOmDDcxHen7KoFssqGNeN1pd6NgY2h+BTvfaGfhm3FUt3q3pJdXfe+0YulLqmj/
C1c9ojeE/J7lClyGF5L2ONgW0Q8XkZ7QwrkEHU+pgsUSbXeP/YzFFcTitBkpxArZkFFlfVWjyY0o
NpcT7x2cct89uwhAe7pdVblHtTixBjGv4tBllkhxRBGz0NLIV8T5QLxaGOx3DKBOBcfbMc1P46tu
OWhuPrhM7GbISwG2rWwc2yTlU7alv8/q+PdZn817C3aBC6dI//jG9OSKosYzIuBkmlhBFCJnomwb
qCBNxgt7yKdkSHT6xtM0zMU+FtnzwC1sffEAqcMyAXf9h1zhqPvMuHuwJHvWrO2D2eTzQYphEI2q
4D16jn3wtmTp5lZkggdJQ7953EGsyiKGz/3H+k6pmVW/RUL4YyHLrl6z8t5kKyZJnMJUBT7UYiVq
7m/mRt32pW0IUqOc+dptF1toGc7pS4dy8AfPagxIpADviUWjZQhnbZWuI4X37GA0hueLMzlahBJx
VuvuYJpMu2Ba0EFEcrNJB1fwCUhGUHmzvrBOtyN/lIJac51cwUoJp6nEWGsCgxnHarafD+pfV3NJ
u9JWoD1jnd40YLLsz/cEZZPqkHguTCElvmHbniHvWVgq+LL5kL4uQVIkEr9yZ68yfXgf7LaeBP3C
8ASb3T1QSqkMDK+M/vBnAefkFH0ny4MWYZhYmiEbzqQ2YBCCYnllHeh0owLH4TFtVSEtGYto7WP2
qtZAHVf0KZ8wKGX7sdHtzNlDnS9Zk1FSunD/8lxYPXkimA6HmBJtmYt8GtOVirwNE4p2lu1kLvoN
KGgdbxDmyiGgBfCRogG8wD6vbpl1pOswQ4mhTjqbIV4JoLdVYzyGFfJE8lNpW+VL8dXLwByTYx5E
cPhixXwvVwr8l4Ej6IYCxmon472ZW29v5rcMaMJO7//F0ELbda6iiAG0hBSroXMOVSMajn4pMTt9
3l8/5ntILUOQ92M4HyaGmQLDvtaFp6IPggqH4/c32PdlXQD3nSihVbJpXc6FUpOGwm52oOxfRdu/
U/gMyN0fqWxoM+BrXZiE8s5mxMYRXLLs/1k33Ui2ucxCZGXU7J8t2u/VUgYAHCoFQTRVF2NPMp/p
u+ezvqSzBKomkj6hRBono4t6l21uDBuoSqBMt64YGnUyhpP+VZr/R76Lr7JswbG4WH/v8zVVzApi
cxG3aC65amOmdPF4nvkMFRMacRWIikzjYz22CkVMSBhWiBDGZlN55RzuODshe3bQvWivQiX/FixW
qXNHRsRo4xG2IwuGjCStIHf8i5iClJrcVEkFUI4Y7+hqNOqh4vwk26MpuqDe8yoT9ivTDKH+Fe2z
toh4neM85L/9lJvMV3Uj28ISn0PeKgKS2kfqvmOKDYJZSN7EvL/MMBFwJIn2t/UhPzXu0XVIBVdu
XdVrJqAPDU0SReZ8jMlmxiRAvmHgpfm9LcT5CXXbALLzICdDjKQOEPdoA0zeys/k+d5699ZpzbpW
sKIDWEuFzMgxBIAJGbthKVIedOpUjb4efTJuqQmfO2ujnKiA6rmoGg8J2LRU0Rt3sRimozQj8wyw
RM0z5m/7ZIiqFe1/oeDogRVx6OZofOvkYLfQVKEoIVCX+AkIuqQiIVfAFv2K7JIr3GJblJoZKxAb
l5rTw9NAAi7HEgOLf74i5MZaENP0guZqSoDp6ggCa+eVd9llXxa1CK3CKKr7COhZ6QXMOAonLs6n
gfCI+C45eVOnQNul6KuBcvCCBVdRF0qv3rKkUf89mQZLgjzQ5ZU9a2fVYmpoQ9KP0ODdDqhCfJ60
Qygahbeb3ey4OGJPdn83panvhRzSjI7sh9voLHnqg9/g19EPzdrpXphY0aZ6bP7fgT6UOSisMEQm
C9wdHogUchYwAXL5yUGPevZAQS5K4ipfsza/TjODLwIh3CPnU2lR8XPDIwfhFjy6MQmEL/xtgUsn
A8rbFQzo7BYJ6khoXAdbeCz08ShrRprZBOpZtcXXFdGCtJklpf/58zdbtKd/bhLZIY0Q5TkSTxmi
5aPIsPBtALemwg4daDq1vcfzyT9mWWtS2DTvlNtf2D1scnRxs6HSPCjgBewcdlMcZR5oRf13muiz
CjsjpGNs2WbfqvhYnj5w1Akb8G7MvSX/rTmDvqA4CAIMLDMnWdSotINz3WCUKpiAPuY4r0iz9295
V1TzrWiLcgXxbgEM+wlzM+GnzUj/Bhn7bO0DOcpsKKJURX0oWgPTJ4UGLxhdShSw2+4hFFdjK56p
4xXFI68BgXzyB4CCRu6FF9xsKflUSWjWjRnRQASO8e+gQMgGjzp1xGMZ9AxZeBJaY8nau948mBT6
yuDlexmiQEwKiXhb+xE/RqBFfhfcwvpHmLTKcgZFXzJZGJIQsbfT+e4MNP0YSHbSp38KmxaB5tNp
lG27UVClvcdK6fQzl7qnVoMM+6M1zAXHXzAmbjMR3mvMtF3YgkYdhr85eE1QqvhO6Z7oGJhrdv5l
1Oa6MkBSWIqk+YIQArtLLQDqe9DtA/j1MzuUM2qcwDUopnbF8xkTPMLfoBsHPamn2Dd+oT1zcxW7
K6MeaBrptuB66d3GakLMuMtWg0XoW7dJczakz3+39RouSJsiIupxsc1PLg8b3/RLowyInHVV/mCL
cj+1VWweCaj5t+9lTf28irlg8fI6fAog0ZqnIPwayOcIM6PBFAqy3yom9NzDp+tw66wKiB+Ds59n
l9dO6Gm+HyuwdqNDpjvhn/OgxG3vNso9J7FpU5tQiNoQUKqQRcBbGbi/0Vh6hfVBSFRZJWSivu+X
QTkrduBKkS/ggEUZY8fRjV1eupzmzDOkBBdJmcKdfVOhL1jyTBhuyk9OsEF8StP0ZIrmqUr/yxz2
/HlE8gaUPDp+fP2fQxnIEb7dxeZ8NH+hykgq3FOAT7/hflCzCwnrrjW4feW7B2UDSsDzXWCjhoLr
b4l951DwCuX6q3sISanvBV+Y/4FfayWzSOi8dtL+lg8hKgdTHSAni27AGUbHbl26pMhmXadhvCsL
KRzwkVVsGu9wtSBI62eT0X4aeSmzVcF09quY3bRZkVtGGFSlE9zr/agGA4fkTveyU9mEaPM6m2Vq
WOz45kpUNMwvs4bD3t727S4L5sg9T8o5+ghfjnHKNnfZbepvgqugbeYHqLpWcOCAAdtjO3pZ9tmS
pCVnlIY+LRJDZpyu4Thy0LmdBnvOQXHeSnMhUvMY1mEjCekGA+LQ7sWw8BMf2xPUPu/pQx+3JnpC
r8rYeHrhwHo1KvjFy0Kcaw+vbIIeVrmJ+zKQfHdIxZ81rRg0eyhlM+A+bwXb2WZvwplihvwxInRb
ipehLF3Oz+B/TeuHWULlP8iwmvaLHVy+MYnTnJcrFRInpNV5f2dz+k2nSySge/qKTg6lJF+LXZc3
MK3BnKMCHOJHe4X285LhiH+WNG3ICN+K57GyL5PRXRYlDQCtMqkKSI2iBWaF/8iadveOmZ1gYQsa
ow30AySFF6upfwPFNdOAHzlzGHvpiv9KFpXH1B7JEYO66QGFtDCibzBgNjCeAKJQHBmWb8U7rENZ
VzAwOgzyvhU0Y1jHRZ9F0CQ0Nisrxtq6z9apjv+TQIQBUp+DUj2Qttr6wNRutwJSu2IGTZlo4UIk
wtZhJuSHDN6ESR+zPX8ZYtvaeKioc1NS5q2WwRu2guEYvPT8aNyq8xKO5CnkHifXBnvVAxApdZ+h
A6vdfLcu0IB32qUCPq/qNmBpTYQvVkMVeBTxt0GA1+1rKDe4pYSmMZVDEkv//AKEC79mXPMnRQEd
IjVu0Ii0CWw4j5wwpemhgflRTQ4tcMDgDAhboLBUhOH2+bnzjRr7Lm/ofubdGFqJ6XMs6pElSxAX
S7Q0v2wsk5quVoNzPvqfNdWe8t1RXgs74Fi1usBuGZPVKExTPZLhAbSl926uZW2M4TzNlj+n7s3y
aFwtB8MsgaPYTxlgBS3VMYszvPPjlv2ussmt3CjE0XT0yXSvK97ByqvCdV9l5IQDMOVGecYGcKnv
fzqBGfKu8TzVq8xwl1ehECzU5F6kaSBstp7frHUi9Ft2mpUxHpAb4ce/7HgYd90fJ7xPKZ/Fe6Q6
cci6Cc2NqmCxQYvu49u/SgXFhCBTP3lsNiYJIaE8i72ws/nyw8z5pgIhxFM3BTq75neTCerXaH4d
ZwTaA2wYUBGHIl+4UyKCHd7pjCsa1OJNq1TqEPDWgvpMfhzB+2zpWvEvjLNsv+yChIbHIeRyS+Mb
SsETh2UN0YImpIGXV0/XONE3/eGFH/aaRU3Doa90fI0cIHJFvC1CLlt6A2btWGmzijf5AsEMPg0+
v8/YkPg4ZxxP8e4HSY6AHSOMkAd40UqM0DCUthlc8jbE2Qd6QzSjhkUD/dYPzuBMIg0RBiKQ87WE
pbA6/MREcsquKTPuw6jW43jjWWGhhZ4UUOuWl+jIAEvll5PS9iBBo9bNmFnmpDu9xBSTBLjxgUrZ
Ih7Kv5j1hSAmP4wRUXB1PuypCdpyVCGH5Dq4ctcgo3NC9FXkjOp7jdaH9JWekfXubSO5MNuFZkfG
u5NNARduj4K+SdR2g77EEFUevHAc9yBvtg57Tn+fXEowMLvXs+eKp5CT6cw6D518/21aSbmBc29s
mcYHwgfIqBuB8moQbEXji5WYbd4CqCSMz4F6+r2THbjIqnqGmFb3/6VgFbyx3eUtiohl09XlatMW
U0f3JRpdmuFyttNNB4B6ZQ6vNONcEo2ucHUeS5ee3CaPCXZMUfsj+i/o3ysJpKbSf1Fb8cCTpWS4
W1MPFSvu4WjRv2fuLF0q5zRQPFRHvtDR2v3u3BuTvGz3i99Y0CKIMiYPxumqkSGjpMaoODvhuoyr
vugH78gcrUuMErmMQHjGGVcBwfre2RFiPJ/3xRwMe+mmahBTJCBlAKShHdPLJHKRYtZVsskqYOxI
Bujid82eIe61B6dAYvbpdztntc7BeesWH7ZgWPSvI4pG0ywjSUwjxHtrxVJOnlUp04Wi2IjwnM0G
DJilw0NQB3z8zNpU4QhSbN9L5US+TkhrlREOq2JbSg27Nr2lGv9gVxEcUMjT2251eXJJU0FDkKRb
OZVPgOWkkisofwxrSCicyTMQx266387GGS15ZuMpLJV3Iy3bEOhzPrGUe/NMfDI4/6vbohSfuqlT
U/3kAURN0dONoLQCGQY/XKUDU3gYtydSu3cxqNBWS0zlHh52q8I3GJZjWaaMmKJAY19w4DjX4VFI
l5AcClgwCWjxqpjfr/q6P3aIEYSEcl8I7HekgbAL6rP0j9n2q+sdf6bb+GJiGrex9NN+Fbhnk87p
RI7LoILh9S4claZ1K4x+YylkLIZik/ybiNPMUdS+XhNAPXinI2n+a2dEbVP1/0zWXh9KocE1Yah4
UdGu0K2CikYDXW/3JihYwtZQ5Ja0A2xzC49kWVGPaquXehzVY2FqEpyBKulg0PLm6FN4S4+c2Jza
9obKutLPGKh/G8x89+9fd+pcfvHOq0l7XcnhGT6BU37UwW1iFOTkZo9YC60oaMVRRd1BvhSVZqis
Dh1WR/O82+cvIQ9b9/vQgHq0Mxv8/LIDF/jS4hd+3wrmV0NjoQmWh8FqVnK3vQUmV44pif8oFfVR
pyqAOoskuFvKBx080eRyL2ZJbdDKvvzQxKBYbSTwIBxNHgFc/MP9C2px7M0nCgz2aKt8QedbJYmw
Z3OKC8dYBorKFK8qlzOTG8p3bVOhBMTCplpg1gZ8OxT1SP3RJLuz0swAv8MD5M6Mm4vC5V7Quqlo
DQbDLhuHm31rjSIRBYORgFPQ+cInlbnxY68RdfiAVSW+xluKCArJQE0t7Bihg++qLR5NZh34gG6C
ZzC5/MFIVAAoJDhj0L4mSF1Yrl+/Y6RGe6dhzI5krPSEdDusidPG0XPZr43YElIyFuFHXvHlwfi+
EGTQ0bSKMP4Z8GHAJ4jEMPo26dDtud8Glt+cUkbcgJHewGuz0b9AqGIANkGCOFwZbWyomQgYFbz0
qDALsHQ8Cw2ks/p0HLRDJuariSqvdD65NeXBo3469DMcRfSxfwSC5UQ02LOnVomEXtrMEQ+UfAgo
/nYZQ11J2LkmusUxCno9wb0POmAdT/lu4mL3FjjALwUe4vVUnrDKLhRDID9MoYWyA87+lNi0Jqrd
fwd+scfVfuWNH1C7taw0bfQdIjDjqwrZMPsVmxy9oaH1dDW99t+wDIhVI7/VkUqurSX0Om/c0tQu
0e9ke3WAnuBuvrGJubzUU9wp07CUqGHe8mBSzR7vz2Vz+woO9S1FpQaNMLks16a9sy6QToOvBgUF
soe78TBlNSLAmIvDSKKkgetA9GF2oTvQblaqFnWX4B15iNxOPE+EA60o0iwQ86gqB6hh2etbLL5x
qv6T83v1GmAJIHyiToq/x2dnGB5vdZN5rKHGqcVrYT9oX5BjNaqh9Uqz15UVQ+WfqEl2p9z5rrY6
4cSPZO6RI9PwxJfvTNGWEvfzG6l/fXnAJLnxuEwx9Wpzjd5+kDmuY3v3tfo+a7IYu2tKzYixUf5A
12RfZ7f02dP9OblfXSduOeqNI2kJpIiEg5ld7qbrg8oVqpXbyBg7e+NZYmFpEg/5HBL+PenWc5Da
ikMt1pZHu2LeuG33crziNYJZ3IcLWkcmsQyvNPsAVRD39qKY5B1qa+BCeeoOqDWFyY0Gt2IyYD5G
+9Pz8iRCt6uL3I4K5rdqYgsRni6H3iteiBN6MRvcbHxJD9u7coqQ7/QHRYNk/VmCaSm5ulxIb1Ht
jdeRvS63AtdePsVct8oVkIek1mqWpbLtIDZQbzypaVxtYvMikRyOBY2YEMyhSUqZbX92BADaws32
DQNgBB1RHWqYnjgY3g3NLuzwuUPMf9DLJ+ja26RpbF3ZAj0nuqpA18M4+8bExLiR6c47MaGrJN/n
GyLAQ4d2MdKQD3Rum3tV/VPbtm7GsKZF7a6WZuUTDwXlTuzH/Ited4NamMbT+E6aK/d8PwVa/e+l
cSrDwJRUO9n0/jLcJZeA44a+/vgxgdPClmg5Ww1FhELLKk4pVj4I810F8chmElSzJoaMucGRLl74
TVQ+7uxfQq5hX4g7CHUUTiypgJvt1vvUhouuxmndPtdJp8NV1rDhpWUWiu/CmccTqTt1bwb0uO0N
CQ0Xba5IJriGIJIsS6h4tQStPU3lejeiMQ1fZuNfDuQ+0taURp/fo6CnFqXA2pWibHofgd9jMDr4
ASG7M6vUut6fdfQIEa3fRVgfB7KjJxlS0PYkSqYFHmTCfe5++HaMgXFVndQfyKFNa8aayITFz5BV
YZDq5VhTJFwbH9dO1GCAf9REqvlB7PWwTbVhpzMNzw5wEsqlfUV9OTduFXDMXhmvZzBy6irFHn51
r74gopy7eAGtBCi1bgvq1mPBU34m7O+Fss2Q53puz7Q9ARnDg+plhlq/M5sh0RdAt721zfUyGOcY
AtADpC3mhaF2sBZV6eBA1TrRYzjImlNbH2aVFJRDZvAAkRM1mS3CnNk9GAW1bAx0uphJ5kMXBEgH
PdJSyO8cfQdmWBvtwrVNpofU/fj26v3XISVP9Mip1+ovsa81uf/gZc+YSLz3kNOkLqzJ5U1wgNrx
YYX8Ta1cX87nuc6HftMhsdD7pQ1w2+n/jbH+b3dwSn6dk8XkGl4MCYQufHjtJhww7+BbKedK5Pvt
pvogD+kSUPhuTRSiKcKNaqG/75mvUv5PrNqMU4ZFqtCc4VcWxIeh/f4vHRl+tqypsREMPLaT5KT9
UIFfnOLEjcv3DDxhAOPrhqq1IwSTIQ9U28nBZDe9lyEaSWY+A5VvKVTX3w/Il+ecEolJzAM31A74
06GS0NzQ7MkQ6JjpOiPNs+POktL1cHPbQw8smvyf9quskQTqvIV0gGKFP2keyGWGTNuv5WxkJvab
tx3vD0QlIW2EIMS2uiVJqcJbTNgOX0o9g75tBVRSGlwYGTJ7eROmNccEq1kA6BErDQ1zxt81qCMF
gmWT8uGCwy4+1rC1vBZ0lEg8D2GspKMvmvfUZh+BQWajGx1kZ7ZaYV6XPuTnrNmuXuhU8qiH/v8A
dYFb8rMtAj7JMErmT8iLzMf4V6OJjNyeyJH1MPqU8GJ4NkUETNVicAxeQq9pD6UFYf5MOrCMkhaw
k4VBcCRyHp08BzPunvOo0Nx6YygNFJdMDUmICMQ9LxGex6Kv1WOgPfZITeNarUu70AmAgg9WTc4W
Nsq/rH6cjMRoTEcTuD07M4AJ3LgBceacJAtNMYDeYjXIFlPIG9orXEGelM3d1XJPf727vWOsSwYd
AncCgDoBJl9/QCFBjTqYMc+sGgYr3+/Zyfl+ldTxHqBhWCNm+JD4N0AL2VdDg1ChIBV/gFfRcopE
SKirF5ffyqFli6vZ9G3wg7zjhNniXshxK8iiY0bnQRZwAxCkr73FmZEJ2ZLvMbk7Q6VLVKPvgWC4
CUaZTmXaSHEpWDKJEYtTfrsN4TdfJmoSSCIVbKXJbgwcpwbBPuI4aIOntbMwTArsIZJSOxWCwafz
FFao5UTv3L5i/XvAez+un6RdPngvl+Y3ExwmX7yitrwj5EXIEaUodZ7Y5PenbEyjH/QM//eF5hep
MPoRz72RPKE2M/nqx1ZElS3iPpdLDimVionDFb5FlXMMKaNJPS/r4ofe6hoTqkiLJgdNFYVHgdA/
fzRmsjC6ZxnRAhExj4fGMoMG+ADPLT+XBpWsmWc3vmO1MLliQc1DDy4hFHg7qokriXUSNURnLzhy
l1KemaDFkZDuNABlkmIM72bkPau1NyRrV0rshY5Klwm1zqyl94nTzf/r8X6UjK4FoLSewHilJoLl
KJyRamMT9fwdHIxSNjuh3zh5cWjKlPxz4SGlRlMbnTaY75W6wn9w5Jjtz03ZRps8vi5BE0mkC7PG
vyd1dLL7fNptRbtom1fFQISM/zYXG9FSKSqfssWaJu92P8pSXvmazHkeQ07jRa9E5N5UEPJqX6C9
doTkEqHBfGAk369WFaL0Qp1lh6aEsS4LUxQjqVH5dyzKybTyzxY5GJvgASdxGnk27Sg3AWetrElt
URktZrOuJsUQ38Lf2+k7Y/E060GFfUBMsrJhwjskfk0rWws1NF2N7Bq+2qBKjU9hZPa7/t0lrU2b
bKPCmjE5eGyzIyyItK2Lt9cyo1HrI5EovCEIj3BhoIIHJ+tlZ8NT+bOy21+WGMFBCWh6fdXhE1Iy
dOmusxLack6HWFbBnyISG3jJ1jwZNGnzGwFhiovT+NembvnVZN8GquVROvpqvk2UvQqBkPZ/MCZ9
X8o1xmseLxM+KAiGM+R/dwGh0agpOt9ky3X4876kGZ6d2p1IjXHSYmyeQBpVdn3NRircL9b2JKIl
iwFSfJuZ5YB0p3jpQgqPDiiyDQ7vSa7SBwRIKzGMBAq4nOJXzJW8H6RJA2FW06wgZW5AS+314w3I
SDM9Ceh1ATI/hoBJW5igNK5f6NrNzS1o2NFlNTy8zZPlodpETpZmmiDCSqYipzIk/Vo0LF7jm9eV
UaI9HnQMdLBTozTeksGoiMK5l9JAfCRZvvKdAKvOyYRgNX3OZYSru7iJmADwUZFo8qRjJF1+s2Rx
x2XHVPIdC36oXHOssQBI+OhCesujeRK6P5V9KJ8DbBaAWruvbSYtW/RRjXuH9MvpGQwx7U+mB0A5
EJEFCAD7/7nc6DtWPC04NLR5sZI+/bENm36i2e0uZQQwfqmxzy6LsPwYQKaHLVTj6nBLWQCitxuX
GniZ9kftEmf5j7mGVTDJh9tc/3o0rMPAR74VTqT1au8OxzoNjGHcN8g7UF8AnBfoLrzzTowwg1ec
zsuPL9IcK0cLoXDoNxvLkVu52kKz+hECJgJUbB3PEwR70TwR5XR3Kf7dMOrqJcmh8hF6tviCyIs1
xRBkNazauy043rSG8QCq9VHzbs5h7mXhs0eeSaa+OA/AxWPX3HG1WmRi52HSfQ8jq7ejuj7gCI+/
ZEJfhnwx2uhAdNnUB2HDH2YzsfNxN/7lagXnkZ6sxGuZEfHU1xs0PDKS1zqehAub1iPmadkVM3bJ
JqCi5k3UHR6t/uK6DQNIK8d0oX0UBGa7TvQ/R9vXEfzzvNSqEEIxeaX79KFgR/bFa72pemTIM/fA
LDyKHuv9lm09v9cHEU+NSVpW9E6ntREuewOKa5UR8cep9vKdoNNTWsjI6bfZ7uyq0+1hLIVDxH4L
Rx5JX2eeFKMvB/q7l+9NdcgfBjK1QylLXN78oWW2MwWfJhq7Idhld1Hces8t42uiqGhY8EDEdfOl
fsqhipoQYcyX4r0/7jsOZVOAmaH8EIWt//fjbgHWXXe0pqHHwP/KfdHC027ACHezlixGgBKJFRl4
XTU8DHtjejVbTlO02k7v49jAjvl2gK2I4k8bfB0E2V7VijOXfv6nwDf0gPjoAb4lSZVXG7/JnZzR
BKqeGx6fyWhFbq2u+l9jeLKALmGyroyp8TZFbPlxTrVjLXWtrEFPd7ESnGuEQt3z73YyEDwalIb1
Nsx++ITfZJJJQAamWVBLtT/KflhKa8spe7t4mQF9rfcdjaA5SrR+8mNOC5k+FOyTzMPyhjVh/lN7
8+XuSxtHKx1WmhRYGZzmSYFIiR0o94i6kfCsYpNjyQX2fYi/2c8RIXDwZB9LdrVYJUiNrmfoAbcM
ZGsqN/gS+1QpYKBqg6yiPGV5cyfbIARbbd0mh+bk7hkNXKj3hqVNfBht/kGrWA4h756jlgLfnaOU
Sag3FPHD1pHGTbFg1ShrPhwVJ21Dlzk36R8KbjunPT097Oa86PUUQK44P6kQhE+9Xnzt+CpToFMB
k37UQWn7/Ts3On2RH0ZLkXLKbHiuLgpnW7c6p++U3F1i15qt8Hx9S/N9u9opNlVcTGs/O3zYtz9R
UDCE+Ylu1C9Tx32jrabDv2UQwBhlsDgmeLx20Cx3MyI3444aDP0nOiEYLSVEMjKwpd+U+sgar+tJ
mVdzAOxcx5faEaJA8vN9ILXuyYHVGKfacL9Y2KTGhy3ABoNr4wG63BUXdA1+TVL8x3Otrf6AX1tp
MEPoed7U6yBVNMNfub7Jg3Z11W8kZOBb5mgpzSxIm4YkA8aDIvDT9aSpMUmXw4wdf1GxaygZteLS
8PsuYG9VhlL4le6CPJRUayJfHP2g66UqWySOpPyzY0E57XVbS152c61GuH65KHhvKtKQ7zV5F1LL
fFxbQlsOtfD/9v6QSs/FOSJ8QOhNmLs5kpKLiMyLdMoeRN2jKyttj18irIVKk/8VLfm6grypSOvi
UoqaUjNXxPcbzPxU0ld7fsyAySZJq7QvUfdRfF8FSqcWN6FqZOFg2KOcrJyuSELzKgzr3qzOTHjU
fwWGAI/t+R7jkd7eDyq+HosNlytFclCbkD7hSNB7URZkusYjri/8PXIlTlriaVLmB3yv5gIRraFi
A9A0F7qCLo86UqYCt7pw7A3Qvo0/S5vIyDaN2UNnxjOkb1nojE8dx+eeUmy86jC8NJxUMpG3jjFR
uw0ga7/skMLvrNniCJxGGgJ4WaRB0Cfkv1E9A6jHs74/GoyAFrnjPfD7JBsiPbX9MNpKumNqxCkX
LxReWNOMP8O/hEu7R5rFh5R6wuKWFxSJv0JRgPqobJ/jEk5s4ge8zaJSNI/QpW9HgDx4YE1qP9yT
2fMYoAAociDnHCD4yWpyFrONJUkVuu5OMKBgIK7OIOSrjnApYR8BxGGH7j0azWT9jQCQIKbUP+jH
688ZIQERRk3a4HT30U2/3UePEzWNdBiupoU5OZgCPg671v6xsUyoMH2ujawKa1PEF7xNi5bYPVT5
N/FAGkxDZdETDT7mxG8UfCw3StCzqG6rRtRn6OiGnIdQ5rhGxWiTrApPABJCsIOqffVAyhW/j8mp
9L8kYhG+PemZA14YcA7PK2wIXKLi5Jr27nZPdfMeURL98k+cQiRrRtE+xKESO8FjIJW7wLHCc7M/
hqYt5gSKJHsUdXDW1kCgUM0MZ/PbsPZC0PcytVf9sFCJIBZaQG44X6jIYHx4B6L4avUlnTKoU7Wj
7Zd5BN77WPN1bhLDou04QjaOHHrWhtFMElkjlX0UhfG0rrK8ipUU57HgV4Hvly9bn5qChcb/pK6L
VNMwUm9ggvHJiaVkpHyZTTL4rzEUvORfflrlOzd0ookI2lZZFfOLHbsl2r1f+Y5oitXpet0HGNCl
/hK49vPSUsMNQelH+QXsUFJ/KU8AovCpCqVZvvULz/bEoWHen5P8TjcsC6IiHwXy3oXUm7vMjmH7
JX8Bl2ir51Naqb74wmiIJ1M9sbEkwYwh7MGGvASdBWkiF0WF6D6g9zvREl3utti3hAvQYVscFgE7
0bRCUt0tSLAIrc7rFi+s4q4MSfKZ75EW3GQ+QliB1stcavfqccEtLPnQ4O+tUXyr0MdczKwDAwNz
A3sB2N+xFl9Gpqz0BuDB2YDiQuHqeZYiDhhpPq79nROkACU05BH8m2L5Q5tHyly6K6GuUF7sH57S
kq7QSRPwxaQwR9a68P4P5XHwFhzH0Tg3rPqH6SYKiT50EGRlCcylUjUDrMzqu+hR2gjgC5H9XEjv
NJTiSSugYLhXbtnjRWu9FGl9hi4HdsiLsDBf6veGzUnAb8Ph95CnsIKbgP0J3motvw0CxxUScsCL
Rb1Un7dVsozn/3sy9SfFe6ZuC42JtQZaiVwutyrjzur5XEQ9ShXLniJvJPblzdcVrbodp3XjuS0D
z7DvwglDd7StIOhxIkiZmF7yqynQgLkiVC7wxM9Ux7/MocpwQjixTIqgwbsa3m3rx631OSsSgzyP
TgJIUqbU7YkiYldiEfVRpJED5zJnEdVD5D+15ukGDUE9dkw2aqVal4huWAmtD/Pd2zdGjxpImAZf
1W/NuAIf4GW3jTRS0Jfrant/zGxB+lro7YMEPBqy/T+BU3vI/S/f+XAtxNXxyL9Dmn+rK666x4zG
4r34rLxGeK0T8nN5yX2vzOhwAb492m6beDwT1iO0oIgIGdbav05Nrl2tjz4a8TgABtGKo3ZkbKM3
u9hz3nXL5YtgtIr3bRx4ImYr6u5IIYZ+SgHvAxErRue9GKxGlIOvu9/FDxipuie+RiaJtgd9o6wT
HZj5VzhuSpk2gPAsGZBk/gFk8WSCMNyuJI2yqhI9in9RCxDouLjkwxUeel65hOiCqTam0PP5CyE1
Faj0sGUCdjXho0p6yEpk5ZsNh2WiVJVZKbC6gtSpoiJQFGsrcgE8PIxNEjYyD519B9zMvkwV9Sv1
3RyOsLW8/aH1zwEeqjprXwmDxPRxn0mZe85c30uYzPdVl4qCvxoBi1KOv2T3pTkDcYAuhCsisEUN
Q0l8C3fqoBP1gxGHKIgz0S7CXQIiSNhVd/79LsRiKNLVM8ZDSXUIvq2YNaIn4SbWJ4mL02T9EJNy
gUK98oVqDgbn2J6v++p9XfOz/oJFCD2bIv6NNn+rjOzINkgHvr6DqEcOBiVmUG1uHT7iyL5ywmYc
iF2Qh5Is5uKh2RALyDigW1nitcrt/LxdcWBgFbNRtGsXoZc/uhpdeb/pAqwDiJqkrH6/UtVG5uqf
a+zfEEd2WiuqhuvS1ChE7VnSwBxgRQ4nDZdQ49TuPFQsEG0rJ2J/wat+oI2TqETKWnTQJcKlC+9C
AKXim21Z524Jn5CDSlckCNC1r7/dveG5kcjxxmN/ECJXHRPLt+8hzLJ0SItkTDip0dql3zNHJUnw
TGEh4wZ8I/qV9F1JXq3VuxxPnDSDcCmKj0lQJ8XyYHDv+/wnix3J4HzH4kkBS0RVGVhOEniYWHRr
9cb/nd4vMxeD91YSbbnEmwoix787TLLLlTDXf/4DyYvy4Vb9naFgSpLvs9+OQH48Ea0hx/EDC3KE
rsaFejv+64fpJnl32YmsI1Q17i+ZLof8ZfYzue7hpq/dWiqAyRRu4COg55FUzNkEcpY/KnoHpPZx
Ox2G/XJeBel9n6Qfl5HPoF4MG36Um/Kv9MQpo6BVmaWFGHK/Sh3LMMXQtIWeG3CLlnrNhXHkRVF1
c0FFPOC7nHL9bkLcmLV9SjFSO4iDAcKuAirnuc7hscS9UW2zTUmzjTeaBC0ugsbRIjBFE4Daf1Lx
rVEvfaMYY9N3FODzrALWVAQxU/P8nMrF/2V9n3kINDSNN3mKIjTpRPyc5KiN8PtaDjuJVAdgAt3g
2xUhSGDFfoU3xo+OVe4wRFeiy4crTye2EcccYzjOIFMZs4B92iJ+U7i9n6P4eIK6IAbGUVdO2MiO
PfP7u1PsNU5iVm7jCwrYq73dWltE6IYKdC/uzdof7ta3rI6YlPGnHiVnq41wXlg91uC+xJVqZkmU
u2R8XaHkTgjxNUGwE6NKDDbxnZfkvdfhiViEkyEZyfETO5apCdjxlDWFOAedaFJzknyZwJuRym0T
6lrD+5bBmckPE1koNBtSqNMhKJ/eOghIeuQHs/KbHzeqo8wfhQffKp5z6lCiLABjbdhhKCElwyYi
uf4xee0ch0tYEHVQksy+ZbYOsXhaBgFDWlbGaOPtCZPVVYlsXp4MtO6Xh6yZsXysX9WKQuSXFBH3
k2HSlIIaPGQmC1NuGiEfwsM433c5NYj2CpFKrZQYB+EKzkUA8WbUrqRYvtdT4mBGtYplhRbRr7jt
m8flYd79eLCjRLAeiYpc2TNhTsgOtO9rtSZWxIFH4lmWOKt//vndFbRNevsedO5q2Nl9HIoNJaoK
xHLr8+uZgQhjPUKUxlY7/1xbAyMloF78QDVkbwmxiYX4TMwA7iL6VoDz/q09kg/y59Sn9XaPOGy8
W2PvQYeiGqj9KNM1kRWKmG3G2pLse/mnqLBPopMcBDk6+HAryuyNyfe10aTlK7tEMvLFVP7auxgh
GyGkf78N7KD8dNTtfHsIT6ey3tiw37DhMPCrvdjqwlphHQWtJjRMZdYJAB4vuJGL6h3WoCJXC+Ah
ytShNMnEmJnRhmR+PkxIfjQMHMOoKNK0FlpqUvXMsfxRpPY2gIzkeWDqLfZJqHhqa/DnL8re4CV4
5EC5uyxo4NTtJ6FeKP+oDqE4PJGa54hq/2Egy8hV0wuYaeuW45sRLTsouFz4NzinJH3IUcetc6qJ
xBBpFoyHMVHiK7s7TjQhXiS7BX8pInJJTO3UnoFnOJALuta8oaMUG3lxxsTzRg91gIeDGQz3KSda
v3nlxVr8xWDSZ+NoR3nVpsFIylcAS8okKAQWPLjG6IgDQ2XMoMTCXCJ5g7A3/H2K4hagVknbBsWm
yfdFf2BMxv1522b6ea/8WSN+/z4ZDCbCAI6rVlDv6cUzBgk9/n3VRm3p5ELlMMRuRfiRUElo4fFW
GxfzIjp4rxTlrNh/RbRQD1klYRwmCuuT+IJDJbiueKavo81EBp+zbPYw0bQGfWqyCyHJL1rc1Afj
ir/y2KGsqBCfuM4iJSHxkg3w5BRgMibYZ7waMixg18MamWRYGat0GyBGSzkSfyFBljIBbQEBm1g4
ZE/rnGcrGt795KO7vBE+7fc47E2CENCOiZ+vpulTiN7jzVoIIuaVg0evAFMioQykOyVSnL2a3yy7
AKa9J9FDU5gcg3/hTo2v6ONIPVu0TH+WqG42GjLx97yEfsvQbpT1B2p43lrhnLhUfAVux0wMVQMh
52/s6YbthGX4vFF/AwNXWxPoLhMYfy4Gh75SPMJinhDRTf5RYH74TwItN1o+fVjue0fBDgVBfYQ/
/uBFGMHphkU6FzPWcUcBIKSuRkhqq0jVG1f4LMWjFTD2ARl20i9vDrLT5eHh3ejVd36PZBSSloUz
nHLWi4tHnwLTihAaFLmH5KTah7SHXjgHTua+JG1zA6q1bumfYPnapJI0+BdPE/guQMwRGD6Hdtbu
2xyS9cm/NUe/bZkG4mBU3La+OBfVKkT6ZABl2kVO9N3DycVSv15UbZ8Zfdwxybz23qhte7aZyGzI
v69NuTtYKlceUL/xp5Bv6L5bGCyc18y0Ws81HU0Xmm7mwV8w0rncZcuLTS+yj/WfPgR/rZpo5g/B
arV0yxk4a25gbpBgrYA0JuDtqoTW4777Cxc3I1K6Cr8fSdm1Z7j4QLJxnlfVEK3bmTyAD8qsn27G
sxHR5IpOlKTMQEyf+QG/jdtd5lFveAK/0o1Udo9tXfvRuRBtCASCYgFrsX3+nXc/HE4rpr64/Nzj
Z7I7Z1H632dAE+5D8JgjcQJiTztCf/NoRQkzTcE2lhCVRPyeI0+K1kJrPlM+qgfUTK6kDtxJp26i
qRH2tXVgsL6bo6qKcV0VaMjeJHIV2ZSPnTEbrSR7ToYCj+8P1/zZKHMpcQmsD5Lr2f051R8Fz6De
QQtDMPHV8SmXjEUvHClAdkaxbmM3LyEuWXS3sl59ZVTT4mq0gYGOQAAHnBZyO4A2oyqWoS4R57PK
NAyc6LxHZkpCASM3cR4d1Tj/biUaGG920HgJJt6cksxyZITFf1UUJOEeAi5PQ0PYmdXzNKd8upsi
yS3e3IqNeib58uugLaiOLp2q/EoXVR5e/PFndhpKj3TkpKrsuhg+IddzMaMZfgMwRJdvxVVclxr2
o/IGuhnYNS3x7GKNqYNAwmgW8bWU/YSVVkNRoLaYoIKpE31AxNsT/VdW8Ff3iPmAc/ei/iE9Qxqj
Eb/hBAL/LFREHDxPO64M2kat+xAWtCOzb/4ODb2U3U9/uVTzzjHF7zRy7/xlSRZTHohfRgLW/A3E
sqLFC+j/lrrtR6qvryXszMmZFEPKsiSDUnD/W49ByhudAcGXkGRQlywH89dmA3UCKkp5Jq737sjn
V3waP2jOGkKem9jtC24lmGqEiJHTBWYyr77XOEvFpQYRyzvLr+iXmgVOSkLjKwuZhyNWQ1XN8L1p
SI1kX4UqEVMygXsHGDnKrZ7G2IRNd944NqMMcS04RxN5D6ZZVAZ1AY54n48AYlbHCzKWZcwHQnrm
/e8E74poyr6yb3JhkwTHiYPtI2Xe8u40gdvx8bmfHYK0Do8zHxMlfGkZo1ZsRZ4shDnPQIaB0FXx
ruFagij4FLBihM7pPO8Ei2f6dHS06zbchfNeHRhWMCgX1g52I9mgnQo1Nq74mpvyDsf/Yho11txs
MNXMrA58YPH2KMdJ/+mxMoy+f3YB+7SykkFQLGsw9i3NOQoEtb6OqKzokdI7UmZYAOmVyuyd3bC0
NwVBAuY6qC3+Cd1IZjIlklxLl0GYbot3/530nFDioVoT2Ubv9+T56tZqdSC6Ofo9vD1EsdCuH29W
YuX9F2g/YgOwE0BqZD+snPPVIxTZyAWg1H5zA1CvLFRpS/jRWKBXfMlFn6I3VoozDtXgWp3T/rPv
mIV2RsSwTJlyvHBCXd903IMIUoRbPvtFBVQ+Yd3RBf2b/6XNlHY9ILpBgqw8D5Cblc9ho+jIr70R
N9/xzoAcrLWG/Z+4le2qF3qm75CADD+BMqSfMwBPHI1HCIzi+wCDCyDtBMYej+3Zpz4M0fLiaXSR
lKopDgTGelsWzRia1ImO582CUiAgSKjfAYP3UWnt+aVOhWJcxK4N8Y5U76EnfVHKG14RFEOgQxx9
iNy7gUIomiXJa6VihWuYWJJnhShv/pAA37gsB+8d4trn5Io11M2qjxRxMBwqggHTw/3YGjFrHFom
IzSL7bNI2RHTtX/7d76Yr/e/MVyIvgPRZIbzgpSyTbn/GlSiunZLhZZ1pvBXT++yvUQA2ytNE08y
mD9JKxtpwoAIaZe4bOVtP8Mo2+JqHca23CM4c2XVGrUBBSJ6jGoM82pq8MFxCRyFgz9kbcuP/djY
LkPC8w9pB8puHZu4Za0vuYJANvH7jmDap7vOgANWkqKFVYlTO0WH+SQXyF2Mra+7+i7EMWUtnA6c
rVYz+c1/JyzG5KZkqeQ59ozo8soyK0Dc8u+LTAiHfGYghNEpu3ESJ0iUVeLUE2WjZFkPySFfyEB7
ZAGYRnHnmAHSB7juZUPcpCXJiEYR7N+JIBs2FpHsOMr/YFOUSJI8Slc5f/X2WHNS82z5ZX2kpkAT
PWcSjawiLLUwyeZSkfxnHIuA8JkWlaGSrKYYp2pKdvMziCQH4JICz6hVcXO2XGwlMVi+zxh6QTfA
+MCHtal2YXOwx8b/WLGkba4DySSy5cKBHnYpRiWuYYmUR33J8OKKPtj6mFrIUeWSzOK3RfgQTU+N
+LNsNZJcPiKfqxNpKWz76D8cDuPbIevwI1SXB3TJ7/Wdnb/0+aDhtcqtK4QxXC4ouy/sfnq3OsjC
tga8aZe38PrAwkN4GBl9m7OoqaJ/jK4asPt9pZ7hwywmAWOh/nPeomsZeC3YXvx99OW83XXeq5gA
AteNGhCWAodhVBUGTOFPzJ2VWqzMPaZBHr6tMICNlVmGQeA4qjc5xGnZ5Dg8fqBkozTZqsA90Yi3
Er6D8QJzLzd4ae5kPItqbyobYWCgKk4dztAmT7xqhGx6AbuJ97SFZzN9bxmfkodO8F2aPTvPPkhb
8x4e4BFd/ySIoeV228NHiHirUjecemGjP/2qDHN0hbmaGFRWQHSL/tjSCO+ims1hwDs185fv7lT+
oyH99z3g8+qjqWG3M8NNcEZe5d97guJ9krmjiy05n3JjCga3uwQbSWuoqRXY/xmRbDrob6aymF5l
u2xC6f+3BrC6nbRp34bF7gIsqwi4cSmVHOza0H8nXnjlbtg4grQK/IBbue+d8gsHcIFHU3E6Gwht
v1TXxMT6kdKCfk8pQIJld6Drt94lX+csqslKWvBrWRCmC2C0oCXm9iGGeDmpzSyyppBp6svKkW6X
umkqKVy3xMV2o3eFthLHxZh57HXoI+1QpapbgREsqsMc0MpU7FLKmnXaT/ckt+CmaO18o5LTIomT
9pDI17PVHnRkD2JphVO7tssXpzhDNzTK6kxORKQKw+9akYSUoyT51Vwx8I4K231SdIm5Vvkf1HOy
dfcjULMVkmEKKW2dQl9GNTJrxwFbgZhwWwn9gd3xYvZ/TSPUfhz/QG12QMIv5RPnAWGJpaJQmElR
goQ63T08kGg5i5EG7xr7jPuRBpDbVIkHj0qcxJS3ktg33cbWUA7lrBuiraWrhTRr3F+rIWCuKyXw
jK0fwN6A+vzaHKTWgFANMEb1JpevKBzdmpKSF0x+v+yc0IL8HB43y9rYDOWZac4LnIQ8J9fRpr/Q
0JWF8Y18fU4ffH0BM37n6qLItcomOv8I/J7q4BdDnFT2Mwosg3tTD6S3aj9gNxw7et2i79R5hpuX
7MUX0Ev7mzbJD3CY9AHzFANGVxotggUsAw9GHAqFk9NuD/dV3tkL8J8KrDKbq6q5kwlWE2EV835u
gurFn3CgRaN5lEvzouKqLHqsU8evciTvEkjnLkZ+odNaLHM5Frti8ARys9YCjRzvVlowbHEmLm68
YO2gp3RtXvOfnaA2GxJgx6PMTuv9qvVoQFOCjB5pPMOOR/4goTvdKWEuDq0E/ozZ72Sj4XlwV6Dm
XP00Nl4YkCOYltXuQtn0q3CoWq0NU/oiNjTej0BvChVrvQpqKCN+bur/KBkuU2eav/04EPWNb9+8
PxLjjtg63cpHnv5b0mYzi6uGONNpKx9tXrWfQkkHoQxwZa4axXcTtytm+kC7PCR43V9k427fJdHF
WlFguEJYF/+vE3bgRvW513hv+9HcJd4Xcz5+MEXqGUVuDWTOX4KCJ2KHgamVl1ZoixaxhKfBKswx
PHPW4OOs9sIjHEEi6wGcI29N3T1VTRRlHcrVkqwrb2/sWzMgdGklVophcnWJB2fePWXSCh0CRBba
zzqS2D+U9b45gPtircYb1SVhhvTC9LwTpfHm+8ykG10h6fwiOPviQvkKRpSMCbFu467MSKobrA7f
sQy5HD1m+3A8e1XUKO8RiD0L60UbcjIhumf5KV72yH4jNhHLqnbhwFirNNdD4YMxZ4A5CCnOaGsN
I3VdqdixlWIbgL9vMmvcSieZwCIQBxRPaxnra+b2dsFWpoJ/RoTyectaJHYmqRRKpBXMZcj0BeaU
Ray6sSmpOwYM0uElI+GBeCFFS0oeAC8n20B/0kJHuk6E1q/lG5ZVUO/Pxj+IqiiP3vKQ9HggeXl2
ajMmYl7RkL/S8zXlnlDsMNDNAMjkZX2NWOqIbSJ72AergxWBtcl0NjqLvhA13eXCaQQjpHZZN3Uw
hlcnMugokvnFUtKRV2rO215CeZ0hrxpGCK5x17h8c5MjTat/H3WTqkMB+UFXJTyS536TJIeBsSbQ
FPQTrQdY+T7RHKnezNAeXIkOMvMjnVJDLSWyaUc8Tiba2Cm5nqnunTZ2Fck2P4cUdCUbEZt1r49V
AXcNxbB1FQzZiD4W3e7e2j+6oDup7/gD06nC7/EwAG73l7tC2GPY7BNsR6e1kZ7PagWZ0ZP2YDpF
fyyL+ffJpzkej8NdJpCmSZpOnLjCZbektisOlav8FlHdjpxRC9mog4P0zAXivhuhvI/+NO7XEprH
fhQcXOGVzcrlm/a4EGe1tWWt2ORsaItjK451naNqqVwjj6QyBmnxWnqBnS13aXdP88FxD0V+g8/T
qfXmYBkTeG6vtH/iR9eIZQSX9VF2RaCduC3USxpMqAbubLKaIRucyxRhVFCylrr2+oWVVWA2kQ8v
W0D6j1yMnzyFSZJDt81hWXANwA09Ea+t4672dTf/xElyDBnoO949AUhMfiZjWvhasuyvoiQqg2OI
oFizqjCqTavXZZqtD7axlzy5ql4RYZQMBbE6zgxAk0umMJ2GAk8etScGDhYJGNM7tTey2Z0FiZJs
K+5D03qQ5UNr6M5SQCWSWiT1q/EiPDnLNeHOB3H5FOFjjfLvwDw/UKj0sLSNPB7qTmnaf5axI1Z5
lALbNwz549UURe+MZdaIuSUB9rlI3Hx8Lm3UtzwoFWCbEFfbcr4H8SEyoAy9Kg48LOaL3UIC6ILl
0WReQsqJj4LOn5E8Z7NsDUpAU3mytShKeOgdBf+u+l7M7Zxv7N0HO4FVc170v4JyveVWlp7xiiP9
zoDMOI3xQX/sPWtFOqXV5mJyCmDmTG2//Ar4Af8CHcYBY8kqGzbPfegreyxpTSi24mqyPDa0WFEZ
KOV3cLx3npaYCrDku4XJbTDCJOh1+joW86hMpwuFaiyBsu/71ncAnWU6Y+EYKilUSdT5Q/w9jKD4
A3qZOL78WJuk8AxccRno68ftlB+vQpTQ2+3mlCfoeGi/3a3QWMWd7NOnbobJwZBgl8tlb47X1LrG
cJ655zR7tH+HmaK79ak9VAgDZU2rXLR28yMfNzoMA+c7DPqx8dm4+WvO9R6nVNBlXXjV/KVAoOUC
YebMqLDl9NOjd57y1u4LoBoicRKHWYc2RUaoKkkJZ6M3kMeTWhn2UVmUXiFTdIvCOgreH+fujEI6
v43M3zgA93vY1CtQsbf+TKwP8tGITqrKBl00djdDU3hm5xbks2iEzgF+tB9YUvSOnVkfw4RtFcHb
gqqbwhtkCoh7CIT6WNMuxCnYwCldEgZhp0A3flX/mK/SdwK2ddQJNwqC5jH1CeQrBMlmO1g1HwXM
ABl7uK7HIFsCWUTgoCTb+HvWB2JeG8606wpT1FnfK6rtrGgn4f1899RqACQv/5VbTSe//yK4ySjK
AU3yfbO2QbVbn7tJprGre+fTYUcCscxZCSC9UkWkVrj/KsfO/9InCf8ubF0V0Md2kB+dQAZiYhbT
uocSvAa5j6mlgovRz1/vgEw5WdsKMfByf1lTvEZ31g297abMcmE9pCJtsPGLIOpe/izDMjBlnuTf
+1vNkil3+sFbomWWnATrRFPbMiD5fYTPIyzEPAkKK/OBJ0aO46jkiibwuiC5aT0whroeI5h7PJvN
iaEbR5DIeVHupU6B4XTCRDK5hz9bqRLBS6DxoUUu5MVBllP4PZboaOvK0PsFf8c6be/c7uGEvMGN
xYJM9alqmKCMkGM3wZmGjMVnNv2Jvp+I3b4uI54/YneG7NSq8+gearkogDJgoM/sNUSaYJPcVrD2
gEmn3k6mZf1PnP8XDuZFDsaph3zpwrOrm20PiyRpQ37H5/GF8ED6UWAPzQzjjphTx9HjRC4xLIP+
dMk3FnAP3XlaqJQvNAoghWwDSQiBvf2cy4+tU2RwEKJyGc50piT+X/0KXYX1pZtWz+kgziOxYxcF
rkJ5Hhzhu1JInq+TlXqLRL9X2Hfzsvved+In29rhG/2x+HvJ6/EEPDYg8bsT3vb/SepWQJML0x8D
kA9HN4DnWI4D18yfVpi0GV7vH2AMmu/lH68Zk+Xlwosd9SPRRR5AYtiqomfWB6WFTO8uwKl7CBv+
+BwM8+VafIfYWEijAFImnDmLWTA6BxdMrBB5ANazbnYQuQbJkOdXe1fbk1Z+9rJk9Fzk+fQgIdZ+
eEruSA+4/+Z/oQx4N/4cqEav5iiyBjUnjlvE26ZyGz27RRdxyj7EMf3FgEGDsbVg
OBuyE3M=
`protect end_protected
