`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mgu/yCR4BivO1YmqpXI2DBUSB7zOLqZqlFoCZyrh++VdpFQVFEx5sH2PQp2y7LVNJP7kjhk1e4Niv2hokhZyyA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QUaqpFOIuIG55L0GPkVfb4Zz7ms+/dupcSlF1cRvuBDACG1bswnxiXi9FbDneQBE0pShtQaDbiNgCqi7L8xiLpC0f3+pDg0Nb3caHMRdVtQbOI4a21oBM99GaHMpfUvE5y0zUc2TGcZdGhrSjAdUcTSr4q63qap6YdJgbeyYPM8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
2McPJAxNfiac5OGiRfyszF0d458b7V/2zctH3POJ2XRR5coll3Wsc9wp7DTaRY71bA4EYS4/CkpFITmqMtTFs8OjL+VQbOFZDvwYZnXza8pZnObuDj1bpn4e8U4H//fmNG31/SUKVGdbZbBJShrheBo/YDYbpAlPRLbN3b+kBHzptK73mxfIRxiA4+QnwM/a2VN7053/VVpYoZ8wy6Z4oGj/aL1eDnP7BE+kRtwmAMxJV4dF2mlYwXLMzuA6i6PicWLDgnKNw/JUPPwZQaWMHLEI+nmuOMyE0UKRbaGdXNjTJQ8BHDIM4TPmxVilrmzin3/uKa7QNQ3Swv3erXdwcg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q1aCDOTfsKgSZ5Ix1zR22GTkTU7ql/UJTMoKq4Yg2N2nETGhJ6VwxittTnJF05OLBF+v9q7TlnMIzoSc4XXYRGjWULSReQCGFFAhMbc5Y6Hbe/FZfo8c9dSm37Wmr6H/wrYRpRfcql/C1cUEMBPSbtE1gKR2pV/R8qHAnJVDups=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nhNkgfiC63M7c/ZpbB5tXIgVPqx5mGzNipbdekNVMkyaWPGYm8bbUwJcQ337tp8KxYl2HKrp7mX7QSzphiae10yq1KY00tIei+hAvTzVuiKDYhDEQTafY6fFSk2/PVP7NBJo19PJYTQFxwobjy1cphaNV6/X3prO58HNsBFmeJZCFsIGiLE+p5Zdq9gT2dXZKAborBE4ivHKEm3K07rbMbR/WhBUA6FAK6sHm20PVZM06t8tV0YIMZPLboD38s6JqUBEcUHL1HH3Pg/aRXxoOofTmJl0FSOj1v7VY3S3UWyK2eubTZiEdsYk0V0dVQWxde0UO9Es1oattbY8I6MRYg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14125)
`protect data_block
CIBM3nE68rzAW3ago85dy2QnnvzhEHHK3DeN0lesXebpKWJ6yd/MMwOH7STx3KrDJzY85X9CI41V
QU/dVIVD2IcL5C0MzqXnFz03DqnfeI7wjJFJlMDfF0kQrrXbrOHqui78hfYf7duz+gitOQLtgHVz
XrUN7WWLXbNhxHtm5QwlvZmtCZZ6Fzezo7e2/EiaI+iT8T7Xbuih/XuGoDku7JGP32FutkLxLtwf
Lq/v+TwW4ndHNGOmmCcesP7KQZwCDRXlCgWwrxVXhDfIV3Ehgin+ipdy9yLsI3bxJuEIi9n+88e0
B97cJdID2icQG8PoNNiIQ2Ae+WG5Lm83MHwR/Hstd9bLWgvcy9Pa5GuVwFqaybZuMp2z9c8OLC/i
lbI9UdiMF4WWg/sy14rQpA2BcY3FI6nSQ96ldyIqna3LfppxRANpId7Jeh4He7CO7MTEcA7c1x+6
QG2NbboIgZcOuSu3BOjk5ZFgVKbNicOiZkZLkcM9Fxe72jMLt1cyQ+lNhQewpVKggS2RK1pFWh6w
ZQgSasfhD6yioX5jLLVpo3B8gp5SokAbTOaW24rZse1R24ZNejRVGeG0fU8n86e4O1y2Ed8l6Zzs
nSx2tiwqQlzeBkdX8IVE7hTcgOcknipGrrBB3QisTkQgTg0UK6aknKZ3MSM5ehqA+4eH/A0Haz6Q
I3SNTzwmaK0G/BzXzWJD/5LbD44YYyfDHwtTou7ymqdwkfud31JCRUUE1Wm0a/lznOiddmC310Bp
EKkYLLKFXkkRLn5l4/TA5Hihg3TnK+43P9QPKdlmnH/DvH0gldvY15RII74DKIHeiyCPtvcGkR4a
m1WI+A93yfu2rDzUWb3LzvHbG2KjjyabxFyclTpd3KWqIzorUKZwgxn7BY1y0oZ09JiBW/QpDYhC
nAD6uR3xiqzhiL4XfwjZvoq3Ps+H0bnP2E1RmjNU09iIadYv3y5MHI3CxmlZsiMJ/qoUnPoZwl7k
6U5Wk3xlmw7YpQ2mhy7bjQecGWFmI0Dj/jrRfUJ/mMlEFCgFaX8Ulke2MkGCMj5vKYQRSxlgl4yk
+AianarDSnaGXvaikuK5zYoppIX4BLhpn0doreHtIjpsRi7NTYVZoM2mukEr2GSbdT7PCufEmFBF
6XSzVvuRILGR/CqounvIxguHAK1b6fOoO9U7fXcOy4a38EaBurM6cqt6BFaJTwov5thh+jW83EUe
qzHDvgA4qcyVxFL/WJosgtUMl3kYrcWokQ4fXyPhsWTUDqTI/YY3pCScBHEbVmMsb/tKr0grT1UG
/LhJAD8s2Z/p76UH5ono1mXwYPdD9r0SGp0D5H8GPCakoxYLO9gGqbeaIG9Bwrs3J7TLlKJgVcWm
zF6W/sIWT0ZVC3XoqtVYxYdynmXPdboMhucekS0VjGe2nZPKQrrrCGLjIQfKTtvExryA3mwbczzs
ECkGehlEQHtOmPNescEvvPNfGQ5Y5/jmDVTEE4MnEKTLODkPvqGYxSQIB7QgIOoodVrWGi6fI/KD
2ep7oC31Djnp0Us96n5pelth+QhotJdHqeAusUdu2aFihUftuXP6SfUWhMQ/1MzwsLozhqkS7gVB
t2QhHA7Ud7Y3WVt9OkCkwak1uqruraToeB1TK6F+Z5k9mad1i+WZHblFDPtaSY36x5BZG2IOX3Tm
zEcb85y/hEMPqw5L5dm1jYO7O8M6WWRWkJ/1E3GEIdJj0UukyFMbwvie62/RS/aMUn816Sfg6Y9u
OjThU+ikpr0Uj404JZuDc1rR2pbqNGQ7theLCOupU+lmYdpkTXfsLIRCZvYX/pdnU8f8zbwGL88H
42JTp4txeI7jvGvUsbxiO5qanoes9JnXPa3CN2VbnzMSAoOj3qRro4CKRbJQJB9U5N77iN2NNz5T
ShceuPSAVrTHqLFsuFLzVtws+ZMQFT4gJenrJ7n3cnTlLsID8uql9jDpQP3VdEVJQs/pA4aW2y6A
BIh4eVisYJvW9Zrzzq7xePm8vWQt6i4pPTXa6Bp1xpDVq51Uby9N2a2/vg5lX5FPEO0tIWRsPD00
8aGbJGa5axX2BHqgzXWssZ3WScASh6kx0mc+O6tSO/+zv5w/HMu096vESzIJ9cmraHIIAf998ECB
QjRzNyux46yp9E6LSlWfr/XLqE8fxBjPC8wjBM8r7KfBddXL+MdrkODxrZAxcWBFvNG5Icku7Nqz
sL6r27qX+aMFRFG3/854hq5aYlPEwfNdSQ2VyDJuuMbyEbsZ5cT3U3Gv/FkjqQ4oeiJsQ2eo/hlX
6QXRaA43vO6Qc0xrMauZzyxtnLEisPOXkAkTayMgUz7RNeE5gCQ69hX+/fRlx9VqQwAmD/rrmoUP
0jTkSboGsxeOXoLshMg4ZPRH8bptBF8/FIta68A6i+qaG7iHbjO5H/XAD8vidY+P79adQgcS0bmE
BsW2Eg4e99Wxi7Mbe0p65KLT9c1NRlYqzH5tsp/xePjMxuKVZtza5XaaqrL7LEERkmK2H1fAcz0I
+dmrid6Lq0HpsxK5HnVP3T9Wu8w1PMMxtKTz5IO632SrS9E+oni1R+wS+uerVZoMCwH1/3wwRSob
irAt8eBZPUPovT+s2XdAY6iAJZ0h9J2iClTJ7A/dZbkW7To5iBgSVm9vqhrnIO3jacMLSwTxrJ8l
JP8yowfd5xR5HbmEzjvqI7m9vlzNpkxHW2YWDaX7FjcdwDiUMiiVRTCs6QEI7ws7jivyy+MGNXDh
vEbXDCKHoxjHCI/CC6MzQH8uZh8HyUpZjpSetsZw04vzFeXHs+7u/LzlmBqlvg23YsjL5K2lgjS2
qyVABEEw1DsX+seia/IbsDMoYIUeYiKV8q3TJDJ5Zt37sxxZqdRSOOu7nYzQcUeGSVcXrqCwdA+S
jDB6zN4yq2KUI/smJnIm3dN3mg4XGpEV0Y8p0vXJ9psjwTLCiTXUyj6H9OnGniPXUbPwEajkRIrY
23gKuUfkeHxt13aGcK7jOG8eY+1bDSZCvTxdJ1qxqUeZrDstfE2e1t+JGzCZGm7EzF90DKsT8AkF
7FOtcOodjLufoczk/71owvaVR638YiXXB88rgISmeXTVOHMfoM5hW6QbajUNHYZr1w7vck0UJL4n
wbYnP5kr1Y5r56+R1Rirq09Y8xf4d/ZogxNu6PtuBBsPICmdIBH8gjAL11qX16LhkfviPUgzYudq
R0rbsJeTcQoMrBtr7D3wCyks0oP8x/QHJCUKnEPANzLyqxH3krkUg0QYl+LRZj+/bWjvRCrLjOb9
+6GtQaY+giNZTrnMUxEddW91TKdxWTuKObqCwdvf1/YKqLlaG95HVYYcxhESnin7vzMJAvoEIwg3
PV0AnSfa7+E+TgtMfdYaAE4FSWLkFKRiM+zqLCiIFWpacYEVc48pJF2C973z5CuhUq1GlA/xKhJF
OhI9Eg4GvSifLcitO3ZSn85b3TaPh8TkrjWBwh9hPSIUFfhVn0Ol0uhAXDS33LR4IdStGvJjbW9P
65WtLrxnYM7jea7S6nf/EGEo3O2qb9Cop7qLHSm5GHTwIQO1gBLvgrZTPqnpoE0TS+ReNJHbYxQh
TF7bMcx617oAYtdbrtUe9aAYKhoiSXDiz3UTAEee8mX5eKfNZkzG4HGNVvGF+y/8x7A9mfXTACpw
pHaSJdE2VuxkA7wgHygmzqHlkIkj7Jcnn+nUWkTJ2200SNPw4zAW0Mj5UxKsSBOw9yqTFVcM3YSg
deSuokifrartMpvVFrIkZGWIIDEUQMVnfmO0gSbqTuaWa7qTUa5dAE0nLIrmLak5sJHzzJE+N1y9
lNSCeebIItNgs/m8n+tzKD6JbL9aJ7rSpH4EIEe+Y1zqh/asCoJREHRrAstLYaHxMVzCRzF8UwEn
lNry32+GzFPuYTJ7Mu7IWjnsTR8QPO6GosFDdRf8hccc4ivg2+pXTarBYHHf4Yc1IDKRWgb9RASM
5yWwYP8VcjIU558pTnMAk3k2+Xczbxy8220NlWbgauT7sVqFM6K4zY3+dSdAALyJt0fuHdaT+0oV
AiSXETl5k9G5+5QD4dzEgNwFfuUUEVCUgev9tYf+tEJzVwgljuhF1dn/8YZDJIg79azetrLVKYat
bErgn7Bn1cKMg5c2yF3ry0/9l8J5tAToluT1T3+2ZDY3IlFoa0InsxD1Xrzwbb2BY1ReXC3lMR4U
ujOz4ipL/LQvkCq6LH+/IG35WdT2uFSfu7pFjEdPFA7/PznnaUggKgA2ROGJjejes9/IzVGHX8WB
G9vfsLWrKuTT5PHpXT0nInqvWGUl3rv8az6n5quSk5zvzoDjRedXsKSnekMxVw9fULlA5yl3zEw1
SdeVn+eQhZ8PGEFQsjTePXg67EAsHIyMv8fvktcSvEtd4DICPwatbn1F15HWRpLQM/0/DR2hVIJ8
SPntCqtVhojnLT5nhx6sxtNFtnANMFrCJlSxTaL6A7u9DxEnviFCdzj2T8+u143dnbB/OJ7N/d/P
c+YW0N0kKthTaORdtlmD4elGvQmNyK6jvK12VtQoa9GCaDOVs/ZAqQqxqT/B8eZu6TwEGJx90FQs
LT7rqdPkNDIe9+RHc9U5BZA4MmHpkE4q8naP3b0qAthg1W5T1oLN72LTcmS7ABORKlOplWGIZiC6
TwUQKYO07CIvEbXsD/TbBXXQVYrtPz0ow79y3gsCLSK8MevvL4m7FduCWeaXnig7Y5SrINzY8qzi
DhmZpX09Z5Doleu20T7r9G3TYjZHN8csfQfO+I41Z8DudNcxqdc+L8Yd6mS1dAvTvzYtoUyKBSOF
OlKg7+Gq7Asmowd48McDSrXNCCUlNw6wDkXcv5N0nW3tVF4MA//hr9hvu4SsdI/y/RtGPvmnrpJN
2ECQCi3Ix0QMwqf9vewGUk18HSat0y38TTG/7ARQQf7cPn/8ykNTORptqQOlredPpb6ak0uVMH8o
vjsFbTvr3uiUu3a8O5r9tiDJs6uPNxb58zF8pHDfZvCfhZH+uGkxK4HwE9miSLq3K5hJUFoWhILr
9df8Oh7x+taIPS2gSigwsh2zQQwDFAITjhw0pr+DuAlxRE/WMCjfv2BZ9lZT/TsPtn8OcNOjyWML
iVzZ4YM9q0kj+FnzfB3HjLvEpxRGIqVacQHK87Q3tIkZtbs8V7LIQKBn32jzi/MYqnQYcYjFhYWj
GiOC2+El6wsJZaPZKOhbXMsTy6vAyjlTI9alaGR+WUdCuaizdlM5dAmRUAY32wwly4wbk/apchRg
nYQB6V3lIKEUU9vYJpcB2CbWcQbZvedSassPndVtm0SZaCwbZUpaXlKlxnJLVMcr8JwHiWIIWu0w
4McbQtmXVOM8WP65XSbPTeH+KnUEVjv8wfY7gxTFGuo/OsyiKNhT94u0JEmvQQHwDpmpmqJn9i8C
305hUpGhAtoNd6yGl5MvmpmxdXkNGrbyI7YboHBuF2Y3LrEWVsqYyzpt3q7zKLkg9GagYcAvl/ZV
yZy5Tnrc6jvNfCpAHXE34EYFcknHwIP7WZz2gnbmMKAU8gXalVTp9inTRqoZhfhBTGnZlj2d4OKG
OAhEVBEeZbWVTbMb6PG8XM2Lal4tpxkiu9kLhG/cKO0TBzDJq29VJHkdr9iT+CurI2c+6o7mGAC1
l6mXBM01Q1AqZ4CCCNSr1ERQViheglsEvPRJZnPJZGAu2dzQ6xihiJfr6Gv0D4NL+u68ctXr5cF5
KWPpQWDhceuOVJx8FzVMbraNpa9+U39Ti+3xIDoKUVLeJ5ufylzClw86IGFPoB43YynbNzJUTihe
EgCRBx24Zwa+5SB42fByiccGpNenllaFcPzZOnI5/MAsrj5FeWu3VUFv3xC+qfwt2A2SJA/RRE+W
Ae5HsI3ZQ9UGxz24sXhHB9g9JwxAmU9rl2Ujf3JU5hK2SQtQDthJh7PihMb7EZk6R5zOZBvl+q2z
f9PnT5AhQeOWbFEFWlro6mn++HGNdZ9RWsiahyLtKpXrmLqGVYxI82XQSRGJgBUrHcQiuPamQjxP
HuXcq2KvJt9Qy+/IUoKF/EnMDjkhD4BrT+EfHuQisfBOxUjvMNiw/Nu2nsW+kFoLpsGny9snzBFE
Lxgev7+JwbK8n+YdAKa3dvy8h/5CaStNBuNC/UsuLpMRbVMWvSTJjwLxEvmALsSKATPtOFQpBWVV
ft8pDiYF/AM5/ZdExVS+TFtSoCXd+rtrernX9sqIjxtxNonZx91l/UIQK0WCnTU4EM1fANIGTFoZ
SUjZk6w+0/khUQALsyRjjdvityeKZWZi278bu3BpzaIJays9yMee604CWOFMqLF25kLXwsd/vkaC
qbG8UuOKQksP61T5QcrijuOkP55RtWcUhhCXiWiXf8KjgCHLUFwGzSGyV7OM+BHhWWPD72CVB/Lp
18+yUCSfMojpI497u6NGA8QXeBM1PbdK/m1VAQ42RrSo6loOH7blaTcP2znXAITZ+Ohg3rYxoMrn
JZ/xl+lueKuws504TgXhloda+svYWjBYTX+e/A+0PxijcJWxhs75AAS3u8RJjOaMOw8JGjmZviCn
mohaRdQb23k+NWVu2k8xcy0DuZQioZdnr1r941MXLvpsGp6wLDDS+Cn4xJHsTQgYwXrNtGwTTN99
3X/pMjXxQhke2Pw0LMG2ctea2+ie4rTHrCuTgXFfkA5xrquzAdlNjQc17E2aWeDrRWtxP1d6wUOk
LRJJjAPxzH5e1AONXfKIIGkf3WMmPOgk2JZzZBjtrRyYfmUPPvIP8/QRUzP0CFAPEYJMxo2/bxBB
b59FdUKSTRkBcrIgvwQA69FLxfnoR9nLHx6hlBNHi0ZNeRcJzZdHkmVLqoylWlJnPb333F1wgSsT
bhX/KZYkNnTG9E2cTvFM877lWudQqLKM5WLe3olUjkzU/+XpvL/FCs5C8eStVVGoJQrrvoLUDjRK
/aaLvlYluqJ4/V0PNd+HExWHrAYp2sNqv5PDSiBkl2f6iFJ7TaAYriGKzNLxdZAWB1yPF+aZQHz8
tAwz2toEeXZvL5+uFdUwglZH822RLEGx2FqCOXVYoqvUKI3wQrGqHs1tJg6S2hTU/WtxSVnvZc+B
96bxmL7ia7hyxezQT7BbqFXL0NGQw5HrA9WzZCfuss9s/HEgtnuryz7h2BUhalzKalcUeXmuI6cJ
6U1IL6N5AfGR3x2cpxCd8FaPTreCEPCslgjb7JW8ktjd25Asc3nCF1XtNafuum9tbTxhTphrkiTE
HKTxg6grA3XmGTyGqQ6Ai+Q7xnZlTDJwJijDX3c4OqjLr6kSRWLeOKNwfn+D4y3Lsb1VxSS/24nG
RoCgaXqL7DrKCXWFJG2c2/IiAF++sTUZiGNlUaQAnCOJRfzVKPjHbkCLoRtVW8jEU2iIwOj+8G3Z
TgtqkZsbflOl1k8xP1yOCod9WsznEg2gUFoxLkoZk6L5Fp1gOKX/hGJ/wUpdoaqAIfdQaIAghHz2
Fsl8s4GNqP1pl6BRAt5Jdwb6jDz+NKQq33H2MGNSzEKz4mzTjHHZa8LNlP6rHurIp3vub4XZO0sS
fau5YLYp5eFZOj9iRBGbWJeGrHQ4jo6RsQnwYpS6f5QWCJGTgvTjhD8BMEe9fMjohHKDt9aNJ34+
oodkjjhf4ulspYg9KO9txeZ6GPB10QCWDMagX2+TW3iLPayg3J45FWXM9CgYzxcDZ/ZO32FDgxjm
I4fyAma3ACvWyRsnUYMKlq3+TWLTTTF1xq5/jDJDyDsdss+Qd4tvuLlwosV7texSKEsjDdWQlkev
D1Qg4sCU0P1Pg/eu7NGbJK7LXEbX0DbZjk0wY7vpG7rcrphv6RAQaIdNc2RZV2g9Tt9xLDOFpDtT
uT1ZnOqvW4yB6yR0MUESyw7oJRh/I7R1IslbtbaYMbfKM4L+/qRDTgdODOLPfR1BJQ1AeuE72vh3
+u+Qfg4BLNtw4TADDN8OO9QbiNDdnb/+XRDRzpr2XI17FvAA7xToJWU4/miEwTWOdWiiSP4CuOCB
8SeznEeztxBWFXYsyBcPqceY63RT7vs5Hn+BOZLzdfH7ZiatziC1Y2EqgXJPDDY8W16hlDrveGEQ
SQImvV1bv5Tg4NY/VSuNvvkgxzOLdnYgCUkH3BvHTICObJrlmSWdQBMumPvc99kxb+AKA5McMpKJ
4mloWrx+Ev2ZSk3L7TtMb3rH/q0gzLnMiNxqEAclbg9BVRPA/FVoN3a5tee5eieLvAoMRYlqBl3D
wXS5eiuOAAN7OSVC5N02hSp+CIW4pr08l60vFoM8aSZEhbZzy+wmWxxpx2ZsvoHjcdLHiIKCluXR
f88UqIzySy4P2glhcqnrEy0mU49qtk1DTFABMzyJo9iO5TcNd8HQQj3H5jMQjhUPHfUxQIrqHN9B
P9c2mrNmKSx/xSrL9tXuLgxgLYLiGROPUJFcWioXuMC8wDWs3htZwSJF/MfxSJZaGefqAcniaq3W
5tUnuPXDZLClLKgs+SWkfSSsrRGB0T7X2goPGS+iei30gr6FQeRwLho9QjoUwsF2Gkte6hAMYNhT
bo82MVvVPc3xNeEjvQMhlbhewLRDOPaBSCXGQFJe8pGVIq3Zx8btetE9bH1f1arZcIVOe2Zvv8cN
xUFXZVM93d6s3u9Lkd6wzuu5ORxUZIrQt5f0gZqn1dooG5xNNm/47mSuQEiKs7jcWtV2cI+u3oUT
qoz0wn1r1ekUB89HVIn6iCWCRxf+QuPgj9HvdiYNnXYfK+ocvDwAqeKeeVjiSB8EjFjK3Jbqllcj
U5KPYcnVe47PebbvveZkcZFW/kRPfqub5rWaP3B+9b07pVf2oOGlGKaqmMLswk+AOFJ3T2dt/PQZ
krtTl8JuIfbHskx+3Q48tu6DsndcvPAzFgK6Gj96Z8SbpWvck1pydK4P22DPoyRoTlSj909Rn59Q
J41w9LISY9PNxJ7CV5PY7HAHkiGegJKRUgqvr/1xQHUBOkV5CsdOtfqeAW3lXZ80SgMuiAcaFh95
FTe5kOwV7xnWgK9+MI4tuZzEvKNrURawvM/BujkD2ePe6Sq0hFBRHEGIwufnb24qa/kLm3/x4EzI
/z7n0cJmDwxSfYFHsVUoMmAs0KPVXy7i7f6bh+8Ht4Od89idf7Xpp+dM/8jmozzlPOD8Q81Nzb2d
yvNp+Fr3A0Y6046pDiADwaw6SE29HERt39xi9iaHfKjDJ3qa10ljfCAwN8GOLDp6ESfw91lqzBSZ
g9zrPshrIqV2r6YWmlp3ATM4TtNtiOaUFfVuBNzE4EQG91GYrI1oFiQEDfPiHqxrLfuX2jt8BoEb
sd4AyfKuMAfMSofLNNl6SDRWuLmTmlb1B3slMD2ww6/GPxyGaxRfLEZd0dw9a/PSI0GJ58DhhoUd
TTV0+2lUmw+OOoQeb35hzdkczKnPiW3wOShmW3jWkTpqAJHk0Kka8rzA8B1UdzzphYCMIozInVRr
U/ER+Em/++145HUOEGMsbsvZZo3+5ZAI/nJo1DLO1NoO0/7mFypfyJyKZ6M1HCnsjJIxs5IZFkNH
0QXi7ERlznXzhKUNKYJUGRFQjBw9ADLyfuF3s5YQ6gp3/fh6g1KmLOQKl+lLrYch2GSbo1Z6hPWb
EdsnTod/IcaNDw1QTE0xDifxLVGnwycAX4Ve+1OLz7sVNoEd9WqfLVys827nc3c1cyPO4iSQbWLZ
sfRvoFEkX+IimEmgJaa9QApU3a46v0sJZ6UortuiM9+0TCh9YxR8W6odictwx38PlQK3L56SElCE
Xd5vPFzv5HoVYGyA48BrIQZR6gUHKGRdBw4i9Y5BWzqOamyE40F2u1HmOB1EvAR1e7YKz67qXw9e
SGZPQjsjVaMclOpUFD4oKXth44wh366Vc3nn31tys8njJC5vkpcW2mpBTHMi9BLPq0zQjYVLcBCG
daFWz0YHNor9gkseqfcOGLUiQkS26ksfEihSPPMBfDjzyb9KxjHS4L8XHizcU0mQ7VKyNq9aklKs
wg2/Efk3M4BejIylgdR0ZVgz5PGH2yCLiJXpYxwNdUq+7I8YDvNus/fEdzKs87yVbxTpWrJR/Ayy
6k9mAlof6IcnvpZIylcVbYKEu8a7Gtr+EL2+ewUQYYftZfMaCxTtJX8rVjTUCPV7LnMTUdIWHR62
G84Ck5ckM/dXGeATMn8ai8T9ac80xkspMWoVB2foehv1qMM996qYnymztpBEVBgu2yWaX5SbCwHC
tCpLfNvDjlkH31KH6oNqk3PBH1LxS1Bn4p+AhiqDMBj4yVGy1LcOoJ98x4MIxipo6pDRO9OTpufD
JE/emlnMKehq1EulyyU2ZAOZoG9nd5z9mhJQbVagooiLKc4Nm6pnynlghHk8sDAC68bFaeh5tZMC
t5Xk/QxealivkrqMlWvOvcqNdRdh3S2IM34gUjuYaMQKes1j5sYozi4aFJRhDakRiV8SrCwnlKn5
1Bh09SVkqr/FIEpNR/q98PKetfonSzjmaP14xhckPDGo0QG1yLOxo+eqH0RJ6QcXMF/JgUtxofKr
i2aaHFaOhmZLVRGx4P3DockMQKN4nnDLlUmzuTFG9oARkYCpClYYYzU5qLTdPjnHgq/SdNsN9quZ
vDJyTwFSxKFmNIZmsSRuHvgJaLtDy6qEZp9ExSHhSlxxZFoJu3I3lsWp4vNCVC9OMmdxDiS0AxY8
96Nh0ra8MeE3Ihc67Jszybqj6nlHWf1gjyXWHn866aFxgr1jjrz4A/ysUu44iw5SglAG5iAKq40J
oVECIo4N5GmrzJkRYvzm4cAMp7sS7w/nifkBjjZspRxspjKHv4Vp1Y040VEWatF/hA8+HFdkSiid
2GWox1bK3nnG0CY1GPvgZGP5Lk7iff8depqncO3spDHAqMatgIMqltDDX1ForMVFYpUwnlkPxGUZ
DJr+zJ4Kt1/LBuj/t7autFB9uBPBqj62TKE9CeGekGVUHserFoFhJj/Ns/j3RaMTD4P2Jxif3JLn
Fvbhp71WEcVnlcBOcs1MOVt9tnVcXIzhYtvI1irzkSC3Vq0wMf2VVXqPTDUC5IbuRGVBGBSkeRwq
upKqc31FlDfbxiN2D20QumBkTHamqzhlGDdGEqwkGVCyBw281LRLQMQb2nmbygkfXcmN/QF4f2DK
wqQHDSvm3QhxVkotKDi2WZQsyruVd7Y4yI+F/OYZB+vc4yE9AE9W52izGDxUKqk70MQIspInD7pz
w3X60ET5a4Cmsq1DhldrLVfQqQpXM3leyE1rMtDJU4X14mVmd/OJhsYRwd9/FjuyyKJFcw+Wc8JU
UzFTWjDN5P82FbgfgtQfJoGLH1zqEvHQRUzMpg90rsJdoVClRKXwSf4C6S9iCSrKptetwhFHFweb
MCIW8ivCujbQkRH9ZeZ+ijDQYGBLBV6PFzGcLjpPKli6WNIje09civLCCvFVL9/gUzdAKIw2n6bL
J4ti/Rg6IgE2YEklRcEHD7JExCgD5i61m+LD8dAFwUjmkfYiM5464BVNy5yCP/7ZjjqNq/5B8+ox
VxoOAlmxKt4bc6TeiX4GUcAphI/WUnXhZoCIIqAhTt8bC3qefnZXL0Bym5EvlyU3tnG89C7r++QQ
7aZUCXjbPFyDB0vnVigPaFJJHv3elcdT8a1GcLHc7F13m1u7iCqwGntkZudGaPbk2LXvLMu8X578
VTMmfCSRP6JzKsUK0pJl32rX8k8dhuQAPyvxU1gwR5VXf+1aDpJDqytalZs1fbjavsA1KpCtWKnz
phr+vBDrVV7bQk9MoP3bTi0X5GLGOMKUACyoH8fIBUWrbqeOng+dcuIJuAwVtzGCKlfmEebR5jh6
fUi39FOh3LBQucAjDyBMRNO4sGeOMWY2D2nzJSJSfnkOJloV0SSBLvcWX+VSKDoT23rQyJOeXzqV
fMdH4+L0dqwpuCNLF4ke0tvPP+pAaRcUv6JugJZ85csbpiV6G7Aaw6occVkP01IiQ/Ksjo7GhK83
wvUIiBpRxM0HpivQ+n9WLk7IONIwn/UdzQEKEd4VvkapGBu33vo7aFe/m1mvrxK7+xIPUvVt3su0
9w/q7IPMpve9Ue+hgRnNr+YeNU4rAf5OOeYCTS/dZBohzxaB/aE76wBRO7EBVfmerEi51yEE6tMr
XFXAGaAILZNv6KoOF1eEVG8DlQVaCm9T9JzFxxlXS6S4G8Bc7a041KtBs7FOyOVIeACWuoqRwpy4
6d43/NVZkSKPeC+PzNQ3hAtppFO/plY6P4v+R0iF62PITyz0SQLI7DaqI1VydGtlAy3AJvdNHe57
H4Hg7wmmu1HPpnRnSVYiQ3bi+v4ZJOLNQ+do2aEDjSdW1luHDkA6j71CViHPzgfIzJXxxwTgQEO5
9/QL+XOseYaih4lC4GkIoCbAtbGn7vtIaQr1z0EDSLquoStu2b8CWLJfVAEnuiKUKzZM05VqJUhf
fV0/t1/N7JV/CPruKXmJWZr2bKge1Qp7M0XpWGqGEFnWc1yeuLX7xnOgf9DtpG2j0jTLXB7YXRGh
NEBpYEnKw6u+3OqvOcfPdQAPnpgCA6dPfHd6sUVwyzI3XGP3ZJcLhrPLtEGn6/raHlz9/yNPjy3t
w6roKN5yYnUb1yOab3YJfvXGa3Ru66UrqnOX/SDRrYwSnGQKQzbUrAUWj8/n2jxP6QYlFr1h3zXp
Vu0KnDCDjVPRYzFjzMEOpKG7RAwsh1xaDRrN9lKiEGWvqRUc/GqsNFlSRnkM2o8reWVL+1qJdRn1
dVTNxX4A1v1Y//SL//QAbnMUz2wdAqUkua2N2PaTIlxhQig2VAnysFV5LUe4jOktrhvw7UIJ3mgX
t5aLb0o8FwRsow/qqk7WmR6LNFAVjUxL7eCPeWa6toh5jjOuBBNuA5wok5Ly+g0bCeju4IKpwDRI
tAS18Lb4eDYdkr7WqmTJZPqJf3q8kShrPR3PNzKuNS6qT0OHHHRdYzwUPCf/RJ0v92glnvBTGEWt
aUXSy5wi5Qu+GFNEmK0wh+Qg0TcLnGBFeN92HtG4aQqqu1SJLQPViLH9A5OJ5XtnmCuDng4vN1fr
TOxJ7FYsNIHVXmCW1EssDnBm2gY1ibMwaoCkcQtelpsUFLuVAurDkcTn4499nlpTyR2TrP5tKdqM
4kF/vSBKECUnV42BVa4SIbPk8R8BkV/tZG9VV/mA33/MCB53GK46OSBt0/xgua44q2HMezvG2bZH
XAG2WrULWXdA5wLbHYZwyL2zfDMdptrGMvbktEu+5viuyjE+z0lbVbo6PLbOJSLtJ6FcMHfe8ZCt
d9JuPFkft2fvggfJuwFQHuAwQSlvPJylI/Wo/ZRBI9D2nJ60QQNYkSYtmPYlOXXWy+kEYkyooKIt
+8m6rl+i0V9AATvYqf0w5xtzpBr8wymGWFQwLDbhnDXtIsZgjfjVgIoMmisTLYCusvFOMl2E7jMQ
t3Z5PTQlP12omY797LRVqXzh82RrBsyiZHq/ExLieAG+R/PeKT1vxdhovaAN/dujzTPuh72hp+4e
CEQUeucbszFZQYtJP7+wVWAp5HWkEWR0SY/XFxv78AK87UXo23GE2bCKABUpdMFR2vk2uPplGeB1
olYrIkTWBP5LjeOn4awP4yjaITxxQRgyROm0IDs2tyQ/C2j8sxVjjtaCADV0J8i9R0584lgzfGkq
HwV44HY5uw2elZ26ygFUBWSkMJOJjt02sJLyR/Dr0fzgq+CEESgOtXotwRr9Ilww38rzEbtjeU06
bt0m4CGp+oOuWFRvOyGtjqeTNWnC2P0cvoe10MZTM+wIs12qTjpU9kB/TEb0RfGkEFgSs1+l50Nh
NMjhI4DhEv7xeH5qlw6pXH301oIKMP6hxeDhqNI6sCl3XKkzhr5HMS98T+XZOCVDoWiW2V+NCVj6
MBu7Z5QgsS1aIHFJV1402iM8e0WXaIaUUFcNrlxJrHHq3mgNE7WJ2eFqozVX/dtFofkZ471Bjgu8
7AMZGajO4AwojVJE9hSeyMz5J/Mt2jBPAk1wiZ3GluyfEXU3ku/37AasiYWanQ5yzmF7ME057lb+
FXivwgMoIqiMX4y4t/yr7oRq3OKwNLupw9i1mIHQ8vujW6LO3spcH5VPgVr3xp2DF90yj/Pl2kWF
3hSRAbX1d6N7Flw0+JcDewj5EPygG2bis4AGrYH+Jeug/NW70aRZMscFVWeqvxzfYykH3fdULHxg
YmHPogLvVglrraUo+wH7lxCVGNbhS9P+mZ5ELGv+u6WLKM8j3ooaaIBLA/Yy/LVlZPN+eASICQcy
VplG5UbX3vVdgwUqtkwzMN8NWIoK+s5T1fwAgChaUpO/9cvjwKq2cSeYXMOgv+n2vRBeyN+R2sYG
p0K4NBK/6rZqDPSdl9t3dWmm7auHfRhBO4hMWGvUVKNxjuUvSbpeeC4tXxM8hLCyuo0Vne5QBWGC
0ARJAehZo7HaqVNk9UOlK0P4hPfF56RTaGmo8rN7NL4CU7n/CTIcZq7qgu3p4nK5UYMT2eNfD+UB
T18yphqZwVdIeU7UWFMWkUicUbyVEWRlcq/BHQq8iniygdQGHr7/EaoMek89L9fxzvT36reiXEB/
2iR1f8D/vbCU87YMi2ehVhMoa6bWkYmdtrXnXiAlRFg/8OI1CqpxLbMRY1R+vYmvs/R6sQA7OJtD
BZzCUTMnvHs5dgnIvvz9N0GGORLPkeXTDVhxN04sNf4SZhjDLMuXQgakLh0AJdegvliJURywK5v5
qb5Vrv56e8YPwHhYnmP3bRlqTzDJxfoNF8uM+VQ/4rxWjeu2v6LmUd9ouQshdoh98Y6DTP7GD73P
R4Mq4iVl6Vay0kqEVFTUdpGE40QcAfibcqrvlNpm/TnLoztUAndUZUxUG0Mk3sjIFOH/U/r1vLbU
jP5AvH8cjgjGO3eC3i8ojT9O7x5y4ZFYAsjQdZkSSD0NQiBQRCxlLD6CwWd4Y4ALjFDS7+t2vd7w
BkGEozeZQsxJhJbpe6vmlLQ6y10qabHFe7l9Nzz9BSq4oW5g9ZNRo/0t5I//tBHNh/Vs5wS35c+r
Ma+0MgVzUG0w9/gWfb+8DkTW3qxhIY7oJEwBXuytT5ZfRVKMAXWZ1l0FSVcbd1Os4691w1Xe0jhT
VoLnoB9eS5PZ1x+99NxzUcGPv7Px0s1afIyApSWxzqHWyZwqdDEmfOJwIt4t52pln29jnodW4r04
ooSBGBaI2Xm83JSbm+rB2WIP88otio6fYII7NhCNzYHHiAkTi99Jxgdnk4iyt9SfWvtzG6ybOEzb
OkJacAftiRIWDh0FB2McBCCj5OX2uerYbG4yOWh8dg4RxdoU64sIyCCt/WuEcIukOTd2am39qDzn
fu+J/wZpNsWFlW2f4Fob2LqUWnRqAiYYILax6t8AJcqJauBkiG0RXFom4j1zTzI/N2JPfkq1w/ia
QWATxujkkCrlZVFLd06ej781jWPCd94prPzDOmsUc78MzRsHA6cyLvUhRQB0fq7ECIW+Bn2XFJ8Z
8IjQXfgmWtt4ifFh9b7N5QAcnXVOPTycLSW7Ml7aM1WT4ZHSJNsX6S1NME9XgP4CtUrRe0QOWle8
9LET7vcTvjiR3ArClC6a5tmz+xNvT4JMOHBjn4K3Yrdx4yA2nbVC8YaRTnmMsSNQfxciNkMrrLAz
3d9/gcfi/aHx3+6KeKUZaJ4+XwapVd7H6y52/Qe65sX886O8SkpcDKy4kM1+3WOWw92WXJ/UgMma
FBDoG9dBzp2HcjSVXBIze1JZJ4lol7d+RCA45QYEcrvRL4u6XbQOXsMO8w9bi8EoNeaOS3UafGR0
agmTIGgRIQFBl5s+xiAgDY4sPUSkZx5YKSxIsZF+ZZ/obbV2FzDqbz5CtGD/FHOxOpN6wPb2mKQ1
MPqnPpmgAvuG00oTK9pJaP7zJ/q+2O/DCmzZyqgXCPGbW9heSTyTDu2ZWGxhfsQCPOY8/AhawKaj
87nMKxjEvaRrRWrqXtiZpLgtf8K1OUkoXOjxKVkdMfps6BMZZZfcIvevpnRpX+WXm75f5mZ9Z//C
9gv76PCiK92uQuSQ1z4fseyAbmrYqwyGS/FLQCBy/Ewi5xO80Gnen5kv3x64igVdnicXHXhHWG3b
dqrSDvFIVis1eJzFo1eZt9MdoyNQrWN5MRTa2CKLjMC1N67mvq2ei2UrxuMloZFChaMH8P2B56m0
fmAqx7csII6+tFbaBssrClO0RZYnUqatfXonpPTwpLly69rFfuMFFRgO6Fqqf2MKp6ReGIewsbsk
T3yIb8crEHTC3wtWpL6ojzcj22pxExAw3DlSJCXl6MrkQdJY8NDI2stQBUYJeRgwPmbVARk7aTjg
IsAEdrGcFySggiDOl4h1eMv0yAp+OBhFHt950XeV8PtbngGRFICpug4v3wGGo+I9FPfRxtymgjQw
S4NsAYj/rD426GbovH/2CbhKiA/LCmAzGvqUJvWuZH3fwBiI9IgJt98l2hUJg8NFG7VS8kGvrf3B
XdqmcYtVbeP42UkVvB6pL+lswhtTPWVwBZ6ntKJRWk6t9Ef/xi4HnzWCz366FDA5YHheu7OnaDXI
NhbQEhiTgDbS0AArIdZXHLDtoDCJrK5zI8StdgcsUwAsjf8TPAKsK+bVAHuOURyNHin5YV6M2dLe
vEAwn3kUhiqj+tors7MKwQw9CvtxxkA6xRT2P44qQHafLASiu42bMhNWoSytu4iFzl0BSLQzGGEe
Sdtgn83CbeOHjXBrlUeDdWsfAMVs0OzwdqCapxP7mgpq9DQxCTSeA3RtiYVWbW74q7Rc/AFuuyHX
Lx2AnfJy8tvdJcHekFwLwKIxLAQu8U3E7NNA4LRdsTzWOJ57vGKO6qIZKXowUmWNCSMX7EmnWqo4
QIkw8wKAxxOLCmKuv3GTWRXvSjB+dUBPfPLHKchdxQ5vU2R3GUY3qj3S+lOPfLvR2phqzMtHO8gl
kGJFiUgtsR200T1Lc1aiIs9+DuOQE9nI5tWbh7RQ8yIHn5uxvPEqXr0mlRA6lGk0qLzR8Inhy0Nb
jUPc6JZAvp0UWKB3YUek0TTN3m1TDLwC9mmNBe9cKo42vTHm+eBEsYAynLClFnBnqoIIpnLJL+VW
uVQlNIUFraj4g+AGekZ8v5iKuAInaNxYmF+XjnMTi0wd7UrlUDuCGX5lap41oCYQGjmq3VBmGarV
WUKYNWcUb1Illh37O/+8wY3at1ukk133ZGhapOfodiFXDvsiRTD8ZhvQKiIfFhOsPlg3IV5xP7Er
gg9fq2yA9wlVYplTiPPag6XN3d7yHxwcVqXxkDIGuoDccNpQPyMsGsb6ALhlR1g8LVoa6/gWBby/
aUPQl+9k/w9iJu2syONCdZmJXLWd/uDsK6+72LlHrTzeYsIK3p3hQE+Phtfgthg1XK6185QyN8bT
uPplVuMlYgZpPpPwPE3GtOreRQXiu8V5Km7zUBFZjZrwjhf02se/7vsZ3VuX6QsinLT3F/LdX7r1
tALnIi+dOR4FMKWvBMoinMDDvbXemqgK3qV4oVk6mW0WVmn7MczbgmzLvct2DLQeF2yJfkCq7sVw
FidLVL6E5Yr9PlCXezGy4nscBk3654nqsW+3Q9H4mpssnMlQjhJXakO91IoW0XMvvzIuRjY3E5ep
eoNwLlSWXvxrgMvRRHC1kwdgjtCDDu/MELlVQR+7hyuJO5ivo9gb6aUjOD19GGC/X0OWA6HXqKMG
9Ek2jFEw5V66xBsc/FE1PEKtFLcKVsFP7ngjUF0PTL2SJbVUaXIENx5xljpOqmHMbsef+q04kxv+
tpjvibGceBOg6RwZ0cBpH2FQ6R8F2IlPBbGXaE8J/hcME3iX0T8gW7dOLkuHBtCRWld0KZd2Sw2r
uzhIKtROoiGMrSYw8tRDBTEQfYiwW9ABC6h17KpMaz0wcUZy9w8sKztg9BPi2YQ+BzqEeYdux+2L
bOyJSTtjPxZmwra60GpQu7U4dIU97RIw5uKXxAL50DozAQMjevQ8tlUqBWwOIP03aooWCWvUGJh0
H2nZWpRCkQ7w9ZJ2gzix3mYk7Q+tgiyoxHyrAdggNXYBpmdstaTTyBZjvBPYwyh+k2avmDCxUKwf
Pd+0Q/KK90bNSG1A2SqoyWa8Usi2u3LwqR6GFO7yGY3RWFjlOTLVIWVVfRjtNubcsCOuR+H91meO
qxIkwMdzwLFxzT8KbJEQSgUMa6ziAydiE8dzrCUX0DJcxfNBqj70soYcSvLvFLYPPvsxUK7XoV0Z
74lVGIR3atDZjS48sk021W7xzTpt/1b2Kr4Bh/zoCMMwgKdMl0H2pSQl+NsotKv5LGT5flHT7eys
/R/DdO/nYA4k57YxdQToi6r61ypSMuDjpJw0dlqOmKUeENpA/W2L4V/vWoCRLqVMUVii0uobeAPC
l/B9R2gpq4S2rI9z0aM+2QoneegqOor75PW4xIc1RzOZS3R1NYzdybJRC2c3gSKy152etYux56Y5
98yAgJJqea5xPhP/S/uabDGLHyUBlf8cD1vvDE4FNJovLMTo0KNjEHu0g39KVu1RWcjt6IJP5/D3
lqHYTuJEGx6deW6mqzW8xbhl3adpAX7GecKc6S8Fk0bvWs7fJdXQvL5Ix2U5SmyefIzRqcH8rjhL
/pR3/RfXjHVeE5+9+P7S3tSmPQd9tu1q7qN4WmZsupy/rISBl9PA67t6r/m9MQjCx6hvjMAdCzWq
wGw0suum5IML6CQCZH1l0ilaKI4+x6gzwBC4kC6vR/BpTiPH29/t8pOswSLmVIi19dsOjFf4vUne
V037kABBVo2U6eNoHfgoaUXjCQyVJh9l3rsrcpUh+RdXReFm6yp7YmQABdWtA+P7V25AQSCzuXCU
6f15w5CGOpM+tpzCQgRJT52lhuu8/Owv1adZ/TOoT7pw2Esl7PNT210wqP5+O15S8yrQpXHve1VS
/G64ss2PMs0=
`protect end_protected
