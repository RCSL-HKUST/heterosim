`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ph0rHgudn/ytYlmITX7mXwt2C41xyTbbgNvdtYoqw2OYH6erpfIi2xkCawKWCHqEYxib+WNjh5YKk7l6m9a3lA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pJ1dlq84D2FpSv4x1Y7uAaoa/hbsFut1DMD5X5Yr2LUQmWXTNPI4hw64duk+HTwlWtEsbLIIeH6SqSP+ovvdGyfxA6fAtVvFe27ejAMXNfTPRfWeOeHTOlr6XmF0O6c95odmUVFpG5qVEJR5TwopK4tCYcuV7nnl72ZPv6MU2S8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IC4EGe3NcygSSVl3BgNfdVBXsnnOG40UN6SjA609pBx9Xdorb6wDvk3EZLAYNuINgezMZoyejwn9IBHjj70T2GA/Kgk4zdeuy92VvzUyn5BHmUDW5q7hAbbf5V4WoP1Q7Hqe6+a0OqYKnSaL/2vU50XsB7kpFtWnw0jpLSO++5S20k+gPmGxhq0IbWl9GmdESzx+yqoo1BQvOSZNM5zbMMyBAsOz1rl8nCPRH/MJT+tprFv0Ghyl2FbscK4cJNziJo6DVmFpfkmRc8i6YCEAUj5Cq6EyBexNfHMu/rw9jV5YBNLtielffzZ/KcHB1i5MJVCIcLjubwEJXd0XCaG5Ug==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NBtKdjl2hrtLgvXuva5rckTs2e6epgsiROZ1jUO1mjZh/o6Kg7uy0XFfeOCKw07kYqpJ6blAFQEM/yvEmuD9wGWJbbva4+Uxc8WN5396n5h6BXcDCP08VXa8dDpMoLE48gKn+8lHQJbAA+jpGgsDfWr8lRD2prwn5Nxm52Khvgc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Di1oECzdUFX0DIRPdh9nbNXDYn0CxWOZci4WuW8W3c2zUBFQCpboe5C0jylxNH719BDyIjSgPjrJdWpsJ2IFviKCC4bCtyN2MtZ6M5VtJWDQobsESKVLds1nchob+WOw/d6WMhdTwXJkGi7sHsbro7eZxfrUBwAi5XcTXUM3cbJhntQJBCiKL1Xjzg1xbsu8nKdvWU1Er+0ckn/lxAVYYtD8uZ/TDpi4eoKU1H77kG2P1SJoO2jFcHVBVhvQ9xCxmCKrCnEnpksCRZlzYrLKCWjKavrokxRp59L0+VruYn1dVa3qt5UeQ1Bp1WtYMo2ne5RW/jHcW+CVl07QT+3Abw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24090)
`protect data_block
1MN2PNZ7Nkin2/j5G2I4+qgSFyagOhy7uSmRWPymqylNm21DGysvX02hQTPllbCVj/55kh4Jjok3
+8M9T44dd4lrHqVSHW6fYFU7Kc2f0ofa5fnrtGdydnjwRDDIk6poesOTBFxFNuM5FNjDYinIJwq9
O1CWxzsBt8W7OSgzeAAwWFFHxxcLwFeewjzgOefAId0hoWA/v7nLYzik66S01OkEnjrZErNBQ4yE
HEEvILEC1Yd6JgE/C868UCk5QQjEyrhF1Nm1L2ueeS7DJjFL2a0A8j2lIeQkciDZHY1Z/EqjEnpA
iZzSCiWd3E2zUCT0NinS9SPMIH38KlYBNlLEuhFxtqSszSRvEVZj+UmZDaNtNUiUviMuG/7DBUUc
Ymm/yLFVJfa+165ie1erMLeZ73zWfmLItqRkhVbsvIfxXbc0H/MEGeBopzVWZ8je5iyTj1FcK6cQ
u6aBkrLh4o05Ye8VYNlJzB1wjKf+7hx0e9Q+zm+Mpaz6FRsIWzBTCwu6dcy57hCgCAynKpnV7m2/
5yQYDXfA+Pf18fHyxZlfYkAD1eNxI0b2tr+9LnYsztkPpwNjfQMmy3CiQPJpN6ulJsuAV7NhGmS5
QqPfkpr3q/8OHRDVrji3RwANO0dMfDe899MZ6juZfjb0vGkNfQxqMFxpaTW9YpyfPDzQAqmEqtKd
451vmVdawzGr9eL1Tph80Fd+ow1RmNx943/I5/MOVZiR22mV5T3Lyle7vp8ZhB48dVU5I3k1x8R7
xQHfnWoZ/0VAgpLFqczEt1Ozk53tAsQjrI9LbmDz6VWd5pbWehpUv42KCusgDcA4YsBPxxiXDFm5
XLOq18JBMdkOhYBajPdLIKv3VFZGvHtOg2+x43JlS8izVxNVP3ddJMGyD/XU+cWgGo3Kg3gk48yS
orJ2OFZ8yjdYe9u68s5tr2+Ou87bSYsD813sUYGeq7M4s2uzZ0dI4EE8DNcOQDTu4yp6qzFh4NmN
xRo4vTuN3QsgzjxZSFslQbP26eXHwYqFjjtFrTl2Uyw3AXRpwqvg2s+qMtQcKeu0E6LROUzR49Gz
bYMwRycBWPKLAhPG6aUR6Cp1PXhvuPUNNcD0ZjfQjtPdLxgOJhXWXFcRMRstn0tg5g8BCTuT/ggz
cXSZLol35esx4Z3aBDHQJbp4H/K+gyZVatWCK7uRZCJtkj2t0mvDAp6CWN6HdfLeRVioDMht5d19
WiHNWSSFZWSYxyfo0naBrCfT+uhQgDI28+w77QKHKneRaWHOoPhw7I4lSC/dGuVHaSp/OlhBPGBp
3SOh/p/2bBLPOK9by8/RMzZBsNf4lDctqJvGTK5A4Gfs0MXeo9/32l4+0u84lBYuIffSwCZ+xThL
CRyqLrQTx2u9kfip1mQsABXGPyrzPoXlqcVd2OG9axL8DUxkOOV641uUsbvVWNFlkN1nRgS8I2v5
PEea7DFNOjnV9RSm709calGat6UDOezB7vO77Z2gBFFQYw747deimhS6AtxQxVV25nM9/U9f53Gk
mns11hWO75ZrT3VsLbSLAX64gRhfqab4LE+NIkcxJ3VxofQchBRgXAkGgsiaM3bSgo+37wkhEZoJ
zJNlaZBkVZCRJHU38kY4xnWSuGdDJSgSqDwMJnYGm5EynN1M2kheWfrArhaVYu0j/qbET/VPzhQ5
+llTB0HdYLcvlw/uM1RcYUzHnZO8xtSFofom373M+AS+GLF47b9vinnoxHdku/AvP8BfTtqsAH60
5IgwjfOu728z7Ax6s76qP3ATCZ/C3m17S7xZ2oYKyBTY3/leR6qBRcGe6Rlhi0pp/reG9DBk3Miq
6IPfL/zrbFb43054OgEzCAP3SiA5Za3Nex0eCnoEJZSL003QOUQtbuexxEBiAgG920b2wc48xSvT
C1QyiRyj4QMbXPmXxmoJ4y5MT/G71gzQ76AEEpPb83Eatw91oRWxTx4xuSsud65v8+DDLHK5VHup
R+fASorOhCNh05XPPRkY+Nbzmz4RFvoQV/MlIhf1WUQb0Or98S5NuDVzurojcxVhB0lG3v96RgFy
mtwBb21YXGooFBGiCLx3/COV2XimziOqP2Y7ac1XFBb3ZZinwr+olZwICV9to0QTPCyR6suu5xwN
KeP0+9tO4PxKC+hLXwGuEBxTbYIjflFPGuck855/xZuj67rPbCRAw/m4WHvUpyRC6EsfYBjs7Q5t
LR8N78kYtUHNvekv8FhjYL6xNwbrB0UpVh5xH7PNOAy21zS1H5qz5EDLKdJCFF4ypksVQEoUQIPJ
YdWejOLZzIedvitVzt2oDbQqg7+vEfMQXxtTNx/NCgqlEUe4HJuuz9UmOWayZj9hzfwwtJf7XbKa
nI+qY/BNELcZZry2ALiWcCJAP4RrKZjIy2RHZWlhGsKjrWNpzJT3uoHvB6yuiiORDH3hZvM5PoGN
ZivBRPgM0cSQGk//V+nAuBuAfND6VPkTXXZ3PUJnBeqDbk06apNTPfZdjgr0fcqbH0Bjggad+kJ2
SGlgg241bAPpu4hs70TgRjHuzdWZ3SHQGx8vc4n36mSGfj9hZsUa35CA5zxgT9Y7pk9o/VDH5xBj
G28w5FZM7d4VI7mTVqr4NV9VaWOgex8mPJgtzbHNPbjSAkhn8NGgI+rdsNROsDmjx44vNkgFjSc4
PR3mfOYOZzNV736ky7gFB3arbjNGiV5gDhkzvelfwEDTBGAxw2jAXJYxNBhjbjy4kljejBIKOeVI
+Y+VGaq3fn37Awb5ucu0C8joS9j8S7X5hq1r0QZtPoszTa+3LnKpt4xKwFwtIkW/owqkVXNEsUPr
HtWZOklZbsm1Ef02IjCedUp9jDNuLJe3klTIJ9b5Q5QSkNfQrnJcdWttzG5znYvupkU4+dFrc/hC
8aXWsdXlGIMQNLcuuB/+CpdHIiKCpANLdqOnk1dH0m5lumiyuVkBoAQqdtxP86cR3nbCfxmfVN75
0I/AN5E9jyQBl8DKBYXgY5OmbL5yfr4SPgKaE6QoGAtS/1m7F8msRbLmKKCOJqyFJt9W6fV5ANzg
yQu/ldqhmBdgghFTuzsx6tRu4Q42PhZcepIAwMhiVqAmVFOALbwXZiXHSRhXtx0vw2zBmv9pTIdv
TY2cgKYK5pzyzvrf0+eH+K+OJHRVrdOI4tYVambk9eHg6L9+C28f9/vM5vBFX9vcXA6nCSEg8KNY
bC6E2vYIJbgRV9iGUqsHNIkoHpL/cbyb90bac3XYszbBtBwExF4t5E6emTz4tqb8ykHzb8+aC2Gw
5MLLXAVBnTxAVxJDCVPkI60tmr6ORE4pPG4fgFgioIvitTUPeHmKWwC19cM+/eDsEVfTIv0Kaaex
4GyVr1q7+1OYTpp1Z3yIFtbt0nb08v2q8mEkNk7T4eo73SeaGAsBWhfSoZ16mF2iTSOcsb1FbLMS
QpqWv4KFqyUAZmIyH5PvIC8GmddPmvObvrqux2OG00feo3dybrnAsj8w/GTMf7gK8vyaqv6tP2ra
/PTNsdWIsigD3qaxARlwKyDsW76HhHlJEbXBgJaFZcztdAKX+FPykiN96wvSLRpRqevbZrGUMH7w
DW9gYMy6vCOD6B6VCIhqSd4wLxGNLH9UhfXcyY1jVIFuUnrg90Hm3p/Fmg/4rwLLixJxovXot/qN
MipXUPw6TECXWJJ4N5kxIdWJsOeg9TZfVabPLDQYsuGpNICsKha3gHUqQZVXtIlFNMUp2qtH5eQJ
LPIRn8Bz2uFj03ZZ5su8Mmnj89ncCCLVPczAJAWX23khYecK2xy0bzlC8bYgn1RRYFgqHVjwfeZz
VNNNnxFnfE9zRoi40ZZwcaUH+NH/ter9Kv5Jo8XcZ/IRoOAaSn05nDI+WhdCIZCCp08sSKUyQilE
bm5WPZOr4ULODpxAQw3faCKnGJ5tyeZmRxRlc8Lr9HHQz010Nu2J790Le9wJk5DoUgMbX2VcFXwc
PQkwMYnFi2Rx8049qMqsWaLIMKTmYXWCbIJ0pX5BNMQORG7yrRtGWipLeZNAki1Qf7PgbzfF81qg
k1Tx0SYsMTdOdzpSsdBnhOwtCLCj24WHIC6gQ3lT05bJd1o2L9AFO4MckFjsoGtUGmW6xYKYf78A
te3F1//W0CdUcNCB4ItiXi8brqXDYVTRFVCMRh+sPKJO87lsovrxT34b2ebbBx+r8Yus+hizCyfP
s3wNoNvV6u6ppFZ8kBKSMgHEUn+4lCKI7hkUP7eauLK8OTrIlXjFa8smp+6/fjmgugwCR3UvkVzO
1wBJE+4xHi4wlEGviG28j1nAF24+feRKWzjc8ZeyGypLVexQTZ/RLkYYeFAi2b3JsXoYHff0DbY5
xtMqd/W/1nwYLanjDvkeuaJ9+TAmDJ4eMnhT+Toe9cjM+DeVoixyAw0hbeNEnZ1GsTTrYlXXun9q
iDD+RGfv6XZbPIpK1ME8q3HjpkZ5Tq714HYwa1tbJSTrra+R4wrOsjw/i6Z7CGGO8o4ovxDSbRL6
K0jFen5HtYYL+6dUQ8UvWaiKvCBt2zvB0x4e6t8rD9jDwiisgMtLgqahaN0C8YS8todAcqTO1aX4
7r72pHjlx9qMzTIv5ELfMUfiLjJ6hbVMv0mU9dUoDKoYDY82Oof3lHAe4noMmlWpRKcuPTMScTFA
xf3Xke5ZrZfWsLeekvAiXTLTUG9EVJ2B0oY+NBopa2mXdi16ZA4Z8XuUr3wNLpiLFH9NcVBlBfoI
P4nz2s8dmbEMC3dWq2jezy8XQsEyBomGImN06D+7zRN1Jq6o0t3r9Y7deSCZ2eq74sDdFcN65BF3
Lr8cBizweEhS/SvkXE5A+xpe9zJyp9LzNkWYanQ5QTDspiW8+IgYuOBaDggE/SdklsF8zGjsya71
bR2W/TvY87JiQa1ztOcwFZVRm7yN5JkUFo9wcMgYo0oC6YtAInihm9BctXHiA/M9NWOs+rVmIVuL
6ZUpVfcSvlWr5w02issG98VnyZF5BJhraLdJKb+3CbezwaoN3Ozn6rqCUHArTgp0nfjV+ApiidZB
M+AHUkbAPwx1BiFxhS8cFu7SZ6UfOVCEaIdPA7LVx/OKGzugMiAHa8Wcn5g1Ig0AWT/noXfEm6sN
LGBROndM54zyTVTj30kSSdNn13AglSLRp3jL+PZtU2EffIQ6lCgYisSe6UGAlaMuC0akcwSV28nB
CYB8ypFlT1irhUqHmEILWdWiO6TxElONneO8pOmv5jEiZ+y1m4BxlwSUcvhOlU/xzO1OIaBk/a0+
Q5ZUjQOlqaytSl19NscigaPCXB+j4aaBcGdCagMyJbdkoglajAV0dIHW82JSSCmM4X9fbnCJSnGO
R+IsSQ+l8YmGesd/T1exEeWwEQvLELP1fpNoP50lfpuU/wFawDM5eqxtTMfZICLfcNhkxPqMfLLQ
3dVwMkdMVB8XPYIuaRkegmtVpyuuhcJLKRbXC82vcf7VS89ruaHerPfk2mlgiQUqYeP3a3tR6J8Z
gA+09pejeIX5LfHKxK+zgbO7o3TOqcdE2tCfLOh9lzNM5wrIHQhaVnfaynQFPAS0oFJuFhPsvrXM
mgG6O+1fk0FkN8MPCJ1aoLEycSuWBpB5gWYad+IQ8MJWqA61WiYS329VfkKgSZ7wnAQovaRGeBZ/
SDg35VTk0wCXzHHI5R7eTizKKyy9cFvY8ra8RXu1aLCb56CJIL2wys89O3I28b/mFDcmD3GUbxre
6SEQL2JObuid2wBTnK+3yqvWkYfLs4JMrSbplj4Qor02NHnxwNQ8fZMwt9G6Lz/utHOJ5CnQYzxq
wi31Xn/nUreVkJ3gxH3uGgWJa+7r4r/5M3xrISWbX5QwIbsiJesM33EddREg4Rvgrkb5UT4T/HDc
Ph3R//EL/kFC+S2MUY55T1+47GW4CBH2FFndKMAYcyGpp/FeeLXB9A4uBO02c/QzGX0sVYWk8CoT
7BOKUePXpAGbcjr3c7B7BJCcPglR2kKmbz8JawtpXBqqsjutKLB69jeDTBQlWYP97o1g1NoituBa
ZGbT2xnW5ySHhe0ggR5tT70DYp3QXLf9t0glzjOomZ+bE9W1PaTxaG/mfC4VOnep1cjCe5yvpG7n
2kXaiciLfAJmAPrOZJrq3cvzSD8qF8f9t+3CJ6RA/+UpZTxw8dHucuHcADKCqyG49VkwAXFa3l+V
Tc1xbZqdGvhV0BSm3nCmt35mFzpROWIvnRdJ4sFw5xPXIUEQ6YGW98qxXFiW2y2bd3EcamEQcRnI
4h8oLc07YUJdtYd4k93Rx8+0KXBCG0fychxdYLMfSrAxl0ZL0GdX0lhmAQYKxM93k0vYmf5zvGsc
Lf1IRSDTmkm+6zrG2w1dDx3Gd/Q9jb6Q+LoLHByrGbWMsrpYTHFkLegQG0RsBsUENMZOUJ3B4CEe
OfHqH5EQumVyYpLbmAnXgaPKyy/zMQDGcixQ7DYq5AkM+Rte+PphSZ/O+1T8Y1/pULuVMI/CwR7u
grBMNY47KBsomKlLSE/X2O4+sJYbH5TbVXI1vPNh50prCpvJWiSS5BqhLKViObwGQ/RGzfUlI/GM
82L3fF8JmFEA51ko0XP/dk91pjODjbXgh6Fs0Yg+TfN2vnIapqqgs3PiB5TVmE7h2IUC/SsPPtR6
P+CmA2+hB2DN3Kosu3r9IUTImlSBnfH6argePCmFOD9VJi8AJ6lt1es8JmXWzB8FBjg2ukwqr2s6
QLuWbuf/I6isCpV5pjrRsQjuPF9Ql/e0YEOh/JwSO2tx+Ca5HnVFqKXuhKuUdhaCbtU0Gqs1UM3A
1QyhCajo6m4kSafR6ttDk/Mgij8YBlVz7oUEMrJiOTFD40/zlrFNmBOeT9Hd36wyewJue10Hcyob
K0EaSdkBb1KeVYwwOyiG6bDtMlvmwmcnuE1vabaADGb9ci/Qt/TZmK2f4HIEF+fY2sadxeuyRhT8
jHbHHG53R4vYBmhWBob1CPG99jTZUk6egBD1RaDbg48zIA6Jemg9+COCE8HisBvvK7nzygn2G1bH
UduUAhVl7jOtWztw9OqgEwx8eFcSE9plDIwFW0FL7/gSpMlVlWcYs4f69nkEfmTBZ9n4lrU7YTCp
3CZIk17fwZ4daZsBBQAokCbUk3uYbK23Gc6G24WiZGOvATR8u8Dl46nBN0jE0gvcj9hz2LbuM9kl
3nTJMGWMYQ0NBuIsz2qLNR2e9BGmghwdIH5KRcNql9Brlal5gBwMmCe1hMbsDU/yyL7hrkxM2BlX
PkZixy8BHe2+isTHBbDgOSw7EgWX4fMROSG4rDkskm3bHIAYUHKJxY2ZrgCARnc9k8aF68OPNg05
A7WzJxT/LuDFO8gRbJKgP0hQoEJ0Rs8DhecU3KlPC7zVTr/YxLM2y47Gx3iw+1ppapn+VlUziGyH
ZOxEp4nwkli6ztQC7PzocMEnDWuWFSIJJdxr92aZ9hrq/eyFeRKhB0w4u6OXOmzrzdox5cLll3fw
Wda1POPuqVYsqpDdsun3vLIKaORJVJ3/3eJmsV1KGZhti6jS6u9sd7Gt1WnLGp5fvTL5Nz070n/r
od77buJ32xNblHPrPp6p1xjgJjets6T7ukni6ur5hnqKGRQQ74dsqSkVoLQL0XtAHnJEDUeXqruN
cBuw46H/R0hhifb5BbOgVgNj/D4IeIlgJwLBTjaMiy/AFS3EzmlmqTHXGolNGmOFI2h5WTM+Wocd
RdZ+FxqCVlWkBxiC0pLRUS7uVaX8xJYOtLoqVmn6/Z2ahU8CcOdAxfWrh4MmmkW0pfjEWixvut4j
eNdQ1EHunLZMkxwCvs1JruMGGRmCHOADNFfcKuO+B2ddHnj2FdTAa97Uc4LlNxhBhbuTXpQGpfsF
7K9E6m5Tm5F8mMCNwfp7KYurMOeYfU3NAaMRvLcyPUKCn8Op+mufkLZ8T94NIHuYzJaOP3wBc9E5
aKGu/ISjp4sw+Wzk375Yw5+OM/8MPtk2GFd73EkT0fh4uwFUmCLstSB9sKVTbO5xIPiHER9WahBM
fSAJryTXfwOwliHmUhy4k4S12tRFg+i1Ex8pWiOZ0dy3l3FTZeCn1moCBwnwXH/9tDzyYxnF8Jzv
xU4NxMa4LCjTzFABtRb1Dxqy6D4UY6/T70bQICLMYtQvjHYxQR0Rxoc+yUjylyigCTYm7P3dmZU5
VNe73E1tuchc/WCuLuXeXeMt6A8bAgwF3f/iXf3McHivrk+cj49bTSwfC6CxrkdgLTrK9EtSFgau
WFNd6SRyDoCxZoaEq0G95PvGXg2WsdRSMdG1Dsz4kyScEbzk4Slw5t9a/7b85SF1ZvO3H46I5JdH
KEGVDO32Aw6fuWCDULhDfV16iysdmjf57XX6ozoFz+M9ftgznttEXyn0GLFuG7LCe/Ai6TWDUgHL
mGkFx7+aNz2OeLUxZjNx9pitrTbWVagc9SB44+Wdlgd9qmLbgx3gBT7InKTaPg2OrTFg4Xdm6quL
SFECusjHFRpA3ESO+nioMMYPMpbeARTwl2K2JDinqnxtm0TnahnkHf4zoayWCcfBvgPwFztELfma
qOySpWsTyAt7lA4mfPFboLqsYnUgT74yE4owpyVM9l6XBcXuatBSfcGG2GMFkjNGPMtb5p9QvOwK
AfGu1SYRebFP6VKHavicAD1I+1Ao6lIM26Av82pM8iCzo6T2wBrr9VExvgxDSfH1iGm28fHDimOk
ZpvAgyWjl+a2lWNr7on4SOLJ4IwEX31og6fdfX14sdyKUvb3SmABuP1Bf/uenqfc3MlksSxrgA1T
UnaL8HRXcZ/LvGrn3KgJyYxcF6W98BuVWMekVOiQMZiR7IzoliQaXSwd0RJeGZn8dv1zG4yoUKTh
pHrKBExOLM9hvQmZWpsGLDTc09J87woB4rS0l/hMx8JPvImizCpYowYQ7jMytUNRkkoh58kOtiQD
+6ekgLHUsDI36d6TsaxDj7P/4cvI0EP1vLPVNGvXzPS4P0oIQsXAKKQRokyqqa2vtBAyFJWyHrHY
lnaTeVMcigSHPYvZetlf0HZjF63Ma8fABWKoKtC7pOhWivNnJjpQYfjvZ3005jGGb0YOc/HIBxi+
vn/aBM64PDVkjCgdZo3fVqteFNfVRht4M5BwlBSn+QmPzRXXmEHGjibdrN76VR9QyrfHGYbYOyMT
FzDtn8Yp4ypzZlEb9fLK4/UbKOdRt1kKhCiZUbd3qC0TaUbTsIinzyiSNTwEttIijwiKIO7WcfKv
13nr305fFIWoeepjei2XNrz2utBBr5EFFgOWFJuxwLvaUUZw39qSN2XUcV1wjcvEM0rY1hx6PuRU
LJ/w1u/ntV4QvW1mO5F78SEzcqB9+K9/0u+UdcggZU/RSEKZu/UQcHCnMyyWht2C1g9mWwSf86R1
bDc22Y9CE2KSA3HDusXPMTMidyduOpDrDp4XMzmsxJ1lcHU2YqW66MWd8KR9svoLxMIXO3MHhnCs
WjmxHiFQb/wib+j2T02PvfAYIk+1/1Woef6Mqfu2UwB+9uRTYttZgOagoj2qVH0d4scj6yTAw/ET
eS3U09WTSaMf/upShufDkFBoQhoL7fX7hXhf/7UD1+k0V5yXgji54LLPXeb2/a/R/2bL/9i41u2I
lohqfuRK2d4j7TntvCoQ6xsxAJRgRheau0nIeEno1Sx7PxXaulxW3mM4jP+OQXn02OwthdSe4vD1
teVnRQIiLyrs/5+0L5BbeTelM7ZfXj2WmkFLDc6UHgt/SAOHKcK77EQ++cmM0L2Z+XKHbh17VtUH
Lq2qbdN+NVqu1dgYT4XXuBa9G8LbQTWBZGnv0UXaAqDgUt1Wja7UmB+4V5mcuiROtls5Qm8nK+3g
vlFleDTJqHUxyKUI+AOdamBL91kmA0nP9Nb4OKW+Zxen84oXkn7Y8G8QzUhvbEOmpMAerADAEv2P
KZ8ZHihj+10GowVXDBMBCvpxJm7UEgA9eMw4Kh641FfKltCTHTYRzbesi9qwsremwbuk/OcCmF4q
4jnPPwYcEvWbxZlJBczu568BUm0RHFq27mKCWTuusPI0MbCof298aAw/EDszS5vEGmwEyNrIs1Rd
TXYlPc1O4rWuUOB2aozcEZ/kY8aYF9cp1ZnRIIhLfo/y1hU5GYz0oxlhAOJ85Wo2sZRtY5kQW932
/7yK+K6Pkiq7KNG15RC5v66OrI+TyxLdLwTbo1T8JmnQcGeGhh6G0Wq2hzgbIaNpTl5j37rWQ5Dw
WibW2jtP0NIVaAiJ1ej5BR9gJWs8Gb76UIjmjgWGjPb9BJHj2/eBXpWxtuNj7f/gAMs7+/dqKdNy
v3824Wu70U/CBIHy1bBk7bMaaaPnB1DQXY8dnWjdsjml22KMhUXuD9A0XQeMvFHzyPz+1obF4TNh
GCcpvogeQz3AI6+7yOPptNojbQXzuqKiE4dtAexMu7O6DzkSrh5GN9IBSFcH/lDjET7CFOz7hrDH
PL6VwllLG2DPKBAHeJvgr/alFrXohvL0WAhZXs3VB9NDHcABcRwXAhGgRlDJZlYvouNKBUxypEzP
b0e3055k3PpS3LVWCHONno3jBGrhzlBpJ+ZbHWkAS8hUGpUescA38pmzLUZ85VFYkrjSMQW7lTO3
o9B847V96i94iFBQuX3J/otnno/kv2SjhX7XSWSAJ3PflqhrmgCpbpbLAv9HMbyKaTAkQDyInH5G
+EI8kOcdYoFRvR0CGg6nsKVQ7HRiOJSg0FCuZ3kmRbmd7dKtPBvFjvYkO2Iw/s4iK/WGqIRPDXOI
PtrkyytBT4zX1RUn3xf5nsz9M9qZQPzH/Sv/fhaXlvrhr+fHF7L1M046LAFuSRwcWh9Ns+gAL5iP
Zi7x/TbFseQ9zi4WXOdbhh3k0bb7Eg+9AdoGsfW1JUQgNvf9JuP+pNIkZmpZMaH8m/2Jm7cUlaen
/HhSi9mUr4myLQSW6wVumfPFGY5TxRMfHmPErRBhoRd0ZxcUui+9v+szPf3AKZ5BbRklBtRqU9he
3sBLSazAB5Wl8ay2pHclJAAWy29WqDIcFc6X6//ExqRNRYCvt4UBy2Pq9timlO7yISIhTeYQ7Y5L
FFG8t7uoAm8NHGiDFHGN9mjjMFNEZ8GezbfbjxfTrIxXP0X9V+ddQWfCSsZ+o4NZpEcc6B+3UsNF
khtAEa2nKgZ+OhBS8BjA8FjYzEJwMLg5+E8+2Bf3JXHilu6pN3rFi5XVtMVPKfDk0thxIKbQLD4M
Hxhcbx/yzXg9FI5kAZTddZXg91GSS2TkhkgbWZkW3a2PJNGdKpFqXLyFKyTzZQhyHOPMZLcLoubI
o1mfwRvvcYNM37YiC2AK+Ut3djbDaXDmGEVerkOP2BpH0YF5+xKq/NM8scYy0eQ+1qToOwMGuDnt
sUP9EG7XCQHEG4dmFHaxuGYYWVTwfX41gYcdEXy5gtcLtiXwNvnmllY95mK6ogyT2UJRzVU6SRf6
MzS0hBLu8+HFR3G8aFjqVYovfgfC/+JiG4BWCo0uYo4Og1AGUSJwpkc3cHth7wMZfeTp57DEUlTQ
6g7LipdAhcZ9fzIc94s49rwdcec5XlV8mLHfi2KQLC8LayOxHLHOA2f9DXEGGiGO9XWkgJ6YwMFc
dYKptQgIddodYl+j/A8vfHBQ39vHhxFzg+3SgbfRa80slGdN/syqGyJ7YFho5+4tHRdeBftFRrQc
BPd/LXGQR2IHJFzgaZ9zX0UzfbTnuhrINmC85xstjQ7Tpw3uIfJCi3jXYPv+5KpuREBlwvfJUPEp
ZHCiRTnwTuasJTFQAOcfw99osFUobppMEm57krnBWal3MeBuDAY0sWds6bgY5xkGE6KUqdjZnMFQ
XgKXDjRMqXcpFz421ecXwdysWi7jTNMLCK+6vdmFZ9d+aGqfldg4FLCEyIopoyhnH3xwIGA1XkPO
uY/Y5RJJEodQLzJi9tRXgtqXeI5FpLeO3r51h5IR/jlTJTpfDqzj6B4s+aNgXCd22wQQsdQl/MK2
6JnPxmQMKnOxmiqIFMiPQUhW6bNkqvACZxy0uftp1UM/QSCHfgoP+i4qxxntw284hVi8unYVDErg
PV0MUbH3OED4gxcaPPYraDJeb0yRgQynfrmvRmWlKeatR8pWyvU09MSs0MfR5rZaSyvDPAwyc+XW
zUPIDLlIOI3S83jwcxhTzUw5kXtIHkElPvCo05ekR0m6581qEdFjb7kDHN8020YiM8g/MGcNjxzP
Eb/7mu0Z7DbulOaERlcpIEKvsFtUU54UKUQThkXnMenUlwJv0dSx/IXsxEzBckJoIhfhe3ANAe/A
awRyPPQjSNgyNMT+C3gc5PV2f4yozLPZYXk9x2IIwOTv/4c2xTWWU1kDdr3M70olO6+MaN7h6OXJ
q8E4TmFdDH1tgT2ENu/ViVtVA6/IBxzgfAHW4ixspjSue2YeSno6rRLzIV9wK/Gqbw0jEmwY35zh
xQN3LQ7vG408HAOhDOwDRRhuifGYHCUVetBvVsQSmlS59AXwFRHyQir/BrOOmUJ/QlnCFKt/dKC8
nkujMafSGoEDrN1nYDa3p+B+IY6GKqNlhjDhdvGuV1BFaDZEcRn7WjAe8mnTXMdlB+DdPkiaZAWU
+KWKVl3mkKb5rs8Zdrmw9GEF+f0lT2UPJtVGT8WfCrI1la0hwF6/mEIarng7Nanpp6IDk6EPZxek
a7NZ93lkeRjbgOV1y8OnD7juMFpCYOIBCco2Bf9n/2y4ycRAunBnwVAlN8ZqK12NOsACxFV2Xqxt
2S0O/gMp3PRO2j0qMic3960xroDvCsvWfZlqQVEWyS5iP+0hFJTXzCe7mODi/2GWCEanX6dYVuDj
fFDxIqt7Ofb9aD0xay0BhxdrCTv6llS+kzcmlzbcUpnvtmwQy6ToXyE/jh4YVGEWg2h/MOhf6mTq
b44LWp/TSWpGgv9zKCFsX+7gBwZ44hOY4IFWe/ksTvjUhMhJQ2N4kcR7XWLRSzMYGizeic6mmXZO
eVgZmaYVMH2RyJXuApoGzKiZpl2SiluLCCXsqJRZzRq0vRsrbtkWip9s59Yg6gT15VJs3SYf0xuy
gC+BURxaCE1jYJjU0yZU+JqouSfg3FplrgWdXaX+FWvvimV05Rh5jE2DljHb0UHxknqrnlylBAku
ARK278u2ZC8tEKc67FHuS/J9/PfBQu/NGzVsT36NXlYXqBAcZrufYN9OyXghZJu/GYSNh4NGhnBi
BAixM2PtzgU9pp9A3MFwJatmUJUM4BEWK/RBSaCeJS4E9daU55QaVxhoj4tzXgGcADuJxj9UQwMO
pbiWPqqlgVNBDlVeqRcAFsWLQQR9nG+cyfO4XqNWAkCKhCuLxEYGIXFu9eR5NCE+WK22LJHwK858
sIQMm2iGIXkp4FauCpuW8lrzPg8sGJJn2yR97jJVZJmy05i2kUnldJGehFYXZMq0eOqnhQc/2QNy
Z/BgzK0Fx5/j5nkkuKGB5MI5/FqJo5xqql2ZnHIwkhSmxIM5CB0DijFxbZ1/eht5FF1hRlL1xmU7
ypIWNYWCNyR1NnfOQezi9lnNeeCEG7DIVb2KueCzw1whHyxpSPnwtzZMmqv2UCdzsrOb9Fy1cLqG
zat0r+hUvL/EQPOEb7849Co4bRO0zRyikRr00bIGccMsJFpVCUks9MlBbocZbiV3KXYbJN2aS+j9
E422NrOoZlkn3K2gzC8Yyz1vpX2PZbPwNJR7k9LZeofpvesRxR4l/6vFzwvJh0kpPuIz37xMjNSB
KNmOwOdvbnLigeRVcvNeT4iZGmpgxavXfogT5nM+Ua3X/yET0AYg9CDgN3AVT5v2397zXDphobW7
ktEvGNlhjQeiJ4XCOq1VXAdbMKEVGN+Uzn7k65IEsoFpqU8cXzndwKYj6dDeN2IUb33DaEYb/JT3
FX9NX47keHZu8Knt0brYhavbLKzOtstMGfb4PkWzAOVCAVYIUue2Tp4vFf6PPXbKJ26Nfx2VGFeG
V37++cS47RBSoJJMcRzAVxIEs1UrqGKN9etSn6xE87lN0Rbdnunz/9HBEgemJDcDoolIwvvGzRPP
/04qwoxmojVzIC8ngy4hCh6CNJHm83oD0ZNt3GEHfWQSpv+FpRQ9atwAkEdWRhoGwMd6E5EJI3Va
i+14p5usIVpGxVHUpdMlzfEifYSH7pQe+/jHwAFutkROUZzMflNle3jV2RC7yVsdjBS+q9JJzN/h
lXNSSYBu50pizvBjChlQ4Z4HNcoiGwqxLjsilJVFP8jT07maFeI1I7C4GYCicHdTCZEuXJmwkW/F
3yAIGpaO4vKi+4YH+e7ssSQ39xj8upgH+C4A85J3LuFEQN1cilbo31YYIi7JUfc2q8NW7GaZM7yW
1t/cgY+goK9y9GAGdLcKiU0/OLVeq6ti+JSAGkWz7lrzrDoCfUew/ZuqxEKBJsYI9n8zk0It/PLa
ATK1hHOysZgHEY/itfaEre2Tt6Bzm6aAPLRmd17YFmqVH8WrLIG/d7ZHY2MhMcOLRm0irM1yeFdN
mGKtfu2myUVKG4tlRtN45ip/NitfHDNxj5tlGyi9rnD1WfGx2rVsjo2aDyjeAwZcRG7mBj0uzBcJ
kPNcoFtNjqZ/kgdkkZ7pk3BHr9dhZkdoKBB9fGGtqeIPiE5uVLvudgg3OeVf9DNWqAlbXajYgyly
J7Y8FkhGSwWppyDvGF8yr7Pg6bc6Bhvlh1IP9GoJ/Iarl08W+DVPLC9EnRMWot0xQmUeJR06qhDz
aQsdP9Ib8H1x6IvbIcqnjAG7Flzdff7zCERqCFgax7GS9JGLxa3ljDz6DWMqprm3e700XpOqgj8F
XP9a6lRUnsaGeYFd6z/HZlfK0Epn2UVJn7Qs5hs9QR2jLiBdliyncf2/KBNukyWqtXpjNI+EzD/y
UgXJtDyw1PQu8S+qN4hgehufmK+65d2U2SBQ6ncABsAkJi3mu7yDKTg0JYnwza5w6KukHRy3GUu0
vt4gCDPT89DElRe9EswyQZTfY8uq+2jEb+10FPZ+ofBPr4Rfa6jkd3MDIandw/gFM7u9mT433Pa/
1Da2zoTLp2UcNOMzlaVQsHplYb2DtDkrC7v2qu8ON01vgcauWh4nrdDdzFZYs1kACmEmYbNdlgJ6
QyZyFY0embZKAKTKUHXitpBeDAxnerXZRshuETnSfpdxeaHCMhlUl61OnBn2IO3bkUTHOzQFtA5W
7BbvpWIbUZ9t+HQ9MAjyAjMszG/hK7chsfeumuHWoo0iig27UD1gMTR6iJMWZtld/ynMyyIjk1WB
PKnfWMIgtCGt1X9gkgJAS6LHd5UlD5CMjor7ifgD8kAjWJKh+aP49A83xWHCsKX//S1GJk2Y598d
v5Kp3mnQmZyjuEEjtWAlm+5Fgc5q3VQS4RjSZ4XIzdk7JUArhDPjMz9rHFDfy5BOPI3ljBGkCc4x
kbFgidACkGCYp0G/H6OWUBoerpI7RnNM9jsqlM0v65En+fZQzUkMWLsq/nJzLhFeZZ2wOL2NnHpn
0KnCYDPbxiocNVd285t8WdSLKiiG5bH4krwnKG1tn9V62IuBexQ7ZmhaijgirhK87z+IyD9qjti3
dmOqpzdcREYB6PNV8tOPWzg0+4QGKM2q56MT5tLKh4alAp6PwHQDVnwYeVcLHx5OXyts98Bkq1Wy
VX45Qs+5m1dH226kDDgKnjDK4ZmJElNYN8xOtnkZ61kVENkLemGgIxT5GfhBvmucuBrtOOMg7lY6
voorGE5sKswibij3brOo/VlX47XSqBWlIEh8XgsY9EE5buPzzO2R8IJvpQzpjOOQukLrBznVgjIH
srQLpHqen3l03zIN6ICsdXTwDIMcOrpC5TrlJl6jMStSPcFnJeMJQ+QpsxX8V0gtDOoa99EgpxNg
WzasYM+Id8qeYM8vSjm3Y+LDRY0wsYOyOxZaRzm1sRCfhlvmBb8m+ehdnPV63zjVn+2NKfg+NsPx
mbzwRIfAb08ttnt8qw7Z7Us4SyHUr16zZzUKPZdxCFhRiP1sdZ9Xulh0AKbnvdjTfMCKmH7vtURF
MO6dZVBQspysrfZsJYwhL81S0qFle24SBKqw+LgkS0xpsMA90HVU5LNV/pQryyjELNIUBMpZ5V5O
cOHiLJt5s6O8lPKIauAca98X4+ceOPmGqo7KdQkbwYsEpIs35qSpSOydQL/u6C+AmOJt6tQUuamE
fOBhF88i/H+gGSL6J2+oWvETQibxX1HCNsdBUFA0Cy8LMLaNRzpF1Ag5/fEDGmr3rpEnnWXfHT+y
Kkg9ENXAzIFA13xV0IZ8I4ykCSxKEOY6gZikoMqG/vmMzL8iOZTieNN3fv3m0AjB+Os+aJtgwW5f
JmILdNYThMxkWfU6H8t//YWAVbmmGI1pAZ9g+GrMNybDRDS2YkJMQniLd+//MK0wMsXFFYPz6RnR
oxRPO61wEAllfWxJ0BCv2Yuc4LLZa2WkjvCu0o+lKp5P3sUSQK4BBpOX4aEIJCoWFc6ZQPXlZHgF
yDs3SVNuiP6iCp0hrsw3auv/9HBqvHLqbG0wmj0iiiW+e9eAmvrg2h4wCwVdgKfIBv6qRSPoIGWu
Crmr4GTOCT1lGVFPOlmb01hug/CszwcrkK83w1VrMX1WUeBmoIoPC4fjWL+QOfMHWj9P0CiPkLwR
dFxjQYHKglbWVDYXaggLvZiNZyot76//uykcFPEbLrdklVhPdCUGu8Wu8rgnXAFXFdOKbu2S41/T
cPgq6a4UQfAT73adkZrADYFaIKvuKJQknkAuUClwSAMsjkVKTJwGnZaPfU5m8a9UmalziDgR3SD6
/rk3Qll5cKf/Tx0wS+KlFyyr0TuzJXjZtbcKX0JhT2eqeHowN/8YmuYwhUAkKS0kZluOzVCMGt3i
qdlxd6+DFpjDfXWC3bx3FbD54HkVVkrfTGoHym6+JPWTvh6MEAVQmSv7NlXmBD7xWs5wGv0SyQu2
SDrozPbtIcFZZ6aHsVcyU/A+9aP+uVMQStJAmm2pNJ183+Bs9baenBdV/kBK9TdFYOn534IpqSWY
vVnPQM4av3C7dRepCe3hzZ/TdsBCULW8SkkzTjh1gYzCSZSlfB7cwlvD9Ma4h+Bd6fE+FQKw032v
tzmNlhryk6n5Wl7cos7oLYzZxmMXj3yA7ROq2BtRtdfP1oAF2pDyoGKGoOTVVZe150RvLXZVXhgO
jJPQNCBrXOcQ1HXVziCpLqfiO5FK3n8iwP93T8jws1Z9as8qxtfLd2KHDCgWwX9oR8ncYMVVBNi/
1PHjsKEOBRltFXSI/bBzC3R8PuS8AjHbcE6gyWX8odF2OoQpiLvgrudW55fGXy4/w2loqxOZTpG6
iXcu3lBBYI1mr2WFR7DseYj0ggBXEF8bG1o+v48QOcYZc7pD/2CeYGnexaso+oI0rl7bLPJBNT8c
tcqgP5SUjfb+6LlV9veOUU6mLoi5DsPornTxQNXNvR6+Ap85hMQIm9V+TjfaAQYIQ+cnNS5w+4Fb
5AODbPYNSUS8hSHGFrAz//fY/rrGXtYbb9Iu6zRelENI9rjtqGI8DibNK0C/QWO69QPylgawGX/u
z1nnHUzMJbYgHKtQiFWKdMMFqYarJf3KS4ICq45Qo+i7hy+gYhrBcgDlriiBP/rHGrLEmQ4DgKDa
SPJ805Sf5zjvzcrujCfri36ihG2wFL1lsmzc1WPlvFIU7W2AkK779iXZe0N2BiwKd+DBzHSuD+PS
Vh2LjxIquxHIlfr+BC56xKKxBoznjoD9xGj0ycTduJ4BID+fV1WKiHumjKqM7ERERXNAAXCMjVD9
bzwY2rjkXIkf5ZeUfMNLg0+RE3x44VJw/Cq0TDFdTGzfOmZyE+Ne/m70Ily98v3M719WTwFJDHHv
dyRmxwm7SvFWpXcCnx/oAXGohcbTBIljlh6d3d1xwsEb/JaaJdh/4i+dYchsmXNmUAOPn4r3OIrl
NXQt0M0+DBAQ/0zTvBKyZfJMAMn7yRb7PW+2+qHYX+LaV8eZ8TwClbPPcmh0eyfYo2WlN74vEFkU
4yJRwPebWDE3SoJ8WZRi+yHX85C6pIBDm/64cWBQLeRYE8WssYClZuFWcu9tvYtODhZpUi+jibmb
II9EHHDdHduzWZq77ruq9fyitJDPfU+0PfA+mUv8vX0f38NKI09eR0Irz38VaLHels45uKy+TOW0
VQzJgeEW+KfV1wX4NlMHxjTHdPSHz5MQJOS8SB+4l9bkab+ypTHsyglJjjmjanEH4Nhu3ElaILeI
aal4O/BA4oJiSAbuwULNbn5k/E0+vPdB12GWErG9V94PFgUy8i8D+50reDs5l1QfcHblZCBC0dul
L9UpPiPH4BlVs5wIK4vfRX8/lmqf9Dq7Z99luB1D+1IXQYRg9q/uI4oHYMT9M3hj+csRrS3EqI+n
8MW1Rg1VotcfKVr3DlSD8wf1QOQTPVY2EsKE67kTOnw92uQrb+wa2cU0vzB+0ieHS57sB5CoEidu
Ff9Qa06/W4Owh81k90XZJiuS9gvmu5JwDuE3BLRUFYB7KYaRDBr1KFBIMW5f1wmyL1iixPZvvDZ2
oVkJK8v9aYxlZWqa4ZCBq5QjXNnT58ZErftvfujwEUdn2REDiVhB6LzoXZ2q6u4G8NT51TMHZgOo
+QQkQEWbvZrwozr6q+WVfzvcw+/+LOx6u0Bfqu4c6CB/QqRyLSrlSZhNziJkutlL1NzhHIGggAM+
lVz8Cj5nd74XuKHhoe/btFJnhZrEanlwUShHjEGIYEbTRNPrITkH4STKI6WIxtKNqabz4TS2rd/4
MMA0dRFlosohAp6zSjigF09lldyzZ7ihOCnIY5TwifENUkwQq7/o0KtF4RxyTm35ITbQyazFUfkO
NWV4NssznQccw++RyGTrS5ZC6O0S8I33wlNaXz2X3iIMAgyQHdRr9vDOiH5U1q/p88mBtvRzqrvj
Huphy77/n4+g3rUhdXd/0eH0xoWEFkRXWZejsqp0mZ5hVo3snMxMl7Q1kPKg10T9gbMnOZ2OihQT
qX/rVxHH9u2F4JvdyLFKEU6o4XbbwBnIK7MoTPABOKoqprM2pehsXEhHUXizBrNAXFMxV/Y44iHX
WsXsg8MZGk1qP5mzWFhIkB5T2AFUsZfX4KXl5isrYzhoPq67E0UjE5Jmh21+NY7apL2MuJHj6FR3
07Rcht+uwWbxlYM5FyXi31pEKQAZsuIMg3vK5onnBgm8rsKERDhsD7S9y9Q44Cip19mmsl0flc22
V7ulfMa0IeeUeNeL/TQeSrl0xcOEXEvTzyZVsne5fU7mIDsMFZHa3bId0y+6mI6vNkGxFtU+RVNj
H37EWSd2hCXrnqvt0Q2KZ/jmmOOSsASCzNizWJW9CovTGEv6ihOL0YVC5lPLIG5T9/aWdhfD1cso
Uy6H2/cfQoy9tZ3NNLqz/8yssDhcDriz+m0b7i6sWTS3IIMtFQYDgEBl04CHkjB9UrHSRh9tUuUj
neduxOnyMVRuBXoRaMtlT2Yl1V1hA1XX1GymAnf0GsNhc6No7BzON96UOf4D3zK4BOupBpCn05pN
onIa46660d23FVQ3CMPtw9RORLIt7yWDNXbO72BjVfm4H1xm8jwkNDKivANpMj8i23BSTIFX/6ss
nGoiCLyQ22YH5ORffo0Rh3EyBzk0jmEQD+TyJvTqJNbbyfjexKl687MURzWJkTx5ShgJHKfNice0
CVFw77ePaCCR+phcHm5AYyDJD/MPAqTk8l5h7bY8lvuig0SFvl8CepgiFP+i5lAvkX9fEHbYqr3K
Y8Uymp/2mRI5VzfnPO7GOmADr4pcSzVRfyNYpe1VjtJc+XJXlWgXH+1GYDPYlqCPjjIXwXKFlp23
mv00uuxjMnEkqkYpN9mRH5ZvvvYgLKHs3AlhbZegLlLulDbIMCPMQgeub0Q5xQGP73JXqZ75rTQH
/Thd1QOnQBNlvd66OOpS8qGiIWCJdxM8FZZn2I+1g3M4OBJ2vmbCiHrCNo9wHI8KnqA8qjIfk33e
fwpxWIEXk00nSFaYV/U1DKeVa6GNn8kbL2giXTSKLIHracDgd8xDU0NzMfDF+Alu+jzeRDTkLsjV
2XVP9McZB4/rdNpU/lwrc0/uwQ8HcCmxJLb/+tca64xwL/gnEYSotPOcgC0tau7qxH0PhKJpUgXI
IS6cPZwMMySEHp9MTDkx7VlpAErmRCO4m8t34y3d7il2Y2GznUUASQDeyFL47sabptEN1PXdg8vo
gucMWVnae4Joj67jJUDKQs/KIgL5aD7SAux60YmMiYvU06Sp51T6YVLR2ALpbtN9xThgVmcJiGw0
Gm7APaL6oJdIYs1LHOMlkxQyczBMcpXl7sMJTRDOgEBTgQTyDva+u0fFndwFqeeKijrlSNPleUW0
d265hoAZZPOsB/3f7cpLPk9588wOhK3+SxBaZLjIIjLJVyJFgrapOuf4gXWtPqO7ijAOofwLD+Wn
5J3RW3x7c6KVdmsulP0LZBaVqlKuWySPS4drFmme71iQADXNzZSSY8U0WVaF7D0tMTIVFTIg9p8u
S+aSH3BimLZTEymP8eFglh7Y5fvtWuh6ryQK0QdM4iJIkMfTmx+KKpFKz71xK++ZOdoOBPU+eZw6
dMAW8KytYblJxFNX26cKhmNDBjzM63lADd0yTTbNe1PWTFFBJ8i6K5+fdzua63/fJKUZIhEDug2g
0DU8vemvGbRXIPOOygYCKJniASmIq6PftZWMMJ3t9Qgdq8MEbtOYXo+IHTjzSn2VZw+txZ3qSKKM
QZqyA/Dtedjy8QZvlego7MGdCGmoZwXQJGXsu0zBJUnAWQFOldcabaW+c6xXZoAXHzZenuJrBdei
Hk2qW3hN+lwRGoUMiUM5hHCIQp9yRAMwjKtk8/pxPvC6xy62KlqZWaP2f7/9y+SqLc2t9NKxRZX+
b0v9zQn1QJHCxb83MGG5XfY4aFGRGfDpRf6s8hh9C9w9bAlNZgGu8mx+rIp0Px0nD/8oAdh9IO0D
1uPcGLYf9JZzZeu8wYOPcjxSPabvZwpc4KWUP0pvgG8EoMRsW9vjIygRoAvKuzhlWMGJ2XZ6i490
hd04ABdR96AaWHkFZjEhZoz65YS/xEK4OvuTq70WI+hCiCrCV0wc9OtX2bG2igqU3GMITowQ66xy
oRfwiTPhiz9CGB82auym1uajYs9owtIuVLHqUUo9bl7R6his6eUahKcFtZYeAG4tkjNi9bszdiPj
LQuMl4OHqz7L1fZe5qVRnOebCJ8Xbw5be2FtQirsDPiqMEGAgzV5XZTGz5JirDTpVohgI64lBMdT
LTIBbb9rioIR7c0Wu554zyE7CD6l8SFQO9gT1OyGG2kkMFui9Xvwr4Lj+d5iedKW1Z4M7jo1ON8a
nhlCSGDGyBGf6BOC1b3PPXGu7YUKhLPwaah/0jnKCVeDDupeRgk3R8jP7M06w+OvUEQI1FpoJg4M
rH6bBpe3ZS+sbh7nco2XiOOOZq0Z6iCoU84HzHvzbB4ZxIQV3FKfsNiJFlvoVbyKM4+Q1sOSabU8
SVvWnuWSNxhPs1Bduw0oigGKzss/f6bKbcupwjfVUR4n03bJmsxsTYCuXpvdgjt6XNZiXnc5eCFa
EMzpXxtuuBztoEQdLUVAkCgxsmwzfLqBiq5Aruho6+DizCzD5pWkRXJdKILpPS8DHfemDLSfzLxg
1PyLhrhZTKIsf+kpnR2thMbQ/tkTG4EtAo6aSZzYcLqmoArDys77rASb/I1TtRnZLx/+v1zaxBnm
wSfhW4u3ujOj1oddePhs84Zg8NbibYV1lPLP0fndLBxkCUwjFRPEraVVgFkFSMIvomondA00Qu9g
KMH/LfmaKXgo6Cv71nA2gTAQ8wF2P7DunzqCbrelNyLmmKtR9+yWWyDbW6VjTasLSjbzZdHvMg6X
hFppmcYiC/yAHGuAZ1gOhUgRbadbX4EeQWtu4DdqbKRAT7TukU/9msBEkIxjm0X3Qa03Y0A6k8NE
bYC18flYwhxm3R1YTehkFozIEMLIeKuNuE0nt51DwJ6gv2nSmOnAenT8KU/Q4s0q2r0BHS3YV2Wl
hq42SZmdn91LRQ+brPGeHFmsxorQr01GmJIgZHfWSGuTZT0qXOYlWqfQML4hPobvd/Jp4l0f9egn
tmvRI+fHUMFZSyrEIhYAc02kgHbiokPx9WYh5ixfHbtctQ0uwGiJ+CY3J+glUdNO+fAOFd3QWVaW
OQfUvlmxGfOD6d3EMieY9KM065k2Bu50ejh0BXm9AlNsr9WPnfhY7Vk07uFtbZukolxYS10NSyNC
tE9WUpLoCzlDxtnuqFyrlnodd7tAC9C+6QfiAyn32TIJyNVX5v0uydHfUJn8+wTmmAhKDLRiC8Dw
eUt+WaVvi7RXK4lVTjXqbC5iWC5rznK838CuK1DM/4kYDg+jyKx0IxxxXlhCoZALShldn7/QwWt5
W9QUKczcLxcwBiEG81reLKa1Owl+m7uaAV5jwCocpp4IItHzG0f3SmcAP7aFi8EnD2Iwqk1UcTsS
/ggZfpDllHmNPwOMnEpE9C0wHBLL/+dVh7d+NVODf+UjjnEhTeJYHTUYVoRT1Gb9snmmhKQkdG1B
/XQBGhnwL6R7SKF7DdRcWmpxkfgJu+RC8CBRvP7AvGbt7yNgDHtpq6Z7CLH1ARoeg1NWSnIaOXPv
RLd5QqVwZxR4YIjYyNi/ioke6NjbKF896t4YmxMPW1nRjb29rX5iL/UNNZQ+FPk1HpuCSr7b4vrX
P3geg6xIoUsnAcjNNPtQg84qxunTaKE2LeB1fcPhmzWNW9sgHRxYKW0rsosOR+NIDdE8T2bmtjF2
BQ63xdEOPSRB8cceB4RuBYH8rrRzbI/4OPwu5ydfDaFKTLCdXBwJyUr6r7skab0rcy5O3Qk/Wr6a
eKnl0TQsy+fn6FD8ZLvFTW7ANdoPbwvLGlMmG/7IFPsaM+1hXFT+lHhP7Ox+yYKZFGmKqZYDtO4J
5tj9rnh0fwMg6H3V+UALZzVTt5wLyTYpXJ9R0Of2Wsw+urymEu9AOp6LLqJ9N+iMZGiCduL7Icf9
6nD7uu3E+2a0xvL+6hQs0rsPMP+nnwlHQov/NT+1bwceXImLrCEkRUAkA9skQgUuWt/r08tIMj9k
YWo4NJlNeEHoRWZoPAKCGgKUvw7Zoyo/qfrYcp8lzQI5krcbcmpDaFwjDY5xA9vpbkA+a9uVoMB9
9hU+1pk8g5eLdQYuzAj2j3UapoTtOhxyH9qwH21yORyfuV7Bp+9B4vE48BBJ25Am6EvSxMhgC6sJ
mUPkq8Jr0eaRl57VL1rqb2PXJJvAZJmGsqSzhhnT5YbQWG9nRSAKzavCvSEL6TGomkDxZzVdjdt2
JBYWMW9roNfu4OlDxsS/Qm6RD1QtBIv0auyWw0axrhW37p+gDbFyfITBphkfzrRbj8OdKcx9JDhw
qAULzFaTjFCJBRg6UglIWd9nHttzvIqfkiDDf29euG5Py8WxZ706SH7IEm7VEP1eVMZfaOP4RTmw
7SJCjg5U43gVF/wlwgqH+Cwmj9QStDHBOF8joafAwrWa0PKjJXktUYethlPgAt1bZ2QFl1xe9MFP
aMx+xIs2DHHF4KR5OHKHSxDKZGUf2zebyZ0FhRpelIizZk7DqOIlWVKtiyXUVKMiDN4YTcfGfKI3
G5JFIa7msVnQSWuf0jhsnc/aY/RFGvIVpQ7a7DvLOIwbvr3sdJqtIP419u4p/GeIxws+8moWrm12
nguNlQ7/EaSjZ0ZZ2kXMkH0m1CYVqhJgcyaPW1sOp+witcIiTp0bSVARmBQAXrpTUNrpITh2VxM8
yevVwhJST2aXeWRoogBVegj5CzBSp7qVtrW7S9EBZST/2M71Q0yu6JnnA6nAOLZF425Rec4TtrTa
IW4wWpGnhyUt/3+SGe8JgbunZPVo8xWnyXovwOlczh+YtV+RKJdIZ9zMEMEXnELRbdzJGgcAGGlh
Zsrq+RRZR31K3MX+sXt3cyevGRFlpm7EJwClKqamfoK+zVyKe2JTrWXe4JnJ/p5xrEa6F75MZL3P
LmJzapV4UlqDE68jFkiXKdOEMBOwAYy25Lx+ult9zoLTSiaoZ5m87rHQVFSVUOgsOldw11fXTzuZ
Chnb4L3V6PB6TdQftiNN8vEtXM8JtmEnqqgsx0kic7BPs+jPi/5uKQ25wa8tz7W9f5MIrrprZRA3
OjRxpqxOzy9wluiGWZ8z7gp1uVrnWTV1jnf/9p06DX53G0CuvAR3BH9S9dEIV4PGD6ALFr1o+pXm
c1rP/aKBqriDd81e81ygvtFjJwP4ENKRDyQ95zgJGfGJA1TE3zziRB1dhkqFAneSCi6vFs3u/N6x
SUbD39Th7bOUeqgXYR/1IkB6upQMqnOdzJyDlbyaX8IRov1xQ8yPN9kj4VKEdYJIwFUDThEYLkwF
j8deMNnXzp8z33fOH3gQN6Vl/x1Yt8uSEyx7VumfD8uuBuWOVBf9eUdfVZOCfUGtYsxMQo1rsc/e
SONHS7P6InBJy3HSS2T/VWsvAJVrREExa9jLxcF1ycegovQiTTw1+gx37dE352TSbRnY5GPJfm0E
3zWlA2pNhDxSDNjfqB8XsEfzqexUhmJexl4Kl0s3IImn+RFxZhWLutUv1kujVfKg/2J2MRlVfFyd
FFzj10bkdWvo7T0IW8rdNSH1UF1WyvKXUwPlowtSnDW/4pzBCXSnxf6/WL5ZI2KPiY1Igwu316Is
kEJkGSBW8EOQ52Edl/lGO5flu6vR3YAqyF59qIn3nXpbIdp7ni5uvemrM9QlIxye19jSSsp+KE4p
E6vtQpOvSz0HSqQGSq9a2hKTv0DVQNeBSF7x/DL8UEFfLhgRjZRy19dZ71p9tK9UeuggDNlI0Jqf
/yIRcAXx9Sc4cNoa0moxKgVhB++ioN9bBPKpSRwmGM/I547KaAzw+npDXnns+tnmaruISLdknB+k
asgO20PUvLNXBLBRrhDLn6BabwHx+YgOqsbsOGZP7PB0boAh0/IjlCi2TxSW/g7CWmR6XCCa4d1I
LOTQwOdbs4mMHSTOwqxkjQ8EST6mJrfIJNCL1oQoOTAoBkvxRBxOx1CJ2cae+orGimUVKgbo+PdD
QVrNHw9HA9kJa1SRPQXyR0ho3Bi+64nLr2BMKOgHwbo6F0A63uhaQaDzcnWg7Fog1igG2UOgqKFs
fMgFm1UejN8CIOiX4oab1WJT4HuAEyRgA5zX11E94ehMIXbwoxGPU48ze8x7u9f3w5HyDEbeeAtY
SRNHDAMFtvt4h0GDz2Bpu/BgUcBZBFX25xQ1DWURIyrNLbH6iyfZ1uJ4fa8KlSKiFbrX7E2dYPsc
gTrOg6BUfH9A+V3CxC1VI1vppNaHR2F5XpgOUHWM+oQYBGi7To74H0kHonCpPTCimRX+gmBpDD/V
o9bY/xuwuu3XG6KoWUhpFoBFPrpxnQUaWnO5dkTtHsBDZODyIRq6Zd7cvstYgFJ9hk847iMqVsuR
l700XkFE8mMLXvSHpoia7vSWSKOMNv+dx2XmdShuIhFxhJUlUqIvmr+LxR0nVr7FewqVFxMLhINC
Ch49TgYuzNQaAEWk8HZZ3F1sdZyMsaWihX8BpqVVkTuy4CSmkN2CQdsy5PDHpYWiApANABEVmwk1
tfH3hT5MeeDJ2xeDIkpMhhiafQwPeO5dStO8gwGLZKP6kjrlkQlFD3XWDpAN8+xYK7J4YgJglLaQ
wESLTH83TskHmpVsgu6aiU2qMWrNp4G15GoAa3K0nKR5R7BKVkBet/+ZzUTs7C4ue9J869tRHDut
zxLbDYsMCda0PpoRPNY6P0pxxQyuxdHIuPbEqc72ooovCXZuTHKHReSLgifmTsNTvyNK6NkJicrD
LOJC2Z3uDNSKM5dYLE4Xp6ABiOApqGPWZdrsPAaISvOTTYCdMIixed4RLN4u88+gMJy0wgJ7SyPu
pie++3bdnF5GssGIj9uanGzD8DkbJwIY43T2pFtiH4tWVhMExGziMGn/IkIau3SlkLJoxDSeTnLJ
+8Ii9c1zU1ATZ2jLCMy6LvuspNmZf/8LtH+6ypLRN7YK8uf+tEb7csjJAZM9gLXrFx+pFTjJnl+c
WpwDB0A01vx5I2j44c8mZmkh+ThMTlNFxzq/CF1MMBtrZRjZ34P15/w+w6EoP4ZT6eqjUvQti7LA
6+9A7A9QnOQl6fYzJ1odBQ/CszSrWFcMBynx7Dyncr+qLRTPJR44oAOHJmTs4PDXtTExYAjRgsfw
inP6oaZ+2iAQ40ovljAj0DarrS+xYbom4pD3VY+pnLIMw7Qeo28uUw7f46ogzhSh3RQYRQHTolMt
mFAEVPq4wJmwuOYaDiybhCqcXJj2420Z/EMoaVUyM4w19XYIPnXJgL+cj9C8I0aUwxXCuv7dJVc/
efHFWZg90AI+qyM54b0qJ4mms8dI0vrpeakZ5WKzmXdqIrwKuLVVbTqwcFNNGGIpONjtyK+Xnuie
ogNvTxPsLhuSjdHebcVd99i+s8oXJPYqk9Rwt8fXogTLxBep2Yt7Xn2KSRXV7+5mOR3UAaxOEu0S
yhAlQL9VPgyl9+TbEKQgINe6RbMypnO0sdcV85ADdboGvvm0SbMb/sWOxOrV8UxhIDaT+VkSjz5s
1Js7YcOYJUhI+dZWKKgVY2UgOc2nJXpoCDNXtb7KRJdvtBubmaSeasTbMiCyclIktDNOT/lpSP0+
wLJF+KYtmyE/HY4whMO0+B1gpXnbVCdgMODfmkIeNAhJUIR0B7DrE63JXcCqaj8D/6Uom5QuuSnV
FLtSKqAGDKiDMkdJTOgPl0PyxHlgDfAfY50/Vj2+Mu/XbETAUgV726EufcQ79f6LUe65luLEZ01l
5NwxcVPQq+WeowCoEakoWCATz8u0hOlqZw68Zw7GvRj/AkTL56vevKoMdPzQrS4vXCXRMJX6MF71
4i0DWR5TsHnoYyW8o50GoP4VsO2O9o8yBdsZgt52fv8HWuUoGPxyNoJyRDTe/f8adOKyn9rGEUih
qy8FbBJLFJ5g4804infUlwnlvafc90pdglI0mb8SIy2n0ePgyfZwIRimjHVJ6oyUO6BYwsU8nRQC
fYmF5LYW6NGWyVsUfmVXx5VMn63gTVrFGLk0tVUGx9tK7t83i/UoErhBiC11wItbf7iaL6zauti3
xJ4oenGWDcnXAXBrFNzP3aGJkqvZ+hu+jwwZJGDx8zu0z5R8SOP4JBpvJJmo1bKpS2tK8aE7+EZk
eFOjgN9swvWAfkbmGgG8INQ+AEyJ5LYg7Fb3aIYgDVggTlXlwGzhXCCkZat27hgWCizr7tcJjWVJ
AFzkJmQCPpmlCC+VbIYAYznxjKLqyzHvroPKnEdWNMNEuQMwDCNk4P/q/uW+rdXiGsAQypka/ile
u+Z6a3WQtoQun3o3VKRXMaAVosv1ktowGqVai47Y2AS6Pf7izo8t0yIC4m23OMppGmHxjpKeHGy+
wdGtbbAy+Czz6iq7KwNHE3RnAiL9mrJghNwk/yLhMpsEnMQCeWBQjUWph6RfLWjqW2EDaqDV+WyC
clD7LDqxo4NvcBFWaPDQq/XKTrxMzij+eH6fcr9vTCBb31zuRbEzE+UaPFc40yd+zLabvRVoGM66
JCbBN/mmDwtKs/sLfCxnSJBFT4hfrS3cRBSuCB9RsZ7nFTafBmo1OTFkp8HXCOuYHvLCcFrxHd8W
aZ+a8T0ZltvfegRUO21bFEnJXfuDOPevt6+uPOwsa7iKwaqh+EoUjjWuIhk57QCvWl2QxLR6xh6d
VYMpbDp47YdoMptMwVJ4dtlHjIRHZaUgw4FmuOZJGNB67i4M9Hu0dw7P6ecmyX1U6CzS8IV1dMn4
uSsM8bcaQWU+L798eMOZa6BULhLCA44TT061VD5MiRe4QYnzcbT3OZAeEa5SRQszSTbAh3Bx0mW7
4nAVylvojR/TJmmXG/HmWTadMv9tVKJ7c9ODTcta6p3qXIrZT8ylwJ7ycBd8h5BqPow6GmewC/Lt
ajw15CoJa12dshjzxD3bdzFLgURYCovPPsqEDje+aYuu52y9Sx91YRq7macL9j3I4+KNiNgnwJJE
S7J6xHNsekQN0dczVsNrhGCQBPiuLERZjhJxSfVHIg5+rkg0yijgqBrauELG8m2Y7eSN+Ex72Pic
WW2gGfawj+56IEWYKOO1etS9Ts8cXZDFqtrwauQSoVNbEisX/XXpP8zIEZR2CLE6PDW+Di63Betz
SSJBZW61o2uDC0AcXlMPLbxy+NAXAJfYVZtsK0HLJ7oKtkgEBSuHKCneVuNO3wpM8gd8OvpTf4dz
zYx4Gf2RkEwxV15VgptVZvAszqdHc/lkABmFkvr/XGOatdVgCiZAo3030+AC+15hxzNr/S+xgWdd
GdhuBzBL/J3a6ixGP2uTYsIu+NnwINvrSHTxdQxcShFcYiiFf3hyT0muBMAmOsuBQZJ9HNAPt/f8
9gnyeijySZIUW2Mae/JByQ081NIgXWPbE9CRNX7oKL/7frKyQsCkDVE0g9TuPdNw7mEisWMZbkLd
JxtTjvTqRC6wX3tEVV1KBXfLGQInv0JURJUDN2fMXwaB9msQElvrypqvN5UzPB28NSQf1lhHCrut
88fxwjmboq6AzlPP+GhLnh+BUbPUtm1BvXANk3GmpqQCNr4ZM6mHHCW5D91WletcM84YePQ38dC7
G1/RBqlQVCITD9W2RtnppFoWAAH4/JHvUFCdk12Q6o7Gmvs3Y7EwqgIFcHvm9xhIjk+kpAY1EX62
ydqMVOSNadEwPLXWrwoGS0UAWpCKRNtP5rChvLVuApe2lhz0WgQ5GDfpAInaYzfrvyuIB3wHRHqJ
ivc2/cJJMlMnKM3omTTLBRqOfNVUA7gxZ2oHXwnjLvEAx1oSoMEAW56ZJqMQ8tPd0OevdTmimODU
T+wDKIqtQz+b6tQh4RTmhoaERVybdT3fMzKokuNmhJCGD8Tko6Dp6oIhUuR1o+nTcHbEUZ7wd+st
XstgXR9m7caC6aiquVbXSdVnjUf97IFvK2tGSfUtNbzPcyFoojn2bKJQ37t2w03LDgiqJZqgY2RZ
u5/0B0EsBpvtNSiInz5CW1K7MUou+BDuoP4DnJRyDZk/gxHADUlaDP5gIbqD3xIsAjHHRDqR74YC
qKHui0gtoRNCazuB6hqJglF8wsm97pMiLaC/aME6abi9MM84/lQfnuAUEJ25QZMS5KvhnFZOunrL
Jo3fQl4AiFUH1uJGD37tiO3wcj/AUVm8ijgiNS0TObyhNH0B1lQDoJttvpMDNEDACYdYM6Ugf/PT
Euf90hNxmPS6VWZzD+qx6NlZAfp1+DLPK7OSysHbuTH5sbOQ6onCTXiNRL8Pqpj+mQZJw/qq8uKH
8vDUlSkMiSxw7uEd5ASSSEaq+AaxtZtpS7U7oQK4XIPcBCuPAKz/glFTGiT7C9n/V1HkH3waMliB
/VfjpXMgzbo/1YBEk4wncD1H48yMxqIe8mnLCuOGfVbzWbGhTcACzEw5WP3fSzzJ3xGF4csm01kV
4LVYm5G95lqZjA9/fVHT1PoiYEX6VCBJ1urvziJdQ6k3qXRcNpFT3wSxlm+qytMbBOw8F0HvAfK7
3aLmshO9wGAJkOwChYIlZjucuzQSnAJmXXtGlHL5DMec4qK59eaKxp2TV2hqjI506ca7q+4KRdaw
5MyIRn3mSoPNLSq1dtM6zmphRQT8myFUcNT/lUtpMJ8TiTw7ER//N2/kibqDK86Et7ZC/LDbWBDz
LGi7ZjIzw1/LQK4ppIfJ9hLC3nN2iYv4YHyQDrR2tzyRKoHfP3VXLBq8MbA11Nd57aj22kVPQgD0
c5d66LMjdhy0DDfPuRzUGnJ36ATEuoLSoV6ZJXQPQKCV+C4W/9dasUFtCUIPRPgh52naEostBx1Z
Iv4+cwuoW6odS0cvsReVOp7JKN7FLk81giwDznG3YI0oDYqvijfsgB2tZ8bFSMZJPQQuKhNTIZMI
xlNbBe6QScANwteE7iRoxZmrDDC85u+Ws3zYEKCMvAvK10Up+8Gc+3RLFI+Nax/ciscdR84aqhEt
KOWxn9JG9IX9HcmfMfnvrDZpFyvmwJ5HIX5VhTMU+AAoqGUWCv6J05pYwXZHHmgvoaTgUXlNBO0I
EerOEFfbBK6P0c+f3UyQ/G7nP10xVotQdXOtVI8iET/Qb3F55jIOSFHfk1QE1TRae5s8C2qeO6ei
KxlCBrWYwfY85fyDDEt10Oz0GT98p66aZSO1HjNLRUsgw4uiwuR0od7Hqzn2M+0jZTk9Abs5HaOV
1ACALKVslhgSVbgo0MxxZ0u4Zx5DlSI6JSR4DXLVxRrmW9Ta/wJbvlOHlqUnS5zFeW0baRM31BLN
0y8pb+uTzOqrCz9DZP7fc6OtvJFxCcbs8hA/zSWc9oefmM9ZyHQEa2GGqo6DvWH0516f3NpXz4eM
m25vgAur6/6WD/5v7I9hACc85O7wF5v3S76Syn4yQrsEXV9WCQRSWqXEexStO7SDcfpxIs2JpaT6
0meYe6/vMRDG/5I7NrXSL2CxZMA8dcaYI+CO8i+dtxowe1KrELNTtta1odUKXPGsKqrFS4qoBtl5
ae7wXFFC1swaZUwShz3gEj1B5MDZJROaXo4Ybr8nHRs1QvWOVlEsRrZOKNxeWOfTwje5C+sO5UaM
akpGOFS42aUa9V2pke5zbPoKoU4f0Y3tQa2p5WPgWc4Ih5xLWfywSLqzJ11OLW4xgWqYlqlvtyxa
3PAMw+T7BBF0SNQKBt4Pj4Iotbk+lXGFTuoNLX2YK7bzjr23cJfalUht5Fw4iwbH1pRCZYpAMrg0
uxDBUaaBHggeiTAc61/WnsvrXYfXy7GS+TT62zllbqPDThPcZVJNO2q+RD5XQXEslTT+HaytmUzb
Ted0rbECC8OZPk0IIpVuvy9gR+08Z+FTZ8eLt4ih0+dl8i245uGrbB356TFC3ZgsCS9Pf3/+8s7v
l/8SG5Ol4nG/g0yg0Us+FOacAbjhT37eo0L7fHmUW0mbGpPqD7pfdzis9cBJgdrhaqQdbOqSRDUp
nIhRz+Pfxy7SfB8aZF9Of7vnCB9x3cGlpCnbfIsBFcnaZGoBumnHfRbOv3AjoK1dYkY8kBDy4wLQ
sfvx1qCGGkwOoIH0jY6En8IttYDEXWkZh2fUKpdmzcf4eLnoAmbgFjSPUxMmb9yFumK8gf4JYA9v
CODcGj3ONUE05dKxVyXpzBBuADug+7FO4WRRfiZObxkm8iQEyG+Dq96tJkfLPOp94+8c7l3fjU7H
0RrMzMCPXiHY7jI9LvEyWB3fmEAEX8pdetMCdUw3zqXpWdFWZnyeQ6hVNBoCKd7DtAYHJnPOUqrP
JVHmH/AzPmg4ar2pbOJ+gRxuKruYKlJG52A+4RaQHBuP4Gj6FGp5+qmQBjurzBxbLrzm6wYDKfdB
BJjNtrqYOh4zgtTucIrh0ypN/k9hXlXFncA19pPu/rwjdBXlDgA/LKeAycszuqPoXdbceMrr0e9i
OY6s2wI6oSAxEkLvdRPtMfp+YHzHrLbSvOEdOwwkUn8HOWKvQykAv0okHHLDt6LysvclTf/Dx4iO
pwekCm2fVUKBBF0GcWjTtW4y2DAA53iiGdueOlf0vCDU7RRPQN8OGSQvSyjM7npxP2LqKM9eO078
fLMFM2zNxg94lQWTA2VEdmQWrFJrDDZiUqGwM/sdBiK883tCzKovZZHp1A8zoN6VqOr5UtyDAYZU
Y36RTyqGaywPOmjoGQhJ4Oo4oXiBElrZzuN2wmgSCy7yN2X35CYPIUZo8cpfoYJyhc774tTEtSB8
auTd9GfWECLanJmqAI6kKjJHhlJhJ0ZsQBP4ON4lmi+wtiNKoXElo88juQWsD0vg8Am5VkjLoVV+
k5K1kmAzkmc5mmcgB/wwH/ABXz1g8tzB8pxYbilXs+aG954sknt6Rl+aRm/cYIqAK83Hl1nqoAZu
jq3L/MjXZC8ysQdp0CMWCNvv9C0Fu9FFgDlG5TlCPsfYWqN9VKyPn3yrbXpUsYlTGL7Anxm7c8Lm
7YeQorckzakCU+mSxNvdP6U0CQVCHnI1KX4U2sjYcWYb60rBTds22yaF4uP5MJwS+AgUr/+txUBX
RuvnLirlqEBdcoo1IHKhiTREVm1CffoKArS/CTQoi7DjOfGbJztObGOfqNVT3ffBtq2ff3TZiZU0
JkfXiDFBRpHtLE2qM8fvWtSW0mYySsN51G28mCVDZeln7g1KOgob6TcnsuJa0HQf38L+EOXO3h4A
Jw==
`protect end_protected
