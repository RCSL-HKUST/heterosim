`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fM08+zS5HtZ++cY+GqlLBCBvOsyndHZb3YC5pf0nypntAOhY/euJaEsYqBntNIyD8ExqjRu+qk4A7KBwHItLTA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f4W0yX7oIh4ZZaOqnIhhXrgjDvlqWcoagDaRAd9fUeLdn1mnGathj0sWfiKqaIoHusebpoFdXg6qTMp8MGvUZCztIAnBQ7XpweahmdwAgBacni+SudUkPsKurh0p/EpsX5Y33dn61g51yJ6YD+H1MHOde3zGo4cDfa+a3+lKeLo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xvi7DI+uGiLJKaEAHy5pRnBCkW2jMRJsaR0WAF6iRTQAt/kepq4OYhlo+HJwymu27E2+k1voA2/oSDP7hgg9KZRXzbI9nuRZxmrKQAJfOiCXphP5w8tjm2tkEODeB05pXlZIVUvmU+FLTyXmd62CGrzUSJx+yZDaht5w5pGlvt1corTMqv/B8ZUedMl7KrP7BDY5SGyZ7e60cxSYFoiDEUlo1/Bbw5KXoPebjo3GQ+ZdTzsAqYMFqN9FKg5dnVV1k5WnzZ4RcdmjwFcW8zCoXy1TsdpjmazPfq2LMtmQvR6ts7dUd5XGMRZ+9mr1QbzWGoClRWwlgp8Uiswlxdn0+w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N/HgrXycqnR4WnVbLERsQ6abHWIZhclHAzrpb8NS7z2+DeAtp5/+akQwLfrGsEzNAJU33iQjsWCQfGZn1qjKvfPsgmVsQ5xDIKLt7fv7hbe+Eq6UWqTm/fSOgHY+yWtNyLWQTiOJCoxdR7RD0WLsQ0TGBKLySft7P21vd6qozmk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gLiCrsuk9VOADqW2Mg9YA9LOzN55cL/sG9r/8aTY/DaRhgzN/4jpD9vOT0b/TrWWnE9QGRssQyA3L2UXoULKs6wLyN5KAOhy/et9udrKBGXmJ6lL7nyqip0VItsPn9945fI7/i+OOnDCHUq7hvKPXw3n8LwgRV5YDnqTKwNqkLj4sFpNlaPnKHWvRSJkAI3QAxxAcVAvUdVxWK9rk8CinXiB0KG/iBmPvdXx/ibLSTSjoGUy2aGtWYnTGY9v3z2xUCnFRIOdO0zn+p5iVJtEvyVQV0we3oS0R/KSO+CJwY8JHEZnQN+aNv8dm6Q67KgZQxi3IEzRcnrUEqZz6yIcIg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 117293)
`protect data_block
qv4I2PA+AwYJLS2RmDOIOAoQ04dnwlq5/tsutbJzB/qs3V9c359Hh8jXsFFuJwwHBGYW3TA8f6Yj
dvB7iHhsTPzeb5eKiQPriBbfxmGPEIPq8DLEr0EHG5IkEXakVVXWcyORdXlle4e4X1EKVaX1mQRm
mmK5QPZxuiT1U1PXm3+0oOrVHi/XdVDpDhDU7ziSm/9x6SA9ixYFwc9nZNQmLKWNeI46IIMZLz59
Fp5Xa2w/G+2lJvI8rSIOFiEYHtX+b+w8W9EQEkXfoa1i/LKv1aLsYqgqf2niNXBQODC6dJ7d1a60
GT+IsptTSSQxxIlblSYoKBxICAfDxkWxz2BTv/rGtazX9siJJ6dRiutHjJ7eeMXaaLBkH04G/Mcp
PQKoCowsMsYfRb/Q+eLLydDNGNBqtI5jdpcJxsmZ6ze4jy1qvQvVsgLFz1tFS3PTsohKv42gZ2UO
kzOy4XqT7zDoXZPG7W73PoQc5/npgC6PILDMCmgsr9+jrWe0btdbjLWwTV0fYAdEeSbSL9oqkQi5
jOpEKiKGJkRSOVfL44SjfNMJ78y09LxlauxH4rXflJj8G4Y5+btKHOVj8ig6zRqX2+5eeNSr/4lZ
Lj0hfk+MA5IXa48DNSi9ZUHMu9U2RpJw4EFZvqoy/SlC5UAZiKoYPJviKJnNrzkzfeZwSx6sAZDA
oFtEC7OZnwfVvKifKgsJhOYY0yx15soBuO4L1IAXbjN1pGchZ20gi4ZnD9KBU34EoUg7HDKDh9dH
kwvpVnVNweptOwuzbV+VS6fFtRA5Yli7OpBEFtN96PO5+9YhyiDDjJm4Lku+nMu8usbUw3kgmn8b
ttaCL99erPR/7pfjDmki/PrUv1m4SOLUL+yR3/ChFrgscBcElXMsRFoB5g0E4nqAqWyd772pUwzn
yzcBVPRuHCTL1o3DOY5OiHRSOZSedehO3ooY8MpDBBZwjtNgzsv0y2rmAb/Bl+1zKLVCM3XCuA1x
bI3Dw9KjD57P1G41kP6uOiUc1I8Trx7LX4wpHXuGUYvUHuKIRFhUFw3W23PSa3EX9f6TtFlC0F50
dUzniaxUZX5CDYeLpYpX+2kItbJy05NnPZmqTZ7+9ccVK26m2cO0Py+vN+xgvIOzVVxHJ2bHNQPr
ycY6UQvqkPBgx/7mkdFsN3gYq/LT6zG8jfBj3SeqENck4gC6RN+SeSYgMFjnnCnfyIVH4M9iUclz
aGiHFZOMBLZFkkHbG8WvENvICl5cCJFoubaoYgQA6O2XCi9t08hX/9Vvog6dWeORHkPasJm7+CUC
4hci9K59KIgfZ2jpE7rJp+jla4+Qbk9d+RDj6fAYlZU8sAlZ/7US0A3w/sw5Dr1Be+hPjudkPSgP
Lpvx+CAL6zXJlQJ4gOsNAQqxmIMbbMR7BCgH+W4OhIBr46C+awZhrRg2OA+mMQ3zU09rvogmWqQp
TJU36FhJvKrVYPM6lQMGVRCIR5vEfbTTahQEngPLZUdH+/Lm1gzEcmK+BjlF4xXh2TuAxc7YWrRm
zoLkCQww+02n501C1h0ceir63Uu82EhAbsRWAgiZbojcXagAfA9fY56YJyw7fNyKWLkFbsyd5eJO
ni+/Ppdv6VZQfchR+DuXmAY8/8t4x/p9pG9aY/n6+y6CBTWgQeLUcrdaca7f3WT6D2/Q4ICgA4xf
QhXNOKvrCSHDqmYDZ0q5JalH9EhuN95lvpBOkX/2x1eIkrBonciKJqDQ6PDMr+spGS9jEF1hMckL
PtRR5zL98Y7X9jU8aXjimBMt8hu1ZCkZV+m8us6/S7Wo1tgwJTBA9ZTLzcJGOCgYZZQVupy4Jr9+
+FdRyyLYxuWCW8Wf8znB2jIoqT2Y1WswzJGzY7hXqhqaJCD9F7ftz5T3/NieQhic2PhrQiIMr0Mf
gq/U8yUxcIfEmbkddSMT6WWRDVzLh77vxS+L/Eotc9pvaEr/0HsAW0tf7F8eyfJRaLPwEj4nHid2
Sv8wpDLSMn/vhFzyC9QpRYOsH0ys1H5RnnaBWaqqy1a8u1rsPhvq/3DQdpDPAupyixQZ3APf9ztX
uyJglkam+qssLVVbTCmh/SkV4ZhyksepVzFVio09eRbUYgYGE9Q0cmycHNSymelNX+ruzEg+9NzO
E2kXuPCGg/+9idQfjuBkWEiRhWb49jH1rWc+TSiE44IxGCmNlHGjAbCEKfi6+YEIiLTk2ShXoVd8
FO+bkxYnQQq4fgjzXlNWrhjRDxNsNcZD2Q0n8bxd1nIPoUOELK3jm5UEHRKWohwL0HgVPK6jRbu/
0vOUzIc1uFJvgBiCHpxcR3PbeJTMpRG9clvrzJcslZh0rEKRW3RredmW1fKDhGT/ZecadNLI9rzd
dB75xFBdQw9+AoFYeMFKUsXLlr8tj9LAf6n3iTvR3fgYGtB/Qz7XsDtHs+taEIQcsxtMEWxmJKhx
eVVk7ssj8YXTEUmA2zSldoAuTFWcceoJmetdvK6p/Qga6pVzbDdtTmGj+mZlyUW6MfxCQhK2ydf1
X2Vq5l+O0uTGG+xDwObAL2jDa0EZCAI5QtVbSNvp4qUAZVE+TXL0aCYqKl2/mfJvIccuoRF/tyXI
FrEVHlg8YOUtelSdvXy4wU8c0C2T9DMmzquZpeFjiq6rgnHsp0JckAczKcLqzfgPHmRY9wJ+RTYH
dzphJKrihi/mS7Hc9m4zjRg/GPDXP0/O/QvMDc8xAQZrBULTSp/hVY3GVoe9y9KObENnHsL+oegs
CntDhBSANPjpn9plYXFBfbj6eSBTXvS/jcGLf/P3R63orl9QYI1EYU0XAojGN15SPyN0vMcP1yft
73/fQwoSMlEC4s/zA9+WnvT5toV4Lb1aLN6I2ARfKoM2sb9+nEg6jbK4ECdYzYSdVrfCjwdCT5E6
sb4XgrXgxFxioJIQhcmWnRFhza8BjvZvACl+OKArCgiMuWOP7gTDZZfihgqoaEjrBXO+MJmQpRzH
M4f3W39dJA4YoA3gZz3KZScRReF1izXPlNsEOZtj+CKIv+P7EfNtT4PWdvhWXpUYzob/kIHRoGpg
65Ila49PNTRx+B9oPL7RPcqWYpMU0/HwkS7fNjZz3R27vQ/i+IdhkFcXc0g+fufMT3JrKQFvwvoQ
su97lbW68XvEY4ttiEYWnBhQGOI9W2lWIn1WaYW/88hF3ahwX0Q6PQdWiQVaXSRplzIoqX37T+EJ
wzN7NQj628A9KE39on8NQXr35qqxxW3NHi9WZF8mfBpDhZzXY50LFfLyHR0emkvHLp5vIwfbYJ2n
KAd2UTaHsIGnpaoNwtZl2CScF66GItaAk+4PkshPki3JPlKDJJS2N/E2tLWwewqI5PdaZaAZjccd
4Ck1bom8tYB7Yxtd8bgm4RZDbvc/IlP9+YGT2vgKx4N8mm3qfJa4JQTe8meutQ6u70rgGuggJxRu
L3BOixAg8NamK+xyGNOQBs/qqCkQ0nJDjxHzyl8PDrqAe0dEv2bYPvOzO/9eGrvjfB1WPMkC2vvr
qYtm4nMDw1/nccJ6IIAxJ3iOtgMsVyy7rqLVLBw+UGKGUhX4wdrluB+HmjNDj8J0xoYSHguDCnqp
bP2XUG3Z7TZQJjO/wcvCrf6I3EddS+K3tfIsmBkjoI8jMeOVvGrZRNSAuLKuwGj7JKKH44XH8Xh0
SqtJds7tFQg8v4nzTkCQP29Cjx45RowSkNdHNh4Dc7/q78LliCuzX+8rQ3IxhtxCz0K/aAH3OO+P
CDXVqBq5ejVz0+NavzAjtjF+URJ2Ar9aajV1gN5Fc5vB3fNYDkUm4Umj7mDwgB5lTDdQJwXRk6UK
huIEBPOmoFrU1B6pdUIO79BrThofWw5JykD3jrUqFJ+ypHWU0IQ2rTeR8joOzMf0K1WuQDdB8Bz1
/HGbEPtLvtZu3Eos+mIxCKCFwmgVx7mQQSN24h5jAuC6ZgirCNg/MBNd+QRECvZsiGG67KRn6/ma
9DasCMDS/nm9k6zmzd5HoFgUkaUxFXhfTaaVPsmUxwG5eeTd+Oh/wES7rcpPx6JIWFYBauwC/24f
V91E9tdPvozRt2xiGK6uJhgRz6zYo1ay/wfxxaeami29JA9x0R+YeI25PPAeQXC83mlKpkoJtCY+
GOVc6/iJcYOJTS59HRo2KtA4oFpBf0N7cOj52icxkMC9x2BgbGFgf5JO0KR+ZzfLs0xWalNd5E3p
VD6J9mOTpwtUQSubGouhUubQ4Y4mcgvsP1+iKZs0kQGvSHCF+8MdWcoFmvGZ/77q2ML+kSTVJrj4
P45v+TyEuEu9mSTdUysaCVqrvfvaP50nt7Ey9qDTUGjFGrKgGlKNtoiUqkBbs68Lc2dYXs2MwSpO
ygLgkbMaaEXOQDxY36liNO287KpLkPcnjt9Ylrb1M07ZqBX4iIKklBiCDLie3qdbzNpwQkQiSptd
WjPVpLBvkZVJmR5ih35qWaCpy6bvj1TVnkHUR8UzgifCpjCk3a9D5WkK4md2lm4z6nyhmfz1ajXb
6vmn8gNfcUYPQFz7q5mdlDlZt9U1j+0jZaTjVuHPqttuKp7EUojIahez7vgwU13kuFixe3h9c1bg
aNgFzD1KQwDZGRK2RB6z1mdk4b6KIQfNwR96bg79V8wtzuIb3YOHZ3BCG8ECXhautiZPcUHvxtlt
LdvC2utcP1cAmFKN71MfTnvDKBjmqKPGsOaSRKH3nBmff1TpKIsLH1wLHxJ4zFgsje3215P1k5Gr
yBN73pYMEOz3OolLNJm1k7vcUtm3w6H7wA3XhdzHpYuHF9mvu7HgUQehUGYOus/TWqQrcaf76kBo
iG7fcpha+krbwyTHI+nPF7CHnzkEkNOCpTYwIcUWBcY5kk3Aw863oR1/qoeE8bJ3WFVVQeQBdN6W
9YgG0l0n9pzISTj9xfwPqPxfFSM8RmXXixs+DgIpOCxE2tznHayQ3JFNfsbtwdrS4ja1+/ErPvnV
xhER8/D9PhqJNkCz6T5NikgMtWH+Fm92JRtswiUIfYHZ/6eUI6CdgdxBqrdaoY+TnWwRDNhGm9Sv
OUHGVgCppaTmLv1OF++q+4FRjE9kGe44AW+dYk+wqOwZD4gWbXJGqviKF4a0RRO5ujV7+uvqgjV9
PatV5+oMGxX2mX04IdxRzrpcwX+aflJ52jiMoEvCxpe0abahUvx3sBzqJANrLdsXnEVP+M7UhlCe
GmxAHu5Z1pet4vUvWDUD6jEI/lW09Hyzj2vvRsaFt8DOlygOW2RZDdG7DW/bOP5weAWOWmGjaZGh
qyXcXFVmIIfBvisH7vOBVI31sWh5oOgnxi50sW9AfV5bLfsuE3QTbBWoz7GtbpmqUso7oemF95Kp
bzt+FCScZDQ+ejzYYepL2Ccr0RbdFnfpefHCwwHpaEyKAN0ohbsy9r4wIlJ2Pltnb/6jIdlEN0OJ
Rkmw05u+wCfqlp32iPP9OK/qQulzCdjpA7g765+RbaVelXu9eKALOe2l0ddiurPdW44lDCea3iEg
/F5A6sJLU9KyBTo0y+ZzrQB4aVoOe0UI+pvG/eEgWKc7dszulrndkjKy5m5KE44G6OpsUE/kbfhI
/qtgccmwHqadMQM8Kye03NLRCbSxwmUPCSnXqIYWg983acvxfZ5WiD6RM2+OaGJaPB9yLj8wpTQ8
IKddK7W6CLesIDu9i0enipQuHHcjFWBz3SBWXiMSFvez+QP3J1PBGe+87DyaM7AOJgkx4o8MQIbh
ukgJT1dTJfm/xnHbZdqYtWZF1gTCp7dJ9h5Or9cdRa024BFRmIwG9lv9rZ3tgCECcp2GIcn7U3ai
4FEoPboGYcPy+9+rOfx8lCZwFxfaB+5Xu3djmQ+UHiUeFCuH3nWTC8o9bE+s1KIfFJfbV0xw42qm
2A8SdQhKGyuS6yqI7WXa5LaIPUHAQhuvKsG3w6GNFYJ7Q24vDZXb3iPPV649hg7d0dXZdQwYoCN2
VfWN9O2npCm/ckVX4+hWmWX0zLJd9yJrb5vGf3av7k9T3MPdJNT1YuTxRwi+OwHxTC8J3MMmySTL
4P7SA6vxo7RcRa8XccjaVSzUe6Sd54P6YNitGzTpBfAu/ttRuInIVIy8/HnAv7sAAnLfWfzWdAF3
c8/aPyW2/X1Ww4MFQk19q3GqbHcZSjJWJplZY9LCsCDepuJRalN6CJb6QxoOqSIgWy7uweA4ADxj
a1ZWwZDo9gcVSNkx++IWlWnFYkdVi/X2YJuI3BEXEOPtfzh0ZScVOa1gAm8emvo8h95Fdc3azUIu
Y1HmDdwbqYXMrgutCJuB3+K/xnVuLIO3ITBTsL2DyLzw6/hlGAiNEb5XTr8ansEMnl8cPQ1PRTMZ
xR7s68J+DxPq5NL9ufqHYrWM/++0nbJABojNfPs2WZ3Xt1/AO1jYvtVRclX2uEqkq8ZAfQBkfLXY
z00Uu9OUBUhdWTAM8M8TdXajXUHkZGTl/wOyJ9RegOodFP9KUs30+0JucBl3r6Tbc3SbEI7GeUt2
FP5BMOKV9SMHxob3uu2CSZieJFEeVBF4NU0bFNmzKtEbWlQrotpkk8eREFo21AHbxDtbDyWzF9yp
MBqT780Whxv96JrQKsZrrNN42y1puu0O+pGl7sHKI/BPwEbanuh9GuC3Gf4IsplkWa/ArBtUaQDX
7ydrMGE8+R/OWD5F5UAJi/3wHXT/uBBPnf4L+1Y9g2e1TH/+WkNsThsg3z41Sa/ZRpBZHwLRpZAL
KssEZJL0a+JtHcCn2A3c26aJPUIrF5puabcZPvAz7Axoi/HUF+ZwcMNEalal5ooToGMCyuR9mcJ0
MtjSWKDJ2yURDG0RCRchwIdcTVVQpgUrTdoodPz9ch3FpT/VkL8SJdB06/ghVvHFZyE4Tuvs3H5N
v1pkhLq4zCajXYqH11UrgSvF+bsLxc6p2STGsH2D7hljqLNO8NypgC10lBbBqOqC+kcFreI0XRv2
uxWcFr5Rjb6coMGOFpJm4K89PRi7BXxar6ILUy9GKYgjzyvpbG0e0LRofO9g66RErcG+Zcn6kqKg
Jl3McTAd6k7hDjmdJlWdBIA1PxDXGLevoyT+EXJXDPNmmgXpmUGJ9rbIJfoqqq5QekkuvGAnQcU4
CTSExfmXW/Lw4E2ZmNbCsYCh0FxPuRIvRnLTw9RWGaiukwT7rSy2BOww3L3hmFOgWZzOMFv8GYPe
rgq+cLZgh5CPHTz3HZBsaugWFWS/huutxABIdmZrGsDNk31a0VJlx9PsOm5SVuR32zm6GeHs6np3
ud9hHA29klh8VqnuQ8KmbqLRmlGH1GNfSSTdZpfWgeldBJLcDS08pB7xEweJVE3N+FKtml6vCxj+
GsTNdRIDBcxrOGpEt2B5ir4N8GUdA2f665Sm29v91W5iVMltZ4XCOZr/SbFm1bbUjYITvWg0R9OA
z/gVEFUdn3oCixSxMT3ftKv32gF61qowqyRAxQ/92UXLa1I4tOy+lgLIp6tFKhh0emnScSBT0Czl
dKW7JwNn6X7fF8HH/RYvtLyDhS+mgUZdXcihUCieKWSYM1T9IbQLKpXWdFhh0RqqPi2JwGeJEQlN
1iBqmgzoddQmvbLAz73L1Hvrs4aQLaq6emfkHQevYPPHDlc6a/jhQq8P27Zo2EcH/tUB+HK81GZj
shuy6maHG9vbYYwrTsZbQsS7mZ1E2T3K6rmRH7eQe5fjL8KzrkCKXdttFg8ze8x0CJ+9UUbvzd2X
67M+MEY+CDx6E2Wsl8+xSDmju5o3LAPh1DuVoQu/52R9tlZU1avb4VwpUO2JHgKlq7vJ23hM0Fib
UD8Q6FKyOKaQELW4lm5StgMVHQE9SN6MehfsQMIddctQ9xa+L3yMk8CkI1DLKdl7QJ68jYXeNC1s
4ZJMPjvwBw3nJYmY6Ux80HPCdytltrHULjMb/Qp/fNjJNVbFdNxEjuyb+jj4rv9YIqZa5/8XLIzf
Zj4x47Btpju9l2+g7F36Pq0Enh1sOnnK2PN/N+tdqvfJuUWlCROPHOx7r5y7YvISbn9fIVMhH+mE
1K9Ly6eLMGqqOVfeP8Yn2aqrVVWDxAm5/EiST28Hfl6c18m+L8xigWBA6O8mI+V49uyE9K8dyrQO
i8yS2bj4kk4PXNAMXHwWS2lRhyKOybne9pl3TRbcDfAYiIlWHCihU2nZKjwU5qp1XRpgFCsuf8CA
lvXegFfg7TD18+ZdWT7Z3e2AGYZX8xDZbSLW0mnBJowmkAcAPzASAKmZTzrNKVJSoztdVt5yk1Oz
KXrqbcdv3G9TbY48AuFQPAnzWT1pufiUix1DRPK5R2gdNAsAPGjBNTsRVqlqTY17sNjnEaVSWd6J
eAtcCTx+rNJDcy8OpDNA5wthg9aG1AcDLOkiw6FtrOlWCa0/54Ste1ATHFPCchXiQ7HRDBCDw0BY
qU0Gf6CF9P7/ppO9wFVrM8QzjBgDLPsPClYs+ITKehOr3MRkaMjEsLdfcocM4cz2QaUYlEKW1UP2
jvDF4KGht6On4AKoeyFc0e14ELqwp5fFjpNUWD+DynbmhU6odG+FMSL4UJ3MYNSHQVIo9YR2xt9a
wrmkxco6u1WkEDX5ARWB6+VoICNCxBhR1s9cnQZV2CiIZSzeqTwbTHvLMZhJ0EIETAxSNCyF9fOY
Q0kSIGn/Abnn6XGI9HlTctY0c+r/3NwqxahBsfkIQavfWtIjqpYxuvrRUEZ1dMZO77CUdixXfHMo
wacv9t7zUuKTyGwSJRtRimHWSuKg5ePrXf+zpN0t0LwwnrS3IU4cBsTDjWJhK9xAbvq6bR0G8306
MmhN6bDsfWevzLMl73J9HymEEVgWTr47uhjpHJ2lIITpRVOxmxrO5lLAza2CHhBm8dAba9F6e31v
sGxPXPByJvpyMTi4jf+o7s0HASZ70WWh9A2M68VHycLCsywKzAYlwVz7lk9PSw2x+cKmRtFI7vGh
0U9mCcnSGVYD9tZjCUJvDsC0vUnMS0RCxTbbVRWyXjfnOjmghCYhm4cWp4IoHOQN2CxD5+ceSxKA
4YY4cHNwARVxhAmQ/leqtoyce9k9ODP/md8zBnPeQwi6Ouxm5YuptnvHZQbIt+xcSbU0oPSgZndP
Y2LOOl1EM1TOvx0tBVjdvUgIWBt3aMuJVOSEJlj5YH4W3uI3kX5CprorNA4PsQQtC2kvpiJvOnTZ
lygz9jFxtCoCwsAvFogOkVQMbftw+hbCoQXnz1ScqshRguMQ3sdflLBk+b+4eSTxA7VPnSCd5mQH
RXgDuo/54piZMJSDHJeLvoL6gkuuInxN0G6/g0ilHJWE8Ar4VYdfg5ue0vSTZbPNjKW/qSP1mE7P
oyGvUttnByegAJ2/PwCVaDc0Vwm3h24YzEF/uvVLYCRvRGbM6+xFoFK5PYSQ3yVsuqmuF4bOwwWh
9oHxP3ciM1kut4dTIFmtpho7P5jk8S2w6Qs8c5xjawgOrAwrz+okGf6LasobG4DaBYkGBu/WE4LL
TbdLGMRxjRL4JxcMWY6PFFbItN8rqTAcTLdNcgn2omk+G1HEod69YbD85bSHdiJP90jVV13QPKXG
N13BE7muHnVxuPqrhVv1h4TgmAMYHzhaAlPsDNn6ygSFRGdyo8RV+DA1xbWtcTQCiN9/+0SOH95K
LcFysOp5nZPahLXmOBgi6urjPxMm77m8H537RLDHiI6R98xFczHCQQTXKWoyZIrw4i4XhwGZSqFW
bkUuQhUb6qifJmiaWgmJuAKxJCogaBp208LsISxw9SPe4JSns8bKUqXE6HIQLeLfE0hcC2PbSvWB
9afLYm6VEMYtKGUap6OZ1ZPvzmnXdEojTo5qZr47SVbtVpkEgYO/WT7OTDy1268BeVQBuphcaNBY
gVVGRLjgbEJClwWKaXR5iGyldrYceBrbbunSXiLZsOREPOAB5LQ9ifL3SK2jMyDE+baZ+Np6uXd3
c1r7rVC9cfHdzejXA5ylfH8NYKFn+b03UNtJwNbLLYZDaQE/J5+YkkmhE27YY53nCyDPC5VeVXIG
7Xb+Zl8R1WlZ10anojZVsORAreCubQzIkeI5FOKJvALxPXT4+qEPZafprICyO8o6CAJvayamo5Je
XVkyf1CiMHJ3lu8AKd/sTCvgXCll6aEL/CzKl53W+1EoaVBravNH8yc2Mwb2lP6qkRg8IIeLW69f
gJ7kQ9kGb0Xe40VYNEcF0wVLfIbsMLTz6tEOlaHN53cgVBj5yUB24qcFiaBHD8g1LS0zjp4XEMlP
xMxyxWPwEBMIxjzbkWcTNTUM8iceBlFzpst+PtX2xb3fso/PG0Xgsm95YjH47ZoB9HXOw1SFkirV
QDGXGya19UCAodKlGo9m2B7sKRlcNpnBjIiS56BaVAM2aeNZnw4qDn/5SewMhlW7zd3fEV/AsY4V
D3VYfNSgarZZ7wnGxYA4eam3z1usSIXYUZo1g/AcN7ybv3SjLf2kW6aoRPuG/8P/hnGq8sWXFSiz
y1ZhtMjNkr1r5PqFB77IGYbMipA1rGIpxKMXrOotpXsEU/Jy1CAYKuWlXUwMdC40ww7czWqJ2eE3
zHqiuwYxXMTUqganyxhCac6KqDG+vYRGadvw0f7pfjNpm8uNpwuZhYAVuICy+N+kC4SuzFFdqWpY
hqHMpHJF5DQ4y3wo+MTatrl7TVNqcaxYwq87W6IhhucdBUP2cWac5BKfkPanT2YSf98PWHa7pLLU
tHSLCAoGP0v8Y0QC9UxSeoxVvmz8mL/qw0opq5GTBx+h5Dt5GbctB414Y/hf0Mb0y5ZP0hZtT1Yy
kkqfy/uTKs0IjkKQrGSOmKg3m4pcksqMfil+C8eXF/nh7UH6A7mdvqngXHytMrxVOcKIznIhZsVu
ap7LxQVO+QemMTVw+QSUdWwXIqargpyeUOT/J7CeBD5TPfeOn8K4bOxCMrNUnfFqoWnqr6WrwVAw
+jpa6cUJQhJbypDMimhln56PSJIl+9nopHjdyZm/F43FHZm5aLzAJzddpO4Rr72c4rxlMQe8kjQG
TMrR3JVbEtv4gDf2eAO2q7BRfARKmzYYaH7wEUN+vfdkMG2zDKWN+4L6zaVL85lvILSJC0MuGJN1
f/XX+aTRTb05DLu5wNw7BbWiTiFs1SYXN6zPehUf0k/3jOfdPXGN/pwwdkN3KlxsiCwJsFX2M9ha
USgc+673EIBeTLwEaIn62J68/eFxwr3S+YJoWSQ6B6wsZ73JSI+oQHPqcqStBbaI7vU2cid4dt/5
5Eh4eMESHUKy9XgV/0SCaIWiHIcVkEOFOog60Bq7SJKpcC1OUDI+as01OiSxXEY0hTsNJ2SS4vt6
KvTu5PXEy0NLWSvmddItBF5NgElJh4oRkiN0JZBAsShrkE/gFsOwMPmZFu69GEhbveYQpm3CKkx7
muscqwTiiRFDN5r0mCptK5wIozlo0VMGISAPFO7Wp7dLXYNi1ZphCFHI5u5xdd3hzSu11JYBFk2o
5HAH9onh+P4yJbQnWf+9xx2XrSRpGyRQTLo6MJOwUcmS9W2TYAKqOjvSxwFT+CzoO2fhir9ZE+/9
W1WdG/T7l6qT55uG8rcsgJ6oT1+Sh2ENpOc580yhLIpOiofVcAAHCUUTyDssDOxqUthrOkWd8hFc
d7NbbshrFP1gTG3JEIZvVcIsCad+HJSlGDQU5+YJO8MQIxQKGQ8HhvmJ3BN3m87aAbsoJ8MNZFuJ
ry2mRJjFlvEfR7AAJ1E38EARoCD7UvOSHoSCZS7zTdLDIy+r70wi4AKnP8vqBHRoJdp1P0uyzWrA
FqoONd1DmcPEcUMFH8HHo+kr8N++tNPjCBhURjhrgLP55zL2sd2adiK7Z5fEMf1WVmhNwbGuqghE
KijadqDSLWLDhaxkEcGpoUvKHqUHsJscq6jLwRknZYh58H7ofkFO13LzWRNygUuaYeGx1ipkZDim
3ascFQnGtGBHSOBnR0CgHzm1NPt/6yWA4T7VcDptwOFsFxCXQi5PcnbQVfXAJpdlWUIQrfZoz2S5
TVv1MwFfag6UVPcERguVe2TjOYfcHLhm4iGbb8GRmB/sN5m9kk2gfcYT+Et8hgQrOVfVeDpLYmeo
6V0BmoNB8NqLVJvV6ofMPv+bcJ3OGs5ip4bwmNKQ0XTNj4v66bNL596q51i5PCYfo0CiQMZhHbXH
DdkIOMkPio4uCF9WoLB2JU6QxmrLNiee/WWNivxeQULu9kZ6gQ3GsPtG+pI0NeilMx8fjp+XLmvE
oeimLnoxQAmu0OLTo6ZVQykZyDKwZnGDMZpTqt0DnNDmGFhUqg04lQ30LJ23B2E6e4VUaC9IVlEm
Fc8swWo9w9bPZrJ0+khTsM+ykn9jRaR3KkgKSuu16TBB2K0XiafkMuhtuXTDXZNPAt8lRtOom72w
Kxonom0lIt+Fp2DQDqexbRyRdrWcm32LvonH3lCra0dYlboYw7IkZYRiidCP9GNBlYhIPALK+cmu
5WIVzEykSsx5wl0tjkqqTf+6waSdcA0PdoTyq0PmCopFAqzeghJqGE5kaEdi3cMW8o542FWzMBGJ
V3PF3IgTXJ48LwVhp7S+rdWb1Vw9IT21iGdkHr9qjuZf9Ayzbo7VgBevrPgJ4hqiRv8Ux0O859Rd
ZhQj+jpW0kXj4LyOf/p53rdBmXApHLwkZ5L5lBsWT1MDQ1aY2edtRKCEllcuQjEoWomkw9FF95g2
Kea/vvHciCeJe3fRGfdzpBkAKYM0TMmrKbyiQyxip2giCPAOwKeM6hlPpOlRgD6rHy+6qOKNYVnn
lEvYWDqIZwXLIYiJti3Evjs7QKJo3S8DXkiJBQNVzDzGORmp21JfFqLPIYqxSCrlByg3KC9WBptc
OYmmC3x6jviNPJM/phQRy/wLXhLHl5t0my3UeHw/o/eLjOUn1m/1e/n2znOj/1s0fE8jivvwdkdF
RFYUnKcsU9gCs/juDlLeotgugYsacavIGgvFAQFqb0wXu0ZKUfj34CuFr8gCa3y4XVhNZHEXlReL
0h4FyQA1hZfwZbY4r84VUNhMwTB8IkZzhegPgOnZaEd0Gfh71g/DLJQBoP/utwlCC7FwER0A+TUP
AD2+YPRafZxtQKBrH0wkHSobG3FTC4SGhwZTP5QVmGmGJt7qdR/d5vftauP5j5K/gMH1hGYk5Oas
F8Xuz4zKbt10kdhLb6zrSJN5/wh7G0MDU0v57Zj12i3ULwiFeoPTuXAsxS3SKEl1C9ZENAa/A6y8
g5AinnD9f/CcS2v6Ar7ce7LWIooc9XI1+EdofEVHI2untALyPDdtlq0O8x+u0Z2A50b4CEWRMbkV
aUDMXuIHyoyohf+C8HGZpt3Bmu5rfMHmjSemd9Bz2ruV4b5AmigUNoFgvu+Olo0c42nbcVbtbhMw
qERmaRtG6ffuIBUPtk88RmxlXEDPJSocjYCoJkqhAGae93CrZhaRqkvdWgBMxjUdi8KykJiEiQ7X
kjmA63OGYa5GBa4TC9SF7dqHtzmUGJE16dYiDcbHtyBPeY68OMe0dWUfpY7XBcxSEiUtS8VsUcfj
YImZP0uNqiOQiH4QHfaobb0dqT34ZdURuvOjBTpztdAMYi18zLGxiwMJ+gah7yaLkkAJ3DnSydWX
8PPidcnM1345sHTLg5fFadgtiQQm29tc36inczNK/KrxQNs6dyxb9kbgdEv49BLIiczD41vso/W3
SK2t9/CFIJV6KzwT5dQrQmQe7rRgTL17e/QZ27gLgYzNMdhNM2WOfRGbX/yMUcDKNGUYbwh/hpnU
4h+Ie+PviEWbmS7vAT2W/OhIZe4xkL4lNWAjRNEUnNpb17AV29F876xT06aWcbfKtWLOK5iTrJCi
tDQWEp4WeCXyY7QrYI98NXRDbf5vOXi6E0KaGsoCMFP4yGyFm6gSRw1Rgc2rF8Qb3nUUYM0JuFux
S4f6/dlA3vDTkZYrb0JjYmd4q7qzz5NXPNyLRoAfofVUUL+S0Kiun/YjzLeB1P9mvMMSOIxPDlTH
7Yry2zerZQenVWd7adYPJhIufXrRGY/Y2Kw5Kkq3SO5kNws7yZivu5VHtUh0dv9NYNWI7Q2K3ABF
lL1T7KIXRmQrVyWue56bfmAP6YBWyJy+r46+nsckc3Kw3C4YjN9asUKNbzGbmN6p0jc3tpCqXWao
yo3Op7BJ+KElccS3/nnYDY54kaaQBuz18IoM22relLXVEZqDC2X9qle4Bri9B8qKGNd6gAaUqBiN
RFceJoVCpPhcfuu0gO2tm0VJJAUFS1o+ILMAbAX+8mqwfInlBIpYlzT3rVvD43wbqj5jwcrPCkJw
shG5w7KOcNH5dqI/gWSL5KvuM5Ewz2h3RoIjGf56EreUm1D8F9AiEgLA9ZS1M799rGsfcOlf2p7n
I8wewF5vUmWyvjUFo36yylm3XKCVVZD9GwBOCNN+9gaa0larYUjZWuMTS693VbKJdfbM1lSngA21
/osEtQLO3Wg5/Veabc2xH1Bk/MXNf/6Przh4HvtQRHZRFHJXUvt+QMYsmD48FVq6UHJshzalkI6q
ADlOkcdgMQghMaHrStpTl2ekVWiB0z6eaMZUNz/AXhglA/HGSMc25GZCkyf9ymC4obgMO1Pmuqm+
8Mh1CkY7BGNgglYGijxYMu4oKNoW+arSu5i0r7aiFfRTwb2uT/DLELevmc95mOxlpFNrFQa5vD2k
rM1foK0qWFTdTwYjxjf5NmkgRW8tLBRmMXjZqFKHl7G9JHhoU5T00wVcvuJaJPKvJJ04um4tSoMk
40Fmvnnh/oAH/MlBfy3sXc4GzmDhU55ZrouB7h23Zhau7RavWBXM93cciBoq9HoUkZJR+9/U1sng
EHHy4J/tBmDlDWNINcYoDQXW1zNxC29MQBU7Lomil52dWU/bc6z6Wagj0hxfu15b8/pFpYXkZSw4
yd6E2zPR+5V3RHRoCXyoMtGC8/jfLcwOWs5mNfCYMLhL3qW11xtOMsexihKWdpIhgb2XFB1hn5Xv
V0u7zmfe7wduWIa+NlJEcRs/DWd/HUZ3DT4uP2uCFv+9D2VZTTwx23Ugd9vXpTkVRwWRoRDteXde
hcnJd1bn91yg8kF5j8cR8hVOB4Ot6jV8Rzk+zW5kIXHsw9r9m3PkJQg4IA2aTizKI6WYzQrDPTbu
i1dJKjorrgGb24bXa8AWBi9OdDhlcvM9fe1bPtVvAKO2ve8q9nVrcZSE7NAk61Gb0DVIvClf6ogZ
MZvvksn33Yt6KC/a1w8VpCbzE7InKOqXf13Y/AU8bMwsIir0ytgg/GHp6lofIOuKUtfgi6qHoRiL
4bpgQLqZSsMx8t6vUH6aGOYxt+u4rrz9o91ea3Mzlj/AueyaMd1g7hFIbLr5fAMvHd2x2pXswO4D
P2zrC6MVOrJwKZVvgkJOzqU+KrnBVOOh2B9x7A9tlsZ2C/g6zCIdXMjHXTGwi2nZcHYMtNTprUKd
OBdtNuBIY91mrSOpsrNhJNcmKswg/zcC1zaIqJuxQzY8q0IvFEx1xDbuaCVyRCy8zEuyJPj5cuQE
r9nR2V89+ohjPQPRPedBASQY/UefiFFn2lrb3NukuIIBmzpancNVTGZohE5L1sJe4BuQXc8gmhDX
sE5xpc+si3CTHi7vFdJoxsOfMRcpppuEwHNHQXyQYuLAPj0I/iEDhhK2ETMvE8YC9+ic5ASQQ1rm
uJTjyXNC5+hgQqUmyudKuvOXleeHQSwn0wFSV3UiVeCLcri+4MuMYktjAVaZ5YnfbRjZSGZsydE6
itiLziw/aAWT7uuoE4v9xOE2DDXIML9f6PLO/51W7ZtWhngko3aHMMfieFpj9LPUrL4ciYKqneWo
BC4XgsjAgr9ZAHEPg714G8m1CwW4CYeu5MwnJ0v9IVZv3au3l240TJssxrQfwSyaE41diMTb4vuL
z/b854XG6K4TfOKP/jI9+XSwEflpit50WIYZsvmfdE6OdYArHF0HU+wluGU0ra201WKyTqkyiBec
jTudBjaooB4P6NIPpoR7cvD6PiZH4z70vDYuya3xP5jj6mQmIdvLb7mPMYcRN4HxoC8jS6ffk4bP
oD7VMpHdiTF75U91TJ/zogZlr/akrQNvp+u+D0nSK6slVAUwp22Rt7L7+07J5gO/nwNdoYkkpBxN
UZXOj67UewNhuIz9ZCVDLa8/DuqYJJiWWgS2iQO9pt61ARej/rchr8lYlrVUenU7IOVJuIpWD2+a
hXMVnDQIWv5UiG40zoQGJM1M7B2fQ3I3o4ylcLl3wL8bYf9HDQsJwJd4NY/yPCxO2UCD/54i9isz
n9YPyyIzbPUtkl2gUCTpl3mNhqla/AchdkcPs1zM3655bm0padV39OuxRPFRXDHTlZz01zDH76kL
5ELbpHxDPoE4nljMtfwvNm0yahlcbvQwVa7UU9FBuQufl/EZ6psTVb+lCSS9cVTMuoR+NNNAWX0L
+eSMMNCEEgoCds3PCK0Yx3g796PvoGrmQIGwVFuSMHb0rxtCQGSv/VdGKOQP2S4N3ZChJ/KoJy4m
txPLjqsET2jsf6EUwis5kQk4p0NGY1avvuEMj18Bf7viZL6dWIwe7w3eqeWy/fP4Gbiyt6ZYWUdq
XBaROARFRBblFrsbXCUPtka5yennjHkjpPuJNLi2MOTyCCEZgNy/Z6R0IDjzLXRTWbbogAOCQIoK
4XHkjT9Ed7pel68kAhj0Do7tcEO1xCKiN9HXU2J0pPBxeAqXlmb68K1C3lbg8YcTIgbccBYPaHXV
d24kWjFSmb97vWu2jlvZA0AozIlr/xh/cLJyO+tcp3I9aaKXBTIpU5cL3YpF24n+5/o3hvK471sv
RWuNtDsbyrM0+rCV1VkzfJeODwE4Io6nxVcMGSrKkVS8wXD8JKjHWNtzsfktYB9+yMNgC80y5n5P
9N9U+lUxW/eNBUFAhuoOuAOVpXqwzG2a1/kO4y86tTru2Q6kKTM9XtHBXKeK1vVMiK7vF0MTPehN
NRtbWG82rgVedmmBfSApaQykEqvy1g7A1I2ruwBB5edEP4H9rvXgEv4xBRc19OI7aufevVoAbZpR
3ijzAaUYsqGCwmf0USySteQeqFaEA2jKxIKsTnY1+P/Nmqon0VmPT+wh+wGKzm2RSsQZfjcve1wA
FVsXA6mCcB7sdXg6YQ04romDuDzYoiVpTlaGBSexA4kBZAZHx+DoLycKCX8zCqOWmYJc5JdGFrf1
g4DtbGqxqKBudowh2+qrGMwQq5TnYH9Dcc7zCFYH8njNq1btPw9kcRbo/oE0FdAdcdVwX4GGA94H
RPbPWZ9ZlrYENW/zrvLuoJo/nZqebeTs+drY6vIPvzBQeA2bqOXfey23azpdMwm7yeJA9xgGcrdr
cfeN3r0qC2RljZxHL7S0CffPK8uhvf/QtqjwqVVw+YLGI65N9P+MdBbXkWaypf3gOOrcj8trCJNE
w+7YTa8KmEQEEfgO/kF9EpdnPF2aedwveMsodIxdKBt3uRfumLutxuhj4wkvMWS0lC2j4HnrjY2H
4JB3rroBYrzSH7BzTf5gq7RC+Ib6dpBt8+oVf/e9bS0raTsczwbfYsIGLGA5ZASd6ahBg0HHyAo/
gpin+mbw7EOjHnl3yqzV2ZWKKQih82Tge55DWxcB/kVRU8EkOg7GjDKhx1PFAg5VO+JkBiZAq5z1
joyzLq6xKJOz4pOAZSg1fkoMI/n/H6HTpRwZV9kL1eZPBU33udS0prM3k/Wynka5nMxItPiftF+3
O3V4eJZDZr7+9I/nzdLBGnJ/MSSxVwK0p3/uiplzX5y0pEXO8et3+9E43BLit69xPt9M1n1akRB0
5KQMzODuwbWMUYkGe6Mkfp74O2lV2a24eifiU5SnwwDzqvXZSPGM5wVqAxT/BRa04J2T7OOEtBSL
FeZKqTUiVVfyTyWNrVE03x+fRl33fYBmy+R2OLw8ohURWsOp3zwCG6DzVw7I9Ri4E7lpdoOuBzvs
4A0og/aHVcbKIZr2qqZ0cHDWwRGFMPsSh1+Pg5kVB81G0uFMb0o7I5V/pQYqcktOiKc4nIr0C7gs
ovRVIl3iPaVGPYH5eZ1XEIpt+ES6UvfiF2P1MjWGwLyorPnYshTjrSyjHmgT0f1pQA95t3T4IENF
cAMkVfdM+0NP8efLTZIkDgiUO1IVwUV4aRhVAoxY4DJ+/nWzrRSWl2uyBEJwfJ7nfg0P5jOprwnx
gbmvCgnTArzpbp93iyjXeucHo0PyeCUVoyorWBRL7fIRUVm4gk7ppyQz0zo/UIy6xza74nfYpYKa
s74KycUGHYJPc1pvi0O800LkWaNcjDX42aWwY6gYP8/sCvlRYZIOeuX1zj2oSJZ7nDI1iitgqLOX
QyxID3B/0ax1ct7enGWRW/L1fyPyz0+QT61w7dvoI3znfEwy875Gh7fbzlvc5L8DxSJ3/KpjMpAw
XuMGlVHDGQ/Fhu/depiKRWdSvqRX+F1oQ+buL1N36f2Aw8oBdf4WuU7Z+Ph0oiS7Zwy5ZSm3jSJG
Pg0oSp+A8J9C+f0xcIto8pluhqlC0MwbgELmIqHuy/uXym29mM7dGsjL6Hozb58vPtuoD1qgcddi
/x64DCICvxCFKXhsheVdxz/lb2yGMUFRCzNN3S7e5yLU0th0fDb9cP+0kz1EuXqvxWxBBfwyIo8A
Oh6Y6KE94NPuP8D9oc97SSx/1uBtnuuSTUk6MT4yPwYyChs3jWTvz+P0rk8IPRXowtCwgAVogQSu
GUeH0hHRH5zfbrbckG4oyXaWD4BTGSSBp2GF3Pxt3aJfMiRmKfQ/qlbXqrWksZjaJUc8yyNb1XfX
xQ04WnE/b/LnS+jRK+94KXd47+43trLUGgxgRuutFXABbH5jA0Q5/h1FVm+9dHzRgonul+TVgHvQ
GH3Iw6Fb/EgrYzBh7sXS+KcwiWPJZiqVagM0N1RBgBgXn/bs/beR+inu0h6Rtd21gTlf/iP6ntGj
iZCkrJBc6xYOnZ2kcoBaiOGvvgMIs0IHNleoDag2T4jQVKsfiR96v38k+992onPWyH7dS+mc5do9
fAkoVKtEuhqD97agnYyBsYImEft/fBD9idbamzAreNxgQDNHYy91FZLBUu1R3txk46uVQ1YtQ6Xv
yfEHz3mbNzvZ6HZwhwhb3cJXpMuppWkmJ8hrvTRqSoBnWX/NpVw/jCRHL7BN0TLIlabdmQNugOhS
AtEBWh9klZJ+kJEBT2NVFlrKwuHQI64tXDi5qY+0vpl4cBaJvyM1J6FWdAdtaGuKgwxr6vHExLuj
tGJEksQ+Xv3S+/mlzJWH3aj9AMM9v6ZKoS/lwAqx3gO9RXTHkQjWQpYpoGvA3UtRKugZAZTV756c
JFNmCRpcdeX5HTWVxHdk1bCsvtW7RffcfVNL09CnLy1QMjFSLr/UqGVU1+8NODqUIF5BqNjvEvoc
rMRKbwTbOZVq+IihgshycJGwgedG4lfPhD3EO1BZza9n4kAKmv67PgE2ZOolG8Jdib3lvQMhsdOt
YUweG+jljDOWjxlXEkaB+bbLb6IG2YcQNyZDQ2XLMy8dLg7xFbefGyaHjCeGIgSnOQS6s2rH5ny1
nYZwZExE82ZzTXkQkl9mLvV02gZ6cvyxPMlcalhj1SzAmWDIHmTVnN90ktJxiPJvcAi1y4tL2VIN
NyG4RuAkjhe2LD3KOvjS43c/kf/P9dtVne5dyHaNEmuaXpH2He5FATbi+K3c0JYjuND8KfLlFXVk
mUAitcuRz8DEbUXuSp5NOu/Q7tkFN4F+vbB0oDUDDMEicguYLvbFb55qidPujE23QIr+1k8UsSIB
QKTliIKn93bg2zppHPDIN9u88RlgYqkf0NGKyedSeku+GZ7pO316pxngrkNQr3UKOluZbmvsiVc4
a0YNg7PiQTuf8z4sjsMUxxoEY2SF7tpIqqnLzrAZAw8p3jnf9A7BUOv/iuT6hvnKaK8DsE4gzEd5
47uA4McmK2gzSOhsKLXKIscpVRNiykMTR7rJ+ja3+BO40gmbq1BIlOLgJX/Ih0OdSkRK0CthEFRx
JJCW04x+CGQEMPHotElba6vBeA4jdvBhBYxSUDCJD5i3/sDTmVwWzelUkgxL6kKevrB9uge+WTch
7SImElNeluJQE8e+4yMmc96SwDdExkLkXWfvwdO54RD5ogJtRxy5ZxlBZlyCzzotQWgHGPCfre/7
12dRdc1fzcLE2XG93C+APTX5dVxZVc1qV6qQRXQ17CrAbLIbuUs4rk+fqpf1KsOt6CFlTUnQklaH
mbPy9DqHiBdbjt0ff4poI7NISme4B2c+98R2ZXJaA6ntRF4DCHaYDhu3lCZbfzRCxrHz28aOMZ5d
2hq8Cn2NR8tF6g2HIvdistcOZGWf3LCoxZdkTeiERfi9K0bOVO5f1geoYDiIf6G6/YVUHcMb99Lw
CKKWzrPCcCiiZD8xBvIF0TnIJjtUFNzfJOpaEM8Z0DEicZZV1JLET5RfSE+n8yy+jaHUbf1x7/mH
rm2n3QWHDEQvgYWMFJXPk2IaF5fk5CLM2hBc5NbGFXjkZp57ZZ0qU+3BZzmr0kusK4KzgLofMg6s
CBDQnJKwcvK1FQaETUVtI9s1aLmz1mfe4ZLGlu9m0PdB3GJJXHuG9I/aG/AerTu/+sI6juyRwGqf
SDT2+Xpc1HaVa9ujnQqEydWDyWkGfVnIdfPtWKOcZcYQhGzz0LlGehJtIKOJuRRSpvnEEyXZBC6m
xIfXZ/mYtXVl8axVRd6y7T2Boih7kvXxJKrB/gn/ZZsBr1KYiK4O2arJNZ2yDx9qybC1WG7j/qxd
HdKwFBoIRAdhPQlRxx5dGCKPZmPBKa81JseD1eAx4OACfPqwXGzA2hGZICDn/S7ahj4KGN+btt/u
Hx5uM04vZa7bJbm4N1AGKiegZM5UwUMm2dwpB5I0J7t05AF/UYySmz96aZcFlnxgwQ2qexng8MQg
wI9IjhNTTb40j/UDBswlYMAbWMDqqCKyPccvGS/zQ5svGfcWE2mix3KZHLAtnccM11lm0H2GwcQn
7y406Spa+mYkhX0HsJbjx5x/ylZjMMktIRL62+Sjw10Trxuv223gEaRffNYdJMr78Zz23VhK5FrD
erezNrvQyjeLjJPllbF/m8ceAG0AeCSMNgocd6Ge8Y/wp4R8mbSVPSYEayWAmJQ4SxMNHxiZvnJN
Z/XgRKT2cr1dZG5cNFKHwQL/7R27lz8qo60neSxAa0h04/RoucWZlmyEON446ApoLkHle46gUuZL
lR3Bvp869ulyKfq+giw9L04N7T6n1lrPH1ZvkFcygZi+v0bN7zCMoWDYrLqaCnVbF2n0qHP/pUFT
aFkGiedZs7lHp9jcAoyemI0CH3wu+5XC1jvfG9mADOe3InGRZF5hPL1+vcRRC+yXeMiqsHY6dtQl
MNxo29fAvl7UVTgzWinVeiCxjpzUT4sWsdEnjjHeGjADnnm0qCdan89xgl9jbKTDzFipV0HdAiqh
nZl23qSuoCKVaODZXV+siUS3kL+GEuX0mOssAoV9TEaZRzlxTeLNurVXweOmt2fQ51KRxSEZA+VU
FMrwWDJFKZ/mNWmFkeprljmDjfrNS4uOjspvs/v8aYI08lPgULB4vrhgd2IoYevcU2PpIjWAXTls
jyWNROimyU46MKmUR4CQj8KICxSztoHrSTt9CNOWojg+mNAtXckg20/+k7g4JfsuO8LIW0v6norI
kCOnum3f1Euerf4r8hRkMuuN23DC5UqJ6gOlj8OyYdxGwQT2DrQpPe0/njhY7JFZ/9bbB8xLR86x
LUE0LViJ4yKO5/jFh4Zr9GWDAnUwCXodhpM49PPt2nWtp8dKdDFeXUi7EI8E/h3Yv6hfv1OzvwPD
2bhaqiq593/scMudml94NiowYuX3RcOxawMTLk+2+OjBPbWPAvZKJR+xuFXOfHDPQEfWDTNYckhL
rXk9SLS3FijRHurtHbNHSElBXlRRSbAHDCVCNVVmISJPxJ6JMLtkxf8V9+jNZO7ntJpDjD7rQBAC
Sas3twJI8ZZhr37Qypwd3uSlQlEIN+/mPxA9/cbGLJs/ueXirAXGT/YdFAeky42Wga9wOP6YEf3N
My3m6colR0C2uY7B4eW1PhY596ds4ECYDtD0pgCW4iYPLfNJnfqJDwhSX046oeOyXp2mc/T2Qp0X
AZJ4NmsNApMylTuyFvtnSaG009I4umO+IV81w235mdqoun1pRnlQhpffjObKZBz+YDCk6qukNEGZ
iBRBRDZqpy77NnZbT5rY17dWut3RaHtNA1d/tSyz0ziwV8X8h7Tsv6OxhSl3nVXwBzo8xpW6yPe6
AhhePcoXfCNbuEtjsKEx6bbhOItBChbgkfiRm85207ODIT31kFfCXDb5MTTiY0RC2HWE2Gsqm9h6
yoD2Jy1KHnxMEvgJ5NGQvQr6csGa7yLsA18+DtmFO1V6+LoPV0sI7RA9z8++xCZV65+0QkgHxAa6
LC7617gxkQWGRIXe05JxevAOBXgpvB69BsMl5Jp2zLJaM07oht/D40xiWkbivC9Ea5fbU60wnwU1
hbt91Z2XCp5WNThz61gYPUlIRAJ4bYaQnlkn+mkBnU8xquCR98BB3PgapJ6ThtEI4sXWjNrAWDun
gpLw89+bQB4z54y2C78CbG7b6atwfPXwO3MwiLVVE3ZwhAQnn8RJsd+OkNQLKZKP2j63wMBvCjP2
Ylq/ftkMmRLDXB7lyF1zUzeoFM/Bqm4AHTZJJS+4uhvPvpzPf5oG16emz7xdhEN6WcUKmHdA5ePZ
I45eNiTFbbfJa91oKis42zA9PIdq0umxizwTPzsWxK31JvbDz5RG77hNrr0Nbi2slXQv8eggzwe5
2iPyT2KCrOh9owGHvI3xsFAdf/FMM8IVxrqrlaj0xTO2qIwcYqW8ifmiNHvCpBMKf6+Pzzi3WKBH
EdC+hDRuTsK7IWnP+POVOIlOf+xl2YJuR125pe43SadDvfjIYsdZf6Z7TCvrignlz45QO+tRjETo
CIrdWFFT29AST3/+V2nSEKVw3DrG3gwyRDYFq5KOj24xa30Ax63CMAP3hSJp8eiRr7oQAjh5f4PD
zEQLhD9uo4Nw202LiDEH6ifmI1nteP1y02A22+sF8Dw0po7Rvgeq3Hnu6TYZ/Sku5OGci+k33Wvw
R/GrMQOtne7raUp58NWJ95oVtEwrJybQCowPj0Mu91FnhNiegoXB1J2VSeAjell00l6q7qEX/Yy9
1b7FT7Eiq1xLV1mShnFmDkOjcsKqwfgfvBH/SXWgG07tSP8IhtoqbjrrUnOpBgSQJiIhCFnz2iao
8/+BN/hkyFOqGwvxxxstED3kBR1aaC1lHGxdLjhB3R4xQGtwIRpGCwHNNlyBraz6HOtnTWB1kmUC
VdU3CEqoe9hwQD2nKcp5aRJiEVh0Iocox0hP3WvAYX/pKP1MGRYe8dpMEG0YF+oVw7r1eYHQdEr9
seZIQhoWj+cNYyzmcVR48cU0W1B9I9mYCydf1k7IHfuZwjfLtfT05SMsWv0GKtFKzDgePHAWEU3x
fGShVQTA84sBnVKkAtvET+w3w3IL3C5bjHTNCU4/Jg3kVUWM/rUyAYPCWyg3LXswCUmWyP1UVccs
mT0Z2xlcv5k8vcoCnIfOJsgNb6Md22bMm4jeqLPzDdDlFFsRsvpqLYMnT/EugiF271Q1RmxCYdbA
AUEzdNeXmilvqCgeikKI5gsA66du1JCuRv/0shiu3bBejvt+emj5rINfNTBZCIRCru9XC68NKok8
dBpOMKX2og4c0jFtDo8kzCbxB+TWjCdsfkj1gWuVkFsnwX2IHxMEgHBIAiZphuekzMMBZfJG4BL0
pjeUGkrZxMQK/yXjHSP2EuVq8Rc+kStwcrdiNQdq5+LEEv5LgJbY+jCH19ZZisOHEKLcHsUhOfna
45mNf/f6N6kLUbjKuXsNyIAt+goQajDHvgMVFv2HgEwq6t0z393j2SEhF+AHFZAU0R9JR1nD5Sdq
/VXbbZDLNE0hH78wQyWa57JicNZQhHR5SUel5Rx1yNN6lQdyjcFPOF46AYFgsqu/kN8TQF5YHkMx
eoLwrlQHClo9kz/rVe68hIA5Tr2JMaYo08UvkyoKL4zpCAje7c9c9jhwgFp0yPLaJY763W6VoAiZ
6uf6dZscbDnnfJTB3CC9QY35pB0GHAEE6oBmQzyExpt4UCqdom7VxorulzBX9IlkQktpoIHwyAkF
gXnlJj/S+wF5lXTIUGCidyFTQPVSXzyJlIkfJZ7NftyNzqrz/NZWhsZAEOn0p+mQaMH0hqdvcQ5L
lNjvaJdILtx3g9b+ZbsmM/2J2vYPf6nb3uYKuK9hWefbdXxcGkEacXajqmoPI2iULL57kuUKx2i7
luC+Y7ffT+xDT1gmI6W4DIc2sRvEtlYQupvZoW3HKGH9vk1u14IMcFUcz8scT2/pD73a8vKfnV6L
WhlCZi9TTvqGTXL8nPrjtyFp/5mmbR+Dl6kk9Clm7MU+n86sTDqi3/PxJXVd7xfKnga0DQ19tZcA
4R5bc0mrYg1vfiFTUBG7nZIude6TV2qWIWzTexH70E1vp2ANbhiTiEzrpWaPIXfoRvY82o3DBGgd
IzxJtxoYceIPIy7yFZZSOfZCVCCxJhRa/MAXtW9YiQZaBErwjSELHoR5PS7mmz2Fqds012roNXG1
40eYhIwLKczs1czxj2ZvPgp5HJleVlWqGYwXMKk8nErpcZD53vSoq37iCwpC10UJYA1JiQOKwyGe
slDdFsz6KyAMcwJtilbL8dGCAY352DQR6mqqbqL+0T/7laiCWeTkbb7KrdAyhAjCcEQVCYcpneCV
tmd6er/pUktPOhm7olzPGRvEtGFw5yyP+i7mHqjdtSxoihLmygmCEepsCuESb8dtQ2rkMsBE67d4
dSxxK0K+NEY85JO9psjo3itmK+ms2Ytf5B4hQYtKeVx7c6Xj/MNtofIgNzWYE+Mpb8Uvl7vcS8Xo
Ays4R8cIUtMaTT8ZI0aLrCDApwvjL8l2wT3LJpD/AWWftrT5nDiXLJARnbz1yzpWhB9BWOF3oYRc
YF6PElIKWJMnNb7P2EJlOtFEKmcdQoSk5n0hzJOqvPpPU94jin3ZHacX8bSC55tHXAwhadSyNR3D
BaVRTLG84HFfpKrkWCEyWdXC8tYQHIrLGGzIWXNYkUdqG0n9rZA5NeqAILydRW4oJR4lzDtr51YD
C+5B+5a32bhY81ARxjRBgkx7Ai7fah7yUTQ9pgOhuU2BrW1OppZYt8ur6Ljj/ynorIRw72VoKqFg
QCpJcbX4oq6/jf0dI0kaud9DraPNL68GWBWwNVxcKM6LJ+07OU3rOCFEF5OgXqg9C+8rOsGZIorv
WmdnJEpHQJalYQLYVFv1uNIUi0ubU9nYyrcxvukd5oPHegG77bwlYF8HQrj8y6oSuxyFHp+eFvtv
XWCZ1TQ8RdAE52mjqsxSFOztBxGinVuL1aQbCd9Z5i9TPxd2eJwfHCziBBak5LEGo+y+ajk9MXue
qE8fXsw4PMEUlNFVVEFTPyflidl0jVWmg7KOXqgFp6APqfME4lWviMwSdJq1PyqXivAnDhaWJUZu
T4YmVg/WdZSjkl2bcX1DUPiIu0QZ+wRCfR+qcvvGQ6xJw9M3RHTH1Qgkf4jplGBj+OOUNrYszh2Q
ecHcYK6rydiV2PXo6GrKyPForBk8iSUB0SNqsP1s+gx+DHY69EfSu9oBEw8zk45qDKjGQYvFbGdi
Pa2WzIXRjk5XISZ1ldwlijZvcm2cPTlJTQtUIBqNDuCiMVSkE9V8ZRBE7mb8dV90Gb+jp254HVPj
3Nj3GRPaNR8EUCZ1a0wEdcJ3qGzMb/0UQf9+PgY1SggFehe5+j2TRgBqNXCzyi1xVSG0sYkVC4kK
FSjM/eiH61Cl57i9k42PCshdowXGPBqZ+Ro1YJv+NgQEa01ZPcnbrhCUTt2HRR9CqIa2VUQiIdwO
BjEDfrxOTYuN6D7Cfu+FZoUZVz2q/xmkbBVsy+rDiZo9ZRvsWOXmaUhtg8YpUBwj7uc6JniE4lj7
RtjBdLHI4SHwuqF/61bBPCVriRBhPdPmg5nCRP/CpNGUfIeH5D/9WsMew+udx+Pn4HOEd6TYRivK
wnBy5y2vpBvPrY8AeaR70ffvldNyOnjwjPk/paHk9m7nFYU3Jl/RGj+IuYhiQLgRsMKyMx2nOKbM
TwUE9gJ9ktfojBL8zDgcXu1F9rjQYJkUkIyP4vB66D2qVP6VcTyEhuUb/Md31NYA7CATbhaNHsRt
Zbx4NkSIYCX5UgsvLK6TAW9+RQmqVRyrPCtNe1mjWntden9JirQycT5LQKpQ7fcIE7kQi+wUDF23
Kk5vIQpsVWbvynH+tLanrZLRTXQbAhskyEocLYV8I0iCU+zEJPdAmdMMoKOYr5o0yJh+lTRCO7pv
+bbhLQQ7PujZoHimSuLRRr/U0EQ2jP1HNyH3J3ts/oZJ0YlRzr0/iq8F74jULlmDA++tauITXGju
1lilEsehJV0+7dJR4XyooKQltcf+HN4gv5r3Am6lUbUQZwhU6UcRfecFsm5Qdo54YtCYO2zJ21/Q
go3n+2WmTXZUDDmssZ2/HjQbKsvXjGJO8LvvACLcT+2mmay59wodmm3VddF8192FrV6SwHq88j92
b5hdo3bHl3+noV9RNsZoVqd6I0HocLKFkcIRL/ekh935OgmqXhj+aY9nszoooP4UCW45K6qhSE+V
3QdGX/RMXRYT3Tc9VX4zGPHf9WxKOS+HYTLi//LwC31YZ98lpI5YmDssZF7u0PR+ml4vvNe5AhV7
dYesD2B5IZikoPSWHCjUUGdMw71/WJjGc2MRWag+Oz0jgMNwDu3qinHD1cR+tz4j45hBM17cT301
ZRTURqwE+aQB/lettvvPXxu+au+AwFHgjV5x7EagA3is5M47TytScwJfB7SDRcXZyCjUlaNMrcYr
QKLQVEYd5cxr/zeNkFPSFq7bUmGJiX+CFFeQB6MNQxQ9girEogC5PnIh3vVkZOisvpk5YLW+Dgkg
/I5WBJXmBkK38UVfZ5WGjrPt8LDAElTTLZlaHk74govgMu8dcxMTVbACBdiKCTi7Iay1st1g7Jdo
2q0k86hQSHA9PwVApAxufzoCVVwfzF1tZ/Qgf7GGRaHn665iV04+82gIYZ5lpz8lQzAvh7z+q1oI
CFUl91JrTuCi1QnHaSgqDPCIahOz/YF2GG8DfrteN2oIi/FoATW995CEB7vr0e8q/nbJK3abKQgI
paXBUgA1eFQG2ekUtcva5fmU8jNUlJh90ikR3OA6j1C8y0V66av4Ul5aJ+mewluUWSfJanrVJys9
SekzwR+WDmUuxFGaMKpje4M9S9i7vkDH+DxSe2FC2iu4zH2Imizuy0JIeTZQJxdfKYEPXWjiIm5c
gdAYHQSqCEg0x2E0PMPAIJn/Fx7UdGVyITPOU68GBFzFrkB91/PR4YSQDTSyChZH7Tv03v133Tnh
NBnD2xLdtKhuEYEXnEQIHyqvzV6vrwFrSG3FLPABsP/1kkHU28Nvl7qSHtgUZ2kgc+eprfxCbxUp
YXXp/PBGu3wrpW66ct7WugxwjvgLoSjzQNeGeT3jV0MnGoevNkHcysjAAwlJolFvjv/vYkYYpm9B
OZln6FA45pW+SdYml4vG6LY61KS++3QJ44YSXeWveO9sHrq6m1dqNlW/aXoiXszcEnXCkWo1ioHl
r6Cs0OCJhbVK+ymznspVpjilZp3ph0GO4JmIKrWyiBdF3bH+41DFXNC7+Ww0htRyh2W/FPC6/vJF
8hjT2l3agd/JaEK3e9EBw73usFJZ+osPg4zUJRzQM7D6hfykzLFA9O4x2LuSPYUZF0i1AEwlrr2D
howd95hmRV3HdU5sqtHzR2gJfGX5Wj+eylIJl9iMOFOL3h9aN6acAOumQrKy2uAUM+hcH0v4TnuG
Sf/VTcDji8HAVPuXYUBf1r6CQEK0bUwubmbOgA9oPii8j0gK+enqggH5Si6sVrPD10l0Bzcjz5Kb
0z3IGbuypjMXhVnYx41WiUj6IGICwR5ravVOpOyY6ph8OWFxTFOTN/pqVCCjrtGQR3OuRD0iX8V4
oFrSmy3QU0Ntb+gG10krrdFU3esBJFlmI+iAnKklICTNe5CP2nFAeL5DTcpsO38puwMcDJ1KVqWk
y2gKOCDGL/YIDPEmT6iOxn2cw1m2CvaFKiKXHTCoh8UcEVFdPFeINtRjXL9RM9ER0qAojZekbiRn
BJqAgLH6GxnF5D+2c8WgUxvqANkkAll4gOQfUHrZhxJw+k13ICFiHMjU3tIptUYnSs6EC84ih7p5
gjhDazyqaJq1kREbtTTBxnE+7aeBcy73k5+7Z6i1VMLso1hdisNWXBFHvU2r21mKSluTDCPTEHRe
VWKoVgsjhuGMpM5yrKof+2omzRXrA4l2W42QNY6oxP4V1iuy7GwbCG8a5qT7ZLU+7PrgDVjY5ieJ
BbxSAXR4EBTL6e+5BDGoiSNcQjRevUI1LothvBtrAmhM1v6VkTi4KJ3HJ7f2k7OxCDdJzxwKUYst
b7AKNYVK3QyXbEUdRFhu2gqPqcaNArnswX5SLNO+BSotGaKDOlj6kkZzWGmWUBwHEchu3YkckVMh
bAEmTyusU7T4flr+PQNu4s+NX0cZeAMVMobe0jhZtneRMDEmPVhzbxkhLQ+2M6s8GVzut/kQuI+X
hWyqOb4k+tJlzy6bunK2zFR0W8A82S0yFhEdon3AM8Vv4Y0r7zhBZEuGBo9mCWMhXfJ8Ik6LM7SU
5peqlGVdDOS+UtRHNNjz0+xf3p13/qQ0OObqMpkTYN5c/dJ5Az21grllRDvSBpK3OYZQkmS2LrrB
8W1UvtjjE1n1NJyYsXbHQwEVmt3xTd5UDice/CJkXBrJyNgw1GiXH6JNKNdjwfRee2TUMbeyCe77
6ezCS905pLGPiNSJN0aCJX6C4yPP3SpRutNjC1im7Ts5LeDHBkQA7VRmb7IyazVEjtk31V9IlzD/
Wr43OToGYlRi6x5mVzhLHX3NwIAXfdKnzCAxvfRrIwuchp5j6tW07DrpOZoqRTN0w9gzAD95OOWK
ZKJmd3cVUz+7iVG1bILjVEEs8/nQzhzCbjNVr5H00JHM/W2kL8p9JRwYKAlaKWSdXq8KgUXNfiG6
d3sN1IKPci5IbSQ97X/1MMO38yKjLL0gVJuhp8Amh6uo5LRNJdpracpQrgHiQ2q2BNv0xos8nZWp
A0ZFMNN46egmh0+D2aO5HiI2BRmhJgN6sHkZHj9uZ8LUmWRSMDXQoAvRcUFBF+/9UJBzhRzsN0fj
/zuXtjfo9mnMu0L5p62UJoJW3CQgmO9W7xwn+aTwjSg2GHhb//sGj8qWj7SrVamilesTuxsujLeG
S/nInE4z9bToAfZ8bFFcC1sC3/X5yt7DOlfZr5Et45/7xHKOaBRmb9uNZjIipJmhm+Xx6dtJN96o
QAeX6grxAEMvJSTtPDhm5+nVGmE4AIx5F8ES6oCsizlN3KZeKmvxoyEFOFT0ej7R3h1P7IGNxDvN
LpY4Xg8mZCFZ/mBkPtpWEZHxpTmpc6EKbyksiuQFCWsPbX8QMUGTGe7KHFOO6i7NZbmLwA3EhvbG
VFHnUUY16kgS1CMue60AodiTYhgt5zqHlRMEnZd2iKDF+ytvY/R9urXivAchzHNkTO57nNylsjX/
+Ce+OwXcy34o/BB33wn+df0tlbC/CI9Hnva3uV0pbRz/TTU4g01mm+JIjB3BHNXOnlNSy8/p2+Wk
2vCX4MaCJgXqWfu3jEtgnZBYTDiccJ1Usdnzurjfs87alTMQ66AjNbgXPBx5ixRsXukpItmdrwX0
8b1ObXbHP62LBvt7aSBJNywCfww7WeJ6V9Pvm+YIuG+I22wgEnFhQPl7oItu0zvqy78zTAqlgq3z
f43qvNIunwiPDNBon09b7ZvPwHEav2C94s5hs/SaqOy2jiygeas6ztPhQnKdI9MeYoiESwCFpcMl
bDXz0OcUaaqOcsQH3kyqVU2YxrjWzotWjxuZusUcaT0ch4x9M/HxzlZOoSQxh4ZG2MCTk+wNmsxl
2LxejfWYp1b69y+fXVQw/dm0N9lYKjbqTAagc1ON2aGsyVJVjs9qHuvSeLYWXv66U0Pp9wIZW1UZ
oxOyzTMZsSI/RvD7kuHaBgWscr3Pfvh7Ue2kP315nHRSKPDuhD+NYsuYFVMXFLR10CYmhrODbsKg
jn4O0B9yC0Ei6lsF1ahSZ5k5sMUy5wgffx7ATHECXSoJ2T6/Z+b9pR1N78XExRBw9PbZzzbZaYhr
fc6yB3iAnjEjgJ29Cm7SLAwciMaesR2dAtuzqOMrcgQlS1QwgWnTU6xqmdHqs7kiM39iT9S2mUMP
mKuRpbakGX0BI+UjhLOiung/S6VMd85QLpQSjEXJtsUU+qwY8hk6QOKgx7Gmi/1dw7jjYglVWBFT
UF9KzVuKDdanhwJWeeB8i7k4hJGn0AN4/gvseDGirCvlSQ5m4VcdmnIiNShalFTvm6JHsRM/FKfc
9+Sf5JhoYZZHuntWaM4lutgOsURULos/orA2KrT/S00PIwl+v9RMk9WtcEpc8L8P/nTKsQ23OjLb
/beKRRr5v5aSa1p8hGGe0k+y+UcAIB3M0NKNf6AjMBJuECmBpyg5Ytj/i9A3tA4Wm3Ww9ILizjUH
BqOX9VGxuNh3PcJR0/tZmwL76VyGr+9BmijdR67XTncvpskzwj7KXK5V5COibXd6svygUAVP9TfL
WbDI34iUr657W9D6hOwVV8G8oWFUXr/iOduw2yKGybsqjERutZBEIDu3/cqK1RYMjNbUUibZhFES
6UkZF53C5CXwnBLUKNud3tdCkhRoFg2KosIdZNpNDHS76djpV4i3hM2gIqX5K3amEz0fKEu9Mueq
ppexY19QZqmBBJTEnVuLz1B8/ugN7PzaP4NXex3d8mGjrbiTp4QkRKnVZ+GEM7Q1PUUrqxd8MyVY
vS3VBBBiDyLg/FqxJ+baprnmBH5+Mz8toDiMsx10mNm9VoiuBV7ENUKKwqd7TAkPCSEK5KKdd3Ju
e5xqfSYOs5sKz2aUR72pJUzl9Z9uoZI7U2kRtj0lm8Xe82kx9IoM1tuIYBmMRXnZ9XhcPRh+8miA
QiBndWHFy0wQo53ZTHHyIlOQ0ig+MHqX/tPO3FGNScc5nxK8z4r0dWMzFloMGmRIJYjpAnanqonC
oC+xwJA32ThPazyXq9nJna52pUUHnY1fCjZhPpSxFXiXk/qKHGDbn2w7vjPUbhnu+B4i+rrEKEWV
LyWePRF2SseOr5Wm9NcKoKD3mF+Tzsorxf8A1z90s+ORjKCl26vDNCbeaHsRJxpXWbmGfUZgVKPJ
1kfPaNVAwoIzYuqhsVyDhnMpH8+a61cbrjpjwPw1RP7QsstFMRCuCQoo/XPFIgubeGhdeFGmSkV1
Khp6Ay5yGOFrxIPE0ONSbQjL1lk56aimiVfZ1Vc4/06H+qA2EUaHFnfTKqHC9qhqVsIcZJzxEawZ
Y0KTxVsd7U4bErWqcUFXWsCRmtuxVIPcZ+dt+fhgZ653r+X/lu7ZXHaS/5Eek6AvIRLOIzu0JiOo
p59/3gKRt9N7WSIikNEehS1KKPh8slH90YqgUxfDDcHnh4WHS9J+6nP/n/MJkzWeRdbFBq7JVxEW
w7mF4d9n0hp7vlNmosutQmvrys8Y/KFEjdJU7O2Cu/zejseHa8hvzOZJRHKXqsE9jn3Xd51tO+pS
+ZiPoEVSzYQo/f2fu1NnQiqYagfjZzYillFErHN+At2PVW5/12vDT5X/Mo+D5fCpk9c++T0QX8+C
EwvxhEzokgN4wUrdJx16KuK1OCeRMFlm3kMXhKZI/8OZhEBOCEMUMkz5NI+hxOQs/YIOjCGNfw/5
O+GAIWLfKeLT2c84/svNqceUFz2byNJh7UfOSx0VbtQBaS3/C3A2YGoU17Wd7829BIq+M7DxdXlp
wD1YNYmZHQDYbxHTLGPyrVkaTF+m0NRqzKjOpg+MMemO2ajgJfgswgICg2wQG3x4c24jpQJWqzc7
Z9B/IcBDJnd/HgHWGHSvAGmv9uIGgQj46Y2eWmk/r1pVnKaTaC0Hoe+On5oibvTVT9bD+C6kH9pn
d+mkqODbIYofK7tMs4t/LC6PYIraGD4JwwAK0PM8ZYONykjQyIKJUlzVevtk7/wlEpEMVItkC36e
U6+FjSfpzYGFCX5Z+WiF9rKvaB6uM0wnnR2sVU/TCAJlsY6Ehn9m8SonY4q5KhMEf2szv7PMJ+Ow
UvCA7cA+GaYhq5V75R7VBcNL6rgPvZBTRAv5IYrSFVD8b/9boLFb6r38D94zMhOLp6DgCd4CST5z
GtlO9KVjh3IxBw+WiulveiSuix79wqaCiTcF7MTyYtW1WqANeZA/Ed5hmqIdpoJo3i41oDzrhonO
e/MPdtofl+dXneuOdM82YfCk0ArCfcBwBW5uelPxYoXF25+y2RUFgEBUyYKOxZBO3/rCahyqfWPG
p8XBaccXpiddODRFpXFzGcC1KVcPuDKP6TaCuWRUE0VltrugBWPXcdVDutFrgiVZp4/2KuJ46qbd
GczAMKlM+rAzwcxGd5qHFn7jTkcunAetLhXq+j56/vmikVe0ncFbK9o1yadZI8gYSpwl0yNesZat
9cSukVkswbohHpfQ6kKQeQBSeyAojWzMhNwZBPOjMKCsCOnyyXA2o04z4inSZYeGFHte0mXK2P2Q
fnnZRmuDwFkpPjBTNnmIXBZ4qtu62fLMvkeYz1s1PapPLuOWBtm9LCGjhQ3IfBP8JLn0xgK+BvET
Uq+vCVfRutsnfGCyT3HOlqSaoYiYl7bjUKG0K3uje9jmWIQtlbh7F8OFRA+4lQ1MDOn0nwTHSDqk
uv/bJsxNnxTcO9/tjQ7dVwkkqDZhqGOHAnZabp9TDRwe3To3s8ANorrzNpiMdJH3/ghxm/i0tjqV
sg0vm3klLHbg46NYyr0jxfPaSAQw4uW+uze/yzc9aLnYMH+xHuR/fD7H2y09QWfcsP5qSW6utMYO
+zf6xPiGgfj2z7NJ2MKMoxq/PUAEXuuNg76zRg1CaQEVdqCgHUkwtraXy9mlMfX2dl6dSq0e41K5
K+ZH+cTnBJjOgUzpT3qJMjgOU/rgFC5KL/cgFd65an0PhrHHqs6Hq2AADOaPyqmAtC2VhEGM9NkN
kisUvXHrZKjHsSDlkLvUSwggB5lD87jXKQKjsPfMkfnLFSYrhHAXfL49kvyvgkcuvoPeN7YLaOOk
ssj9XqNXtVFqJfR3ZOCMpp7BWlMMk8pZ3Xw83MqiozQI3gnrlPLpQNfKZJZmQNGL4YSP11vjGAEB
dKRQuhA3lyHVtAM3X2VYTTdpf5xDbIpe5hY9c0S36ve8++wBAyo1rGxkxdXZzUVlFvU3nma29TGp
gHNTl/DgOI9OSPZ94cAn7TGckQRp4lNHuNLPNPdXQrp+g0b1sPpkJnhZDOqeo1A+8QqZzL4f+gBS
OoHbGaWbnM1OgL/o/P6nOsvngut+/Xh42uotEUa9f8bno8spmibdXIA/0GBpzACae4N4o94A3ITw
Ec1Y+xmL5J6gHhJV/Ug9/SgSeV6iLoBPaxzpg6K7w14H+okkQNH+7LEHlHAQNK8wgUg0e649fP5/
2BgpuWVMrMKMoOSIf5nelU6Oeo4u658hEUU2lPfQJA19LN7OeoUqpkt7JT0Ql2IX7oNOAVotFsfu
6al6nHnX3SZb0dpK1RmWCv60b9xxlSYS3ATgbVXtncsHLliHOYKWTiZxOEROB8zDourigSdyG4ow
OtvDAp2LowGvVlErt/vbKiESI0mAfy4QhSHqI+G+PFOY6YtSQ83QLYgOnl4bSp/SObwMwEs58Sni
eZnq1nwxzvz75W+rBUH6aKBN1IC5KoadNEltWLKqaVCZiGjOHEbhGv/OKjmFmOnTTtdoo4J0UCOY
7lPrzW60QtJdtXCEwfn80SWmpyTpZokpORVpMdUP6rvKeiyOdsYsPP2rZZxQyKtGdpo43rniB9AX
5q80RoQUQ0V0q54XOXzLGqxhKSWOQdV3/misGpm41MKMXh2X5b5GBXi/eD3eJw8WIfFxP+87ri6b
RgdsxTAMFT3+oQW2F4zj4ovP3Gc5ytsxlJHuEpaBnoCoPDZRANRW9mzTSXHW1SVouor1DoRXWhRj
lhavoCn9Av9keQMjq6j7hpDYx/L9H7+pWqpyza9AezQPnywKmXYOZP3FxERUXTs2k4r3BG6YQv1n
/EuShYv0KBC1xGZvsUlKIC0VonIPOcokQWetWNOjC/wAxEranKa2nQu1yeenQa5c1aPLUfWKidd1
gDyS84yWFPP2vX/hKAjBZKecu2yphgBMCtiIH3DryYz1RyMzHkEzKaJ7sLs1qfpKXEESQv1Hn1/F
rnQCjqS4Hq1NZSjTcC7hfTTv2WurQBTNHVfLs/mLVNjvIP/f4aOlEWCHpKdMQQ96eh0RA1TztILF
1LRk4opL3iHXp4Ey+unouZTHEzX9vBm3Dpepb89atl+wGJdIUor3AQYyPz5qFqE6itJm9vKtjGPA
UcVV9ByozVBJ5Hzi2h/XV4bzEmqTqzZIiyErEBLF8GlaJOow7n2/qnsNA+38EUil11DxnpIe+xrs
UN7v4Z5H3s8Syk9JCagvZ0Y0OxPdVsNpF2QbuLOllFyD9L42VSh+73ypSfdIRHFYaFv2nznpa8H+
a+ty9GCgPcUQ8oxp+KvjqY/qPMPRDhwbqQ4smjNXBTlzojAeI7Yagw5G5zbNckHulrvHuV9vYWHF
vQNGR9uUuo8E3hoJbR9X7xKGyLeHYAIdYWUZv0X/suB9QvE8ubd1njnAlAIqgfM6a4XcSGiPGJzL
aEavnXpBnym0sz1xgLLHDv09E1m/rNK7EhXfEeGYI9Ryv6/Rl+JSIa3zg7tqdBaf8PH4zEF5GOVz
FqlI0LbVG/iZqilJgdPB00jJFsHYLvFuBNJKK1F2vp7DU42EdqikKdt/QWr0EO36WdrfAzNFrekD
svPFWFXHJ9fyWyTl+hYjiyv/ImMbJ1SOLMLjT529VjZCSZsI+JAqS93dmdBEbpgTgn5udhkmEjHf
Mad3E8C8peH7/iZ5C1G5UaSHiGi7o4CCZfqQL4xzIKeZ3Tm+Jigdynk72hxGlWIQDeEamxT4wjOo
s3C1SqP69XNuW642h1O1zqGea4k/KwYemqUFEiijUUPRmZhsbmF+Xm6ACA0giCEbfea36FgdC6IO
AD5I/DaWdwBj9GNoeh0sTaVX4B4pMJERgszaQeHiKtX149bQATKW8/S8rAotYa2rPrkYxfwPW504
8u5QP/vNYYgKy3wsqgMt2H01S/n/Tzic7DyeOxdzYNA0AGlYgiameGPz6mWstD/T29/eun3UvXcW
pncYHHidsYRJ4lyBg4ACsH3FOV+l3F3EYOSQkx/ngpoLqaPZ/bx1s/liZwNngB6xJ8OQvJchw/2x
q6AYal5l2Q7UHYNm4T2vO09sq7JMs5IH7T4FjETUjx+B5qfjJ3vYL+A9s6CNlFw60JKjKVkYPRyq
tZwUtEU9e8qi1G5hQ8lAkqxdy2wPd5wyvayhq+i2JXL+b4HMwkYlkbhlH9EmcHO7F5+OL6U+C+VR
bEj3BEHY4bHw5a7zLUo/JrnK7wjCuPmdVIFNAYa3Zf9JioXW3XUluO0tkHWAa7Ca7iD0k/TZsFKJ
Z8P1lhx56SjpYinuVAq/oWl5UVHdmu4eLNWGEJsb53hytHPnbkBPaQMselZMy8WD71Zcd5Y2lc5K
WZUhkQ1vibaINRow1MWUI3CJJh+uQj/oD1n3F5N9FnPQDxYVOmejQzUVLv5c0OBDCdgSzs43DMnW
konaSFlWlyHCCiI4Rajl0gQECJZoda6QqYd3GE7OyEemliWBV3Di9sT6MiAdetMdVYDp0FiOQA7D
DziatJWiU/AdLuX/qVX58FIGG5zmmd/ppzdZKRMSo9xPJJlKVyBawsjILmm9e7cwXJ24cxnUF9I/
CMDWX5mTjiRh3LdmUcaysAoAnozEYw7U0A7jZIFp0+UYjb5Shy/Aa45IV4RjpZq6Gk+ADcmPQ7xH
gqdW0F6N/9UqtRtBatoQj6zWrPPOPrnLovnJYiWdMSYRHWjVmzfffu4d/F31EHcNy0o0m+yGTg3p
HBCFnSHYkI/uhQL4qTkrgePUTEAM66TzJZbaSzpAp7LOGVK0s+YWxOJtSBnqvprafXYdli8ITOto
8FtGQPK+X1DLAVjfRRTbZYVNC1Y6Te9Cgj5j1Ai0sTOgDQG+dLwPSfNVwDjKoVh1kgZc/DOoYzs7
nLEZQDU1AzVbs4luI3jzFiDO+WhuxD/zNWHCaNuMhuGfSCs/szyqow9t+n9IEJjvR+0qnoHEfO0w
pOu0OECN3Hliws1N4eM1XnEGpiw/iy0Im1WJd5Et9Z/V6wBu8B1cKeZ+BDyrGmtLLR8h7UYPIvu8
Ii+sNbUBPvJGWfHG0VGqoP7InlftqXB6L1dwHzhCcyaBXjpU3PHtwJmZ3AUkl/sf+3mFx8CGnGV/
qOsGU2JgjVB2xs81NDtIY25B1E+YGdujNYDlI9mInq/VUObDHMcptH7zruFqDagNPw2r2bZhP+vE
fkUuM15fgteg+k25meOCb9Oi11Kn4DoWTi15c//LQYZ45LhvX3n3g/ckljF0bBQ7nPH8UEm5H3rV
We7N6zK0RZJB2fJIKoSJ+Bd0yJsUmMSEfS3qx6FVwlYQiK+nB0MMQwARf677i7ihYYn1E2FXexnJ
4WCKAZBJMWfo6lzaSoxsqD6DRRW4+GHJN9s5+A2dhOprteB9CDi8g6xdmeoJnL7yOmEAToz6Q9um
2yNMSlQXINzstwHA51ZWJJ4rsHNqQDpAgjhrBDqRsPIc06DclfE27gR++vWBJTGqavLSIYqEOUJ8
WlB2w6FnZUXZNgHGxyNiC/fUXnHbBTFHpDW3Vd9VbXa7cJ9yptuXANJ04oHOYgGbgZaADpmWIehI
1GvPw69WLUjbv05WR+YqhwqfV7VcFJnIMNvO9uLFiCq29/6ARgYeebTReBlX4knJBLHl9Gai3GPl
FFXQT4cb3GgzS4R2ttHdW6dibrzFGJi6sBchIL2Zli8NxcpZX+OkuqD67OVYdAT07bInK4z06gJq
H6hUO0RlDOdd1OCaVwuLepUg6XOuhPROwAUsUP9b6z7j9Wdi6u+xeYVMFKnVmx4YPY0BQTg6shUR
gd8d8Qpr2nAkFBcooxT82t9vuPIlPvnzwW/66kxN+v0HQ2ua7sR6hoymGbvMkSchikQFiIUne632
A6cURLYT++v+0df0wOaRH857DFhxP+nnFWMU5wX174G9UqiXer9UtvTLWU5EuLtl0LDiy3GKmhKa
qo3zp8AQF29dTMYIjyLnM2io1SPYUXIQ9LIUCapfQ2Q4snER/cK01MEN6i+j06HdszhQVlGyptzd
KoePWZ33EgRI3/taeRjV4MZu86nuz6XzkhKu3z9zaR9mVIGKirdBT5fI2XMAgbUPBNVqEdyLPyF0
R9bgwyaFot2b93gXT0Xb9RtLZQWEmYW06IHTehhffWULV0YizHxrdWuPQ5GGNOdJpM+NQ/mGrzZg
I2IEaLNFjc5JakMuvBAlnAQyZNCBczMsXpLROTVl4HmZsW4Jx8vc1ntjBVQ/CG2MIjOkaSbGMitI
ZH/s7oh58do2NuLvryHpsQ2CnArMe7mvkdjqaKYMTJB4BjqZf8L7N04HBhBN9YHFNUaYMzn4lJMY
UzoTho2pVrqqTB7Zfg4qd4GmSrUryNPFFFXCxZ7IFgJqzyJYiPdpGmDZN0sviwLZhr5p1GwBll57
nhy+7xBwbLxUUjnLsZFdSPlDsrmOquo4AMsNDof0RYypmsfNWg4ewxiCcV8KHzYDWZGxy10Pelts
s69/2Qkr6EwWoGizgwulDFIVJV5x9bfYpHe3vmpSGYMfvB3CCGoAlicAt96gfibMEB0v/wtXCQ1M
biGH8n+/V8qFwFYawxa124KOiSfZ4fcOnWgqk3s28Awm9J6T82eJ2t5Wf1khXZJ+ntBHEGRX5k4b
4tEckIMyptQ084WjRmtbDs2MzVZa2Lu++MyqaZryFFf7cXI2eomp7yKXwV+3Bens6HOlKqXcEqmW
vXzFsfnOaLgD6gTflO8tJ07n7yDvt/GwrAvDt4gdBvh7SoxWTPB64X86X60AThD8S9niHknXkunI
s6pJh84WQRWJ9JC2ICU3Qa0DFcDLv/RVbS5CLGkd8l3gtHBvBpZa1dxxbnkGiumV+3fqSnIO+oNH
OpGaOb4lJ1CGOzLqn5aBlEBeJYjWXAQz+VJglrQF7TSwZcoVsvM0ZYRI4dlXiIk+uoIksqSxIfL2
kmv6zVatgeKotSJ/DyedRp1k10TOb8ALgnTFjNIx47GlTINiTJ6dZg9ZT7ailfAVS6w1By2hfax3
jodw+awAAudnt0QrSDwrJ0qsvrZREFMUzV9IbODJRxX3XFEPowiNRtbtLmTpGc6klFgNIXEcRNWY
HGuTRkZOl8fjOVtlLi769G3tU04vuLfv4a8EksjipiHocnceJFJgty55iLGBVD5uAvV3vJNFLfHL
zgILB6gwFLRKtf4h/6imOzNvaYRl5/tCwGMOXA0Uv/ljv/piZmfs4VBg6Xac8dqhyuogBmfANW70
0q2AJW2sw10HDIc/CcxjXFMXXu7miSau3JDF9KiHTOYEqbJ7yjIMo+BJbG0rJYSVIF+4khDtRGBt
tXyMr16ghHkdVKbaipq12CuOIcgfoOrdhJVGNWyHx2jfTosyCUOX5vYgO1cKz8jDJ2Q3eTjsVV9B
2LuqiqeH0DdfECbhGoZDP61MsvlG59qTrNFeBdBTkZyX/qeBtHKeuv3oM+fJzq+v8q8R96FnySSz
pnpY6w9V9En3/49vh2364OV9lSt8Wzl+JWV/VtJBua80vBEj4YMNAMHKxw+hl1UKHEEpWw+dwyZk
vM4DlI7+n6o/j9zesn95aw47v4eYvwzogxtMTwK8KD/wUftXX/uZeBFfrBa6zbIBs5OuuZR19aSm
dXr2ge1qqmB/TN4ih7uSlYScZF7iaumbK1pBbgEyL/zjacdVSjhVNVRLY4AVkqD9tnpw7cemy9+8
zP4FMDIep4PfvSVXFfXYdxz6X6M7zAK8YqUss+de9v70CO15KDxiya8sjFYb5QIZQXKtzQ3wTlEd
Qm/3g2puUPvsaz3RuhjBTANde1i5HF4SbuHil34NY7cu87KskHcV6ZekLyS2lcukac8hhgsGPFuz
GfAEO0xyl72smVCHzeJjlyd5Q5nQ4QOeokY8DmUDahHJI1l3ZXaTgBfXHp11rvWSzOQFL+pUq3Jt
v3gkTA6PHe5qRpoQ60zUlHCxvpVv5RK0dMPO+hlg8qqO8IHSpbA8YoSm5jowscR4G2tVJIdIH4q3
/KDiQO8Ika1pjzlb8aKGn23VC3jZ+6++TN92NpcPhPJsAzTjTlARqt1c4y8HZINoJLGyskyWmr4t
NkN2HD0Cxx9EZW5jbJM5Bgtu5ua7PqVrXmAF3V5h51ArP7nTAQXKx8owAleMaRHFJCpXRX+55U+b
QCTqZRa/XN08q8bxaJgPLzps8eFQEy0KisGoH76B2C0p3JluNHqKpkLLi4Je8COxYA1y3Osy78F3
ZfvS6c0GxmLoiOxsyUk611Yz9JQpJDaHMJ0zpLkzK47/O1JMr7KCdGbL71NVht40SzMcE8z8F4lu
qzBtR2l6S93esvJpp7V5Escp2+Kos5Fc0/y2OJ4M/xXCfE1HzeJ/rTBSezYyK6L8fAUL6M+6f8fo
4H8ASEjh/BgXRUZHJV5OcWVFLqhkA0r3415xshkdYnA/ej7aP0l1/NhiNMgQSJtw7yeO2FwjP6cK
qbK0inZSsvMpQ7olRTkj7leSxKQ8/p64Sl5WlfnPoDQlRP7hfOCY3b0h4oxGENBYMbFLbSYXvptf
byHzN3+O1d08gtnVjF0eZqPQOsDsT3YVHrXiC7qGzYaQgNdqGzKmVOZjt7uS2WQjzrPIz28Xdhri
7Bwl9kfWy809UgvQ3kE0vmM6MYC0VHm5OewunYUixBPDf7X5tRmQH7DspP2dWD2WC0U7aBbh6B0p
05DtMkEhWjDunSipEP3q43PoRN45B7jJ5AV6Whu37xk7IyhOjuxr4N6iAhdx3HuLyaCd3iRModAL
3LR9KKyf3Tj4L0bO8SCecRGLGPtIWvty1+lt0kUMnnBbh8NNglNT+qNdsEebUe+254LvwcxaHEI6
f0ZuGYBmdRftAlL7FTtS/mtpJo+0eLe1ckrQtMcAcz5lKAfBRnC9mlHdpt2ZwpQ5cPs5sssXsReh
w1/10kXU0R98AoweK5/057V9jJApiDwltDxuxS5lqixggZdimKd2Bzs0QuGjC7ea+E9U6J1fIW6k
ERf9Y/+NLFpcx8SpbVxFYIBbMaU6URB/SKL1FOGclZGoZwPtoLNr0muRgAkVbpE5KG9y12kt1jMr
Aomj58yPmNqVtUsJoCD+36Vn12b4DKUN+hjwK5yx/YoxSQfmq78g4ymbKxpS7i6zQGzHNjJCGJ10
fcZrAXCg5HcPZU6Q50MOBqREjbjxyRdRzxkPd3AtqK9N4Y+VfbxiFcpvU6zuEeKpJHJj+J9PGe5v
VrY+AjNSbU9BnDHLMiCOTyoBEBRX02Udypa/W9F/Gw5RGiYDZCp3vItVxxe1bnMm0W4U995oiZ8e
vOiaaCmea96bg4dFYCkKIfLqJcDeRjIDa4hXk7EDzTwXvSpmd4mhzRylpynF8dmFO/24lZDJa8bP
+Zke/ho+lB8nicwt54V1+S2kcjcgMOjueiXHgL8nx5Z9/pX3d75HltvDdP17hIZA2wetwM2LyR68
cw461IJTtxfMrO9CYfIADsv6gNXLGovXC4KeozPtJHk5T2mCMA79uUM48TV4ptayuHwJ8DUwfept
S3YuoKKNqKmUkJzXQ5KKZ6T7WXmAtniKnpnN8tOslGk55+y6n7KqfhrRq+ly9gqwsGLFTlNP119s
rMgqDQqQLpbJgC4MOv7KX/E3m9tdGfASMoIZyPykIcswkt8DP8zV5UbdAwvZxVGziNFXfZWgBZje
aA1mdG7N/T76PxqhF7HWo+dPWjhcSFgiRJtONKCjjGN4qeRmILMrjsDXqcAP2ft/89TyhhP06MW5
xGE84SDjjGrQk8M62/pR1rFfZyLVkCEUwnQWM74AvDTuP7A84iByVZX7EdBqpITO1B6aRAQM8swX
n5sShhIHRCrxWHXjc+yvRPpW4yff4j7BIDMLVRgwGQ/IJwdhRva3GyY4D2svk5UU9ovwuzzp8tLB
UZJ/B6MAlujM9F2+e9JTRMbVUMcrL3MexkDL873bwNwDUu19FO5RRB1h8WJYyDGWs+7dISLbrNUZ
NjwLiGMt/EDOfodwE9wOve4RnpMHmTf2cPIAWqdJ1kYIH8gJaavz5E5TXsrPmnzU6vPrJJo7uJWr
WBID2gAETBNK3HUKWB3qiCMpYPcfASQoYJhROrzlyAcJRB40+/qlXN00IalNRcDaythd4/HgF9Wy
wsm0XctdqWvoGNSWkCyPFHV5ItCVA/cPxqdYP5D6Vvmn3ttVpmz8BMO/e5uq3WsIxPffJLhA664q
clmkxp4iNGIz8FA2fp3jEJpcoeW+Dd+r0jeWe1XBnNQLYzVcKaCNTHVqsQaT56kD7ef+wPE0wdw6
90L4+RWKQCzo/J70A+qd4Nu+z5s6zi9iuOdyOrrVz22KJP4b1IYFL72//l6brZBSMkT9fFt/XoqI
hx5Cu0P/J1do6cBp+7H7n/Z1rl/U4wuvupunkf+iyTAemeAyTtPgH7qTs0LaaaY6A+Y+/9eUAp9W
fAwnIyxForf06F44fPv348uHESnefQiZl8vIPANDrIYJ4ULQ+BvoPraKDOYjv83GiDQlizL4GE4g
yktwrMxKcNOemGQM9vxNoD7wsfkDYq8EAI28VTNGUCw74tcqbEXCt6XpZSlEFqbXTbFOymsTQxTD
8P7b1ITzUdk8Flp0nEVAXN8Lv6YjfGSk9BweaJNIiSLXoZoGBIYtUrj6xjnOY1TUZz4rl2HzzCzR
brhNcDHAcqHbUXMlFQjMkGXpdFl0M7umqCiHvK7alrsgLQ2vkxO42fzpMsqnTtNtvC5DXFhuX7ra
E+pEudd1uXTyzBYXhjbUc1JD0O97eVjjvj0taqm4D9y7ga2JAQ2fKlcJ7WU5MTWOmJRELCgX50RE
vaVd+ddrBikLeH4U4pgWyfL133lIo2QOxrY9Bf0jkuUffUtkaD13CMESCjSA5u/yGmOab5anK8dp
IdnMEaVfoeZEmDRS0bGy0XePk7d4hDY1jXrk6xDbRfg4X0A/tRigRwmYJcacngVRJ7dPnas7fTnV
cO96cAjXbDraT9BTvCdT8Pu8Ry7WaKefDZxWIfhNyhnbL64Vrk5N7VdPn7/EN7xTnOXBlDwvrHNV
H7WWug+wwwTChm2qEUtqZL9ShUBy6q+XLlUoRetIT2Lhtpgjs/QeuGbb6TaQYc2LjYMNF4AOX4Ac
k0gobRftAFr/q344yKN2Sezs5RdjHcvp0dibju+dOTwUqY73uUfWblSWpV36p1bCmqJ3kMXP+qh8
OS5SHcSXehtxl3BQf/XYtlbj7sO44a2ZEIsjIz/5qevK8qbq+QBqfOQ6ClRrwUazQfw69/Q2+B4y
E6hUjuFuz4LkkAmhPzEyX8SUCGZsFceueRiCQ9133QbCqt+949XW9y0GbpC7xUSG/JwteIDaWmQH
ghQUk8Alu/JnRnbjOOB9fqKfHzUhlRd0Wd3/zZalE/ksJii//5GiyFq53Afc+iHJP1mmSOq8gZ6e
9d1IGnrcxn7yTUBCmYRh7e3bY52OKnPotHN4WMrtmUORUgODQgQrTNA1X7V/XoazlxpYIlGwUw01
fcMIwogaoXOAw3sMyAVqXZhiFOFdJyj6ifn5+DjNACmgTWqn6t+WHmt4h+XpTCYsR4uNsTvjp7K9
ifKktJCJC6DCYg2JmQ1p4r04JJj/8ESo3u8orEoiATufWESQ2ZPaOPY452Q8kX8nkGmzrPsMFoxb
M8wsUEb98+0M9elzLovNJxgcp1oua+ATf6Aeaj2Lsnxc/qlY1ZjfCrfmP0sNUgZ7ZobbJnCLvdLw
pAQB8j2G17n26JJoaQXHgwNadHMHxwA0Q2653XMpmwb88ctC7Z+BH9dSJibKaVb7qlghlLnC+rqr
ZAcROkVkk6h9lROoG5cB4si7Cb4+vMlz6ELHwZRmdbIkodGpMjuSbEoaTqKdNfuKGv6aoygcbJuD
lrsRaBzGW5JI58eIzhB9sjEeaDZF2rRp3KvwxHT8WL/lFS2GBb+oS8n9uqDJlenB2eng8lXrf/GP
t8JhtMzBrWGD0cZ0kaDLG2TAAKqZbNbcO8NNzeuLqZ9gcJI//rIFrmJxec+cPSvZ3Hao2paOH/wz
6Ad7iw/nUw5wvx0dbvmjASBqmzssxan75EL4rC9wXvbbjhQywVXaRVS3A+GbnABG0xeWWcyqDibt
7sKpi5yxhOVKAJeQSRqyEgPiAUgaAMFTsCjDYNPi7SJG1P4Xp+uM4Y2/ZVD9HToNdItVy0b1bcsr
WXd4Jhxmmt+VMcIRAiDj0rGph2KPnGzfRyN/94eiPO/f5UGWXrnHPmlZN6TPVBfGXSFSwHVfBFHD
DU57XGi80pwQ7BTiwU7vCXKIceuTXAJNhHBHhrxeoRH6PCQu2UMQL13g8K0lTU3/n8RU1nbPWnwT
edHY6dg4SPRUFRPt3wz2Xz7ChuWnvpUv1E8mvn37bNuVUiuuTDBnsydXt47i9pU0c5XXikDQzKUV
FSu/Tpw2l7LHwW7uNv1ACRbiMYpHfYuOc0c4sq14+pEQI21XeXOJQ7Gs1Il3eQWjf0ljm23fawtV
SSzpkEVjNv91dC332RioynQZ3lb0uB7typiFDb1+NyOZ7Vuih+OJ2LfhyxpqvIsHplLNvyfHZnaK
3UpxjMzZpy2QUqEE1VCiptddEOVWAt4RhQ//6dAcVbb83a0xY23UobBdN3ooh+E/tVnVhI8+2foB
vl2Mx1PlLZHLnXGOZlL0T2k5uAL69GtN+tk+9cxy9DGchv/eexXjQ8MUoagyvGAuWTV8dVbJQlAR
yUBJRalGWlq8CMQLf9cM5IFW4qpmygjJ+E+bsaIMW4LHK/yQpPRQdcn0EWnc5Ay/ZDY493It71Zi
AbrfbdGtPt9xMQym4yqHS7Q857LBAer3s8qR+0ORw2ooeoxpSvHMoXEKGFdVSESAz2RfhLAde/4d
IGrvPP98oT7hX22oD6iusUGXAPPqmwPnGeIY4JVA6HsNRclDmWnF8Pm8RhJ0XgTop7HXmV4LOha1
Zr/F8AH6Zu2CHZ6JMwKdLbIgZAR7QaGix/PkKVwdbusMKzcbYjiYiwgUiHa7Cm+8HYdX4d8LdZZD
4ZxU8Q/cN07AMhawPtAM61IBlkywhg2UWW8R+aS7ZfoHDUA2CSXenSDSScRw6c3WdkuwvgzRpP60
YvS/YI8g7mTARfBx4jM+OsZsqUaxs1zJ0ld4h4DF8R6eG+TWPiPmLxBtD1OOxmtOFDeNmFVLaJXe
Q0uUPVfknLbKQsZGoKzIPY4zIfq/UxoWr/lqKL3aI6shNf7YP7vqqg66MWceCIfgltAjDrk+M23O
4+KUCUMJm5I8J7qyFdj8Sp0CXYxOtP/SONBVEXHCahSCdq2q5sy/C/F0dQIPBBs9RGK5WdJMXHDm
SRcHfXJMU5WXxq6VRppPopkq0HEYzjuoZ0YUbthLDWElEUme1O9KECMUsTl2nA4wW4SkcbjgU+X6
VTo0yNN/6aFdcl9y/pzaBh120MIrvB/wJKPYqnNMRo/k9mXXYxer/UQzgUI2zM/z5rMEj/Sf1RLY
TAGYBinLOxDCuy+nZo54adeuhjFDrNPJYc7e6vmVlnkWYaWw/Cap+rF73H+8rrBTf8ljlztGf59P
3HUb2UP8sSWdSVrMAjyK7HB9ZSn+L3xt5W7xmdqPo0UYiCgc1nJvOFfNKg2tFywbevjr/dx99YOq
ERJa0UvNDOpXQvGhDL5R8zuiUQmuWXLF9hTtCvptdXaZ9gnHW+WEytTA6qObzh4APNq5jmQ7h5Sd
YDJbolqpHV8t4ZZKQDlAct90iGqqHHWmggCPcETTancvXDuU8ZK0oC6Acs6Hw+t2aNAIZF0niqAe
VeIugNfEGGK9k2FkIzK4AK3UU83TI7Glc4phssM6tw14z2u5LDDBVaoRdtvcVFWCZroW0BaXhXcA
Q+UOkhoHtUV3xXU6sf9B0ENkeL/OjgncGgDw9L3o9hQ2H1ab2WVfdsWm3s+eJvLZK3I6D+6JZ8hI
tyR7R6HGZXYfiA9vRRs4BSaIl8nyk8GtorJDJ4hocNRY/0CqmuiEvUMEvFrGWWGTZ8if9eeqA48q
usOa+U76M3YmKlOOYr/r52bKZ5Vg65S02a7+fEBeTDV77fXE+M1W9ltFFZIKI882/1kQR/TuoQ2K
XcXwPyRZJN28YiTMR8gXErv9+cEB3ldoQUddnsqiJsR1u0mCKrEgJRROscwbg6GX6J6Sv5/xK76Q
MPhAbEq6T0oJXoU0Jqe0H0a/znGwEUg8yUVyZ24/2XS+7aXDKNO+N2vaIahg9EDx6u6O4Jv/ucRc
qFj8ibJAuwlzP8BuOo7lLmMamtWlrWLY9uD4cv9SmcC/eU8G1HKlpcRe1tDmtEQ++8/8oS/aGn0T
PwDTyOf/U2z4T/V5jw4Ky7tBhGM0d7lCmQP7EM54lC+5BGXllDF8d7jBSu41l4lwoUNo+mFG8Qi5
SxWUS0+8BeNMFYtNqS9VEOMTvIMJqSvYMZGVgFWd0jC7Rbuwc8PArELEAVq17MAH4sq5NHQNuLnw
QjdfW70gvizLBfUXba3+G5mJXPORou5iiAx4R+HBjsFyMa5fbU0YJoKHgsw8ORRJPPrYn3peiiNy
bhe5c/YeZ8RqmutFrLPEmUZFgpa5m8gCc7Ai1cZPBJfGAmjsDxTAFM6qtCONYoFrYErlQqVqoyG8
8CLpe61ajjWQCksj3s0PjZvSp3kYMUTNGP9nnqTwRCu7B/DFESCRg9dp68BxGhb7r53sLJS8CG2/
8GHg9nVGqRm/YnUCy69BdX2N81OfYVQ8DT+XYgrZ/mXjbIgZ702p2dgzdIUKrAefThXcmX3L/bUS
x6CzvLFxyWFmEsNxVGAqDaeZSOv6x4oJwnHlVk1Tb/SUSfaiy4kiQQv5GLXVPzKHcAdOPQWrez4A
HBZA/GSfib4ibYzzNPGYbVsipwnHxLLbQzHqlA8O12NdUNNjLmotVMIns+MaSjt/QiS0aqYJTmYE
9gKFz6oVQt7R4sYSwtejDXn0ABJ7wCvnwoPgwSj4Ju7vMmLGQbhS/EUpq8iE3WqaUA12nIfrzHG/
yYUWyokfUglQyCLEGnz+4kie2qViwKWcBTOKiJwp3VkTxil4QhbF7r9vydVQg4cZvvYlRvo/gCrC
2vkIHEQboi3S0kc2NSYBiAhPqbKDjy6zLVH8rnzKhOz3cF/6K5c0ijs8WuR7ueQmSOqehJwXg6vh
baYfDK/g8Sd2W+F7jQUV7fYtPP1iurhxUa6L8cUjLq8Kx1+D7DdkzSXus/Fcx/cfM0FMmBUNamvU
+VQu+SUsYpNqm7au7gnodttTRK8jcudaFJezws3OMOznqY9bgZJUx2LVLHqsk5xi44VMu63cC8EM
fDd2/B+x+Dy32X96ILf+9HMtASM9gnEXeExbdXklb2KbylV1mOhZ2EhJlnerK5wTL0+6uQWysSMT
j+2R7so/KoRGPs2+n6FmARulstP/2GgLlcx240spwIeoemwd80nWHdXcSl8AhHxH4AAYPDAEn365
Lwv7BLZ2hXZ+qV3yPAxusPgSnF3gDlMYTPhSCtuTbpHkOS9KJ9lOkFWL1MCjX15ztsDWJVpoumGu
gRNivpU1lSy5McXYR4KYOMGsUC9dyJMUzJNgZA/JJbzKIGPTNAmAqlgSL6AsmMhMidP63HHUYdON
aNrn5nvD0KkVBpPdMmqlrxnpBDUq7cj7qCptfihB6+mxJcK93ZmwQt/l+ATVN6iYs4JVZ+pQZ7SZ
82g065Jgo8AZkHWvFtZTYnvO/JlwEq0/hDXvsZY7UMBAqx0c1Pz6L5Ak6Kf0le4mSzUJS2TRbzVQ
g01V1KHJOVk8HWDAHJ+N2t+VQnOXSF2TJbckvsLOEOAeKri9EbVFotZfMQCV+59ts2V5rZAkDAAI
pc+dBEMy4XT13VA3A7b0P2v6798SVWWoKQ/n13nxoZJbEjMCBjNHwQrtkZReO/yhP1ynJjZo+neJ
/iaRaEBM2ujQ9W5M8XASG/6PFK+wPOkuj7hWrpV7mQSOBUc89wJ07gKOAr6Foug3IIZdp3OVWmrQ
qNe4s+hSYdQzJ3/Zh9jlvuBaUZu9G9Uq/jM2s4gzB2+UTXBC/JBihgW6fU1Xx1YGSabhbZ272kLz
rF01s+KAZ22ut/i3eZ0S/nhN7P01opS8xvc/+bdwqkVVxHPcHPk7xYOrBGRHx7EV+kNd+1Dlpinj
uq3vesvj8sgOdM0R0neXCtxRLBIPVfA4Tht3jvLfMIs7IAEx0CNH2sHlYwC2NI0mCPxjMIGVoL6E
ryJ/A75be1LeKsvOPJt5awCJ8zYnXKKUIVPj0n56zTQxxRBu7ZbRxR882/XWj3vRvnq+UW7EV8uo
lttJVf4BjWJ7LmkxAMMe9uEzTDdLs+GJSQqQEGBLo0yrL7vZcRUwnC9JwendMI47Ead5Z4yyudzt
K2WTkLldqcEDzR2+TrRo0wUtVwF8+W/daPS6bVyAH2qv82qJgyqv1/gc5+uNEvwodtHXkmT2YOz4
1261PGDtpHYhaKRuDqTge5NQzZS+aPYdas1Rml+hDTvk3JMcmv4pXilhb11g+NUWBF1U2cAHHphb
eNAJtyblb90oBxIlry8H2p2qSmj761Zxl712OaV05HUk54n+M3pDwyzYDogUBYyYBZIcitAUXQDy
lporRdk84aBQRczVsPBo7uBKOfuyrisfQCG981RZRWfakfaPNVszSnaumvj9nODNXOdy11/W29mm
2xzXaMdZKovJi14z//PGVO+OmfOEDNKlocT+YV8LXvDsLHfatP1gws2gTg/zVWJ4tw6WsthIzamo
jRi/w41QFNm/zJ7v+EsJthVhIW2v0Ee3P5V7V497OuVDfVomF6U0YvtqdIFY711RSFCAObsPQHyU
jxMmdK4OcqovGGKd3akRkOX72emAuMCdFZUhK+WjmNggpwTGRcg4mGBLaQe8w3l5dnLxPXHAiSZy
HuGr11L3I+V+0PgN5Inob5YeZqprRJQp8hFOEk2a8RT/93fP7TNhsBf4OQDlvB+xsP8qiUPMddMF
wqRP6XExqbUFLwbDDeajSJ1OEpRnWFjgAZMY0vrR1bKiPSe1/GzyIfQfIqr9sohlPjVs004Q5msX
L1szAti0zJafCDqj6n3d5engVviQRz9hzmnqtH0p2wi2OHI8OZvleoFyviVTmLcEzZgIsBg/JMSD
+9tmd0UE4PLbrx3wURu8GdLzIntm0tCre7wZQyuQQEtZHg7XL4VPeP5eO5pQL2ZtDBT3QbFarAJB
Du3VkG8UOnmEvvfBK5ukCcIj+ygIopwJdhpdYzU96rhud0Cq/MgcrYzrzdnj42ouxoobJU4OMr2y
sN6KdvyE5NVE/+rq04xa1xjXTEuM41h/9stlF/mJ7n0DcB/5bdyQC4sT1GSXzND17Vn65baeyhUx
cuKChe0N7lC14V5Ri3Q2cIPq/V4NmqA/fJrbpp0OAkZBxqRsNk30qRCbCg6jxpkyjNiKLHnXlhX+
YUwnClLybnT+3P3Fvw5QnPYe3PK4hAGvW9I+IBIz2jeKbGK78/L0fMjDign6pPD81CpNxFF08/OH
jOdJBwlnp8C2wC5UAiE/FbWimUHxFFjZk4QXTkZRCUovDd69MMtmjEHy11VQzkulRAuCfaOHn2v3
PoKQxGulNBVzg28o3npX/U2wrofI29pCw/lrHdiHjDLocLahOn9CPubV54DKyuwIewyBVKdBnm/W
IIwaUU0+ZVexPKpMYLhOm9vsQWQLJbfNrZ0LtndoV+9j583nf5JfH/5vnjEJ6nUzToXfK2FHb6yn
uaMhojBIRhs5+M3JTovOhJ9cd13ZoBbJIoeMkH422xTy1B+PWGEsiZBT9iaP44Kub5+26ElaNm28
KqC1JGTF85MXa0WpDfIrEuo1NIWHomSQ34Q1o3zNLRWD9Ir9qxdCrc6T0LAn9kya/SKY9s8wF9UE
Uzv/yhjwXk852379twvb0QKtgCsqeWs8PEJh3g6jfdmzGG9zH1TZQKKVr+0D5go9Ks1cMgFw+Ohb
QQxpq2rTeShdRT6mB/h/mLi50Hzm6nbpT2SCOtZ1dFrynsPV6q6ZBi3/V+zUwoUOvz/Hs10NDeiN
w7SiGJ6N6/Qvq47VFU7PP1EFRTZ0HDkAgbudfbU4wlJuuCCxsnX9jQAanse9JtGwTFEESsb7LXUC
E9ae917UucRj4Muam0nQ8MalUti3CWC12+GN7VmWEpt8d30D0GY4dpvCSV+U3G7o59/mdxK6BX4g
wrN8St9tWglwNiuNXH+jA0Ofd/lgS2ZcsU3T4riUfGmJhl6ofEevaskEQIcCLKs5fdovx1RUHA5/
w7CLaPyc6rAHHxlNaVam/tPEKbkB2IrwH4qAjuVD3uSp5Nnz9bIRhLnXP9xi5aBOe2fYIPQoZOTj
Ibo6dRnMkjiuriPf/5o6S9L7pkVfMoF6ngjuUEpuibznauw/+0QjJuVj1x74ti6L96xQAeYb/fuF
9bkwfchGlSp/uLIwwQMIsv4SduVvVslV9sehFNhWHwJ0C5fm2W+YWRtxWK++g8ECMYiC0sqeBEw2
kJ4o35Bd+fwvf7uRrCysgredwUTD6JwVd+SQFbGLB9cDL7iFdQLuXXkYVOVRdG9YGHpzPA3w+CM/
0p0DoVpQztsRzJ+zda3bsNaLf2tDDjiZvGzUGa2Q/wZ/u0QQ/FOO80o2T0ohJyrFJXZG4z2nhjyn
NjC4QAVdRmZMGDGRrLjwUXmU2svpe6hjiTNMmj0Jx0ybApz1rLB/wRGRTvCDczzOhLeIXrYN3Nb8
pCSFfEY5DLYB/vfPKOCMXSIwogYp9gYA/VaQFGKTGHz9D21NX62KoS38CKHZuAWvxccUlplhxnr8
CPN4CL013EW017U+LTQagOFoTodGPFu7SwByRFGgz5fbefH8lZ9Qru8pak+Or3voxZq7hVvCMrst
y+dUeQkrFX856QD9MDCKmXopb63dkjhJZWYjlwY6LKT8RkkArOhNfZjxdiTaohLIyyS9XPL+xW8r
4WeJ1xvu7v/DIR3qYmmCRK2W4blMO9+BbvJaT5Zhcc58blldm7NlfxCuAHZ3iQosFYs595cznBYM
YW+YaKIG3NDa88S6TOeQp0gG5E3RHeki9QjT8w39Uef7zWsCd74MK9KvDUh70AmG1oNnNT+MTYcs
+TF6Z9kGdckrDYtVq/hGobn584lSWqSDOTXihVMHw8hqxPQQYhVpl3g7+RXeWMnFyOVIHEa7tDrG
054jDr/2+UBxAfh97nZ3i6wRWZGWTBfoTG3ttUl3m2DdpJieBZ5mn5PpzRqK2ua+W6jGjIhnShyy
rp2DtTfik/ZM4ROBIZCD7pkJuXOzmSz8CWg36oFf0WDanlUnm8aywbHVpeiXE5qD8k+mWl9Nthov
/T/2BLgt7Y424jtnWsdIPnqamx/WrsO+zdrXFMjg8BjRKwcE66RfXmzMRsRwhUqRjqwowK+9N8Lw
O/OVEg9WLdY+F4IQX1/VDq2YZwi+PRth4zdGhFrbUfurTdmRrtrdMbXzTchVFBbnhPukS/FmRseT
sEFbkoN+IUAYQd/CG4VLfQCk689rdT08T00ziB1lUFhqonJw/L37m8wLr1jjtrKZkSb4UjZW3Ipe
+FQKMALB3ZWmamsxDSNAMR2SP3MeQd505NNA86dDRB/HCC4CVS8MtRlK4vkvz9wRfDzzg5Y4eyHd
zOljRmlsFaxdNIKlENqpgE5AKJuXaQ1GQ0yHX4WWBtKU4mtAdq5mk7qb2wGXnlBFroe1xq1R366Q
f+IKtSA/+dMa7zapa9lzI8fDMPGrgU0/QgfIIARkCyxp2/q2eTbdzZftJzucuyAh7TgUdJVZ/uwj
kROMVbnG/IIuOY6ZRj8/QivnqXGb5uB/fQpXMwUS5MURDA80FoKcJT6FmEoOuouFEsK8frcO9U80
mwNchNrfDWD4SA1wEE7cwAQ0/zL+pegqQuK6DXQf7r/8PAhRr/700YTBWaY64ZLH33ZPWSpnf4f3
P6XkHBIfpuas+jsPamyePMBJiT0hcOm4e16dS6tAcA6o/VeMipouXhTIemxjm+wFz38sH+XJrQzj
Mv7dnPPAywExNOOUoasXKO63q8kij8vrHnf7stWO6ypv1uxhwIqS1qIMZ+fajnlUGWiw8j0suxtX
p+P2LgD8SlxDp+3uHMZKF5lOtdJ/uUkrbeKOXGuXtjd+9Z/lNolYyvzqQjUvxmNTR328btqQEXls
rAuTE2DruflxmlFlZEoI5X0cxBXipq2fvx+2By8sYsTGLWkEXV3Isi1RCR2o4/20IDNYNdHnAvus
VcTj9P1/T0SpWLiL2uN2lCwCm1yRkQLNYHxa21XkbDzvCTssG1RuuhvHz6xBHWKebnoEeRto3kGA
d0TrOyIe4Vfr63S8SC/lrxQ1UwpIIsmTBhwG/SSR96utzWN4ZyMmTvD0l38xWeGGv2Rebz6m39Wu
fM0hqxSmthuuChwasf8ZuHGC0mRFui9/2A8Vde0tSJgJIOyv/QsCwU4Q81rfy08hcpianM3TgIoe
A572NxOG978vgGpKwJ4Yw4GU/H9wljk+pDygrg+WQgaYLJATwEEoRUhAeUREssU9+CpAdY997TG3
ZHfi818kUkMxl+oR7/6b+DQo+LTn7kKNERv1o1w0OYbkl7e/tWW7HAvqaCTNIaoDz4au2b1506Jf
cgpHuSpT2sMfCVnxPar3TP27ZlHStUCqbdAFOuAX/MlgvE+En0Vzw5K24zsO0Yr/1WtfbgBBVZV0
5H74Kuer99BkgkkL8V93kZLcSXa8iKiuFKLD5hC9aZ2e1jBJ/tDmwIea7ATQLxtB9qE3LoRR9GG4
r8f8i/ks4uP+R+JcBpxMLmBN2MLcp9hqT3VHVcB5uVgYSO/rinI1K77y8ltLcgy9ySlxb3S1G42+
XjxY7DFxvdK1clIuhtMt8Jc1uU3TX4HjcQ5pvD3xFRwEJIfPBgnnx+CH9rhAfgstbKvSM1hCaLNu
h/EVq1wZRBVhG5JGbrlmRUDiPnOcwjhJ3FHLn+Nuzc+79ekX84WertvZxZu76AsW22Ft5br5UlS/
FAjc7HjbrKyhdGsAcqyONptITgPWVeuReFnmzw4G60xaQOadFcdLnW5buWfxdKN+AhcfzP1M67wW
v+jIdz26Yc3n7jm8TWvfhrp2NiWxTprnYviSASfk1+mQ1x+3H9Zepw3siJeUQdxgaQEhZOdR6cD5
MUXqhC7MSwTiXiH6Wu8cEnjISMC4fs8BcPD+5v0x2on2kjDawxbotQKCR94u0tDIkks9KBGTF2tw
jIwWxnMnoVFQ10xSecEd1W2E68AzKAlZH3EbQvgHUICFlRqzUVSwpbazaXzQYwNVL0NnockaDEpn
RO7dvRG4fDBUnmbmUIj5PmYQI9ZVItEp2Ksjz0E0siic0X5nKgsRgVgxHqpM9wfyMP0J+3Eze1wP
teGH0lI62p1/j1yKer/YIPs23OAm9F55BnOyZ7MkJsQ/wF6cV4m8NSSvvEDyT+KlpDpNJ+hHk3aD
mgP3jUrAW+B6iFWVdKLOrX8pAmwRhxRvwKnHR+rpJ7TYFkXur5MHirl8qQoHfbo94S/cII2FC1Su
RxY35FgITgTlhBOgIptMLLfIYdCET4IK9fIqllVPOO7PtZuD+djLSavrHfYqOI3ZGYegtAv8lbLe
ZZPAXX4wN9p1laSa2mr1MDP4cQ3IIUKsSWJztkNjWUBhGVM/nmauKysfe73fQsje4O86O+/wDo5M
dHlHJBPWGW08GIsKoW55pp5AT+K9T2XOkxPWWRhv8ss9ufxdN/6X78x1uHB07BgCh7Qc2pydCrNB
q9ywIilrzhQxFftVL7dktIRy2X1vmTTsFyBpRgyKIxb+WJZA+ew39wEdUFsBf2b1Z41GPejBV/ss
ZoJSEWTeZVgAC0yUCZohHLRG1+ogpkRF4LY6zrUzszQaLN5L2xJbpU46/z1r3Oh4/ADC7tJY7xch
v5Is6n0RHbcVqRgJ9d2gWLkCqbOo17nL5EwV2ddONJlWpY4j7XjQsXu2IyJu8PFjFjeLOXdBMrMJ
IXee9tCbrLnA50xQ+oQW2nln9KjqPCa9KSU2f/hjtuz104QbWkHjWebPCxSZOlnl6uooszJ/sZ2f
rIkXV5u2sI2H4mI9GgQrK5IHncjtHdSOULH9zEEvv4dBqB05Y9pi7czPNO4CsiXt0DhIpKQcBDUa
7X8YT4yU7NvvW1h/+8HR+5sPeetUQ8iS3eATNXhd9dcAP0XrnLS+dtlzYP2nGqnjuSW4JwNgaTxv
MkZYRhpuK9u0ilexZAq6PW89LcczcCmuHgCQqhkV6ocSh0mp06NeGQ2KAeasRTGhXDhswaXigt90
npKXS9ufa9df6lf50ZPV9nVPmSpM58wQ2Axx/4Zk5DQx89eLnM2NVHDF5o7nrY9hWWifvvtKUNEg
TSDHfW7tx8FsrEDvbhuVRMt6xEfcTfGOJowsZiJcA8jYQR0ZZgWDVFFudwa3ybVUvnYNen/LHcAA
VA2q0RqR/3A7nC662+Am37oxmjTD5t83SvzEY5CjxifTlhKV8FrNKTfetA3psVNLhDt7LjWnJC7g
odu6ooMXDDYpcAP1Bk1zQGjw0a7QZZr3VMent+hqkcrehrcuDXIjgc2kpLrQZwYoE+rK7En9ilpa
9OBj1ed5d2JDT7SaPb2dG3K0KEMlC0sc0JVzhZI4E64bx6JluyOSUORO/rqS92Y7EjsdtkBLbZlo
mZS/vycDzm9LCKWOSlxgHgmGOLo202WeuFdYJn+qNI/JK392DfrxPPFPFDWLUPIAkHbfB9N1Udok
wfybiu6x2QZX51Ax1JZtL4bHvgA7O0ZpI0QAL8TmzzUSsBWUIR1XS8dLrknqbUZrOCZHH53QIbMX
eyUNrh6cdr3UZSIkVdEhkXuCg0N1AoUJUVF2e/zrPTIp7DhsPo460/QDe1Ed1yz/S2Bm42Ftkmx/
0jo89ZAPCOKDOvghGCeKk8rLLHJ10BzYFylMFMUQjSO7nrqIotrAcQvLQH5Taxn0BpVuEWw7eUd+
ByacZw0zuRMsttxDQnGQiFbr4q4+LG5m1znAfc0xVbJ07kzsVj2VFBmWOJSeLTWHRbmpxDrifBIC
OwsSXRNOsVtYL/p7aJF/lrcLc0CWEezfGayOb9rzDWoncCy5LjVh/unOFigyy+xYedXJcuFU8ZQS
uB2ksE1QVUvxePaGeJtA88zjwQy5tSq1EdYv0iMNrs80r2/ZFv9iIFITPRFkLR5iTAQYJ4fzXOo7
ukDhG3huwZ3og5q8TLY64E8v2Hodt4Dy01aWxjQDgV+wlVulyNnSQpsekjMLFn4M3d46xprqicqQ
0nPHZh5E4AOsJXJB4OFylZcAnxBMj/BuofixhzyEhRWrOGj6uVHeQlI2R8VUL0Z7WopbcN55wlRN
WDLCWWOTRKZXuw6mrlIuuDTU1TwLz1GUlNzqD9HHMaxeWbKJ+GYrKfI0BNwfLeRptW9pwRtw2bHi
EnABEVvzKp+hTfXiezfeqdCnOirKKKVeEOlAO8CraWeDb+xgO3xEYtXv0N7w5wS0QLB09f1YpUup
c4WrhC6BIyatk0/oJQoztzLJb8vxTJZo/zRqLxWrEG+hjbIOnZzfX4+uqsdvZbJTtWlkvaD5Uoml
IrPavI7a9UTuPfv7VptLwHWht+Sw5aZgQOEVKn1yXVd1h5AQhHPxVgpP+TJ7Hyg1wMFS4lvM6LQL
MvTRslwZvX838OVAP8yWXFgmlKw8XP6JzPh2uqWEc4s1AZW2PT3tRf5TzfLsZN9nNi9QF8jC3FA/
yIAZKk6maajXRSSOiVqQ/Q/2vfKU7tRBsGMk1eMht8+S5iiasoudal8HR3S1hV0viXpiVamI6dme
vD59SQqt2kp2pLuNjCsC7xgnNm3iwgZYpSuNxqqFUGOZ+pjWbb6Ym9tYh+0ePY5LWTDLBEuBxJo1
0U/DREw1aAgFcJj78EcXdxfmfv9cLl4NhCHDs6u2J6xGk+C55wiXlBr6dGjsRLuJtvxKO7cPH95/
GCPocUqMeqJmePQBxc2yWiDb13mS9tEZM5d6uazQFCO7MzD/NMPZ7qQmcb9djKGh/5Vx2NUqPClD
EjgzFSlJ2zMIClouQY9UOU2c+9stW2i9plQZ09v14nitoaC9IVVFx2DBHWWpplN5GaknEQWxYSwE
CTozhXHk1oEMOs7/c1m8HiaJUn90cV1ao1zoV1knyKQZSTvshDl6EhV/Hwcc51QWFbyoEpc0IBJp
OdQXceAPiAK2nfS9LGDMmfXpNA7Wo4Z67IVuVXuYAQGtzv//bTu+erUu3WBXmW/t+p1sAUfl/1fU
ZctDO99Aq5y86PLYEqTSZ45hvzQ54C/1r+/ocQEfk2nM7Vc1JuZ+cQfoLTcUHCyi4B2HoIJgBzTD
P+qH/ITAm6JErQOqNRK1Ig6OSuw+f3bawnJHSNt5MEiUkEoTeFX6RwKckpkWHS0kgO7YMeOvqBXP
fIZfecypE/c5AdJIi6u2ytI5554PZBAmsLPxOA6DwX2jnNBSSDqY+Cje/BmLJ1pDkLsNVDDKriVe
uSRYYECBfGmtTnxJSuocJpTF6HUGYSpqxMsA7nzIYDIb9X/idzQc1GKaOSJsEgEobysTvCQM/ZoN
wE22kvDvogwNrnKPIQpRC9zRqjawfe0XXP5DIcaDOyAgId8/CM45H2V1p8EFhLrif0XIe/hwQ6OW
TLjiPyHHyARiRbyLxTkzaan95hV3UEhtdVZEQUsgiCjH9guwGoIzTFjUkyEsxztup/FLjxYNBIZM
pI1DZ9dnUsbNpOteostOOVhAJufbp3RjecOGB1Cns34y27G+cT0jNSwttJS0NcIA4DPccUxS2Xgf
brwk+DqxLskxvUAprEdOWzsldT2gMnGS8pRHtaVqDJvjrcHlyKYamA1QFtnbpHQVKnmcVBkJX33j
Qi0Eho/hlyDcojbrMINifNEnjIAsqMQZtLlXSu3wbCsV7Gi+dreqt4HKo/JxF92G/KUUB7Ufc7A0
CXZuh843umUKFii08KZJPapFUZljDv3XkASp0Mxp9ooE/0BqYoReYOXIE+jFiJBWdD33e5KoZdeo
sHwDmteeckLecqSx6MF6n6pYUX6bGddCzUJMB/WVKJKlt0sxQg8G2Z1VE+J/CcMBLlbJqPD2qF/b
olshjcDDh9tul9O/t7NWFUFJCWKsW0Pi/SwAx4f3Q4slNXGj0qXi9VWzIy/ohlsafdCFU5DYmKe/
rZAMicJYSoBHhbXqE99YNnP7tT3PHQjDQ8mCe5FayZtqPpRt0SCHPBSu7acUCwQOV+sxWPevJ636
89zLEEzs3AvwAn4jHHj50CRBRejfs1VDQU67vw95Td5Yxpz0zQfHdWRQWIrssRO+QKAmNMfeC3uE
VhqrnkXsXvUjGrI1YpgmbVUCG4FRa7JktwIWDRBeoq4dRVq5xFldHbPZSNaqW1dwaDqJx8deMKZW
+TGkecXn+ftjw6ePNua9M92mEcyM4DRInKc0Plryk22/vc2AoeTqlUkQWJib4SKFTAaiwQf5AQ4U
0ewkkbyIoAqD8K0dKxb+1XS2ZtI74otlPULXf5I+heRrC26+YlN38UueMXtN5tlM4boot4/A0nyx
B02CwwVQ0HIcOui/q8JmIOiDZnCPc1OaDj+aGY+/Ub0alNZdgKLdwgKa7JfVW0VqInvokCQW5xzv
ntgBItgm+Q63UIdBBW2J915cNmiNRoYU/iF2YOcI0QyERrdR3fB/0cVi2k7CejuObiNLIhqcRAD4
EQfl4gxfD3YMBygXX7SkEG4pR48zj/73FJD4tF6YH3a7B3sBUtXJ9UkP4mB2i06N7SIV/5ccRE2z
yZIcHvreaEJDipuA+Qf/Q7NagrWEaYQrZVZNugkKy2Ex+gyEmnD3zqdLCIc1z/3iHpDAo/RWbuQ1
OmDve5Q/ZEdIO246VVWWkcD6bdSQxxNN8MpIZRwrdzb7W8w/isSPOKO+ydLKfhtaHTBK75zchah/
/eeWUcDa6ywpNfRnLEsQp+eY3KhmK+cSK9IS3MMzKP8HNyjzkVrdt7tmiyfGjGJGqtVUFzCoIOCj
v9o13cG4I6yNasLCBku9fHHjSCWqWLlWr02dZwLVKmvKYg2m03bfonAkYDl5SFWdR9K7HAy5cKDH
11F2EJh/BCFS7MHA3dcx5W0m7MNtebkQfTen7q/efQRTVsm3u3as2Y6uz6kysphjcbnwfpDZWPuz
wmPZCrFPX+/p7dC88beVQs5Mel9FcjDVPjwTqtyYTl81AqX/sGC5R908h55B/lBXdDFzEc0rkEry
2Ot9vDBctX6azx0e+XGikHUkFZBv3C30ERAlwyBBH2DyH7C5fCCbIha2OoQMcgo0VIBs3PqLIbSZ
pfv8GrfTbn5PEy29+0bppgzzQZa2JEpf71qJVtp/bDPDYDZ/CvhsQczW1mCkdHbFdljfm8HpMyPs
WsCOh8JgEUBY0peBDcrNUE2MuHUCaUtHXTTN/iR1T/fJzie+WOnTntxmkI2+uKnKEMuDVHqnwjrP
9Jbtc3cFaMWFfFP0bt924sh+/S/lxRF+MpVkC36jwT10e+DZVUwg/390Pmy2dhWwqJ+cQqLxVX52
9FrhO8kkH9B/QabjwNe6k3P+lWb5J0vuJFKoV/x+GyB0HivbfI2vaiphUCLeFy4JDf/h9XUJETZR
V+DIT4bBY+/gRinDr7kQhCdrqZvder0Uv7u3eEzT5T467ubEpHxmtAogR908n7kyVvS8pjSvXfFp
Ev5i3TkhUvRiH/ICNNL7mvgA2FQ5KA3SHBFJdQwysL2KA6aB1U7OaiqB4JZ1y1CYvf4U4/sRcXf8
JelmwcLcUM7wOiS0NRBGBhYrISuaQdPBYsRfPYIzkxXq/h2plQzvEPjp9H8Ws9MXta+siOhlerov
hVQDiQSVyd9MLROVCG2dTl7c8Jh7STr6hWeUvVrT1FWJogEd5Vk3SW9W+53mgerWvzkDLY+QZ9Fj
PKCoB1UOQnTWl+/Ua/bE8W7JajovqVW74SpVfQQcPt0UJ6evIPvhxJZ/JfflxwzCSwn9UQZhCp0j
Vmn9mlC4TACb3XYwzubaiGNTEVZA9PoKDHSZGXYGBn4zETmcIIS8vk+jY2TT9d1umTzvk3w2qW8i
sznUm/vNhcckd9aNKcp47WTA6nMXxKBSz9kRU9YaSiR2h+lh3rqq4DD7iuHCkWVv44sKz/2J5tOd
SoK5/LgpVt5Kjp2L/y4BPedag8TAYTDWjg6Ty+vAU70LDxx6gomEhjT7dOGjXNr7IdPpa8EzcXAl
kdmHmKUcPxSfajTEfB9TEBgvCPhupk6C/oFLcbMnyEHGBODV34OFsvxkOu8c1sGLFqHqCroM810f
SgBwYc1SGVN/qP2fLWNfmt4U5LmDIU4IDrwdmHW0YoD4Qv6fQWciLG9TtwO0onzGe87i3agTnRP4
8G2zO+UZhqWVvawiEJQBMFUi7hic0M/l7VeDLUxveOpFJoFhwjMP8RuIsBs3JDSUIdPg2tTaBCz2
iRWxlpxsPVF8esF9WC688InbMirdWl3Tmr5lPgfsd04bWaUSZa+dKE9V700SkVzDqUZrT6ZS1yzS
bHt6BVDn61l05EYl+8uQCnaYzdd5eFXjmaDCQEJI2VCv6utRfRhCg0CjYS/iCHgwpLJffkhkw8qz
zvXyEqCtL9PseMsWB3TbVTTukgWeB6IVxSKoxi/STDjHvP2wBhHv2qPwyROtxFRfrgTi9277UD5A
EomsFurmPm0/b5XGjlN8YykPM3/opAJTCwESSxIjRly5L6G0cts/F/usqeg6PSc/FUSwqnlQSOFc
P/Kvqmixzec6h3h6j5J9lL9TdXuUB2CXfOmJqOUo/f8vUgOWZBASY+wDNE0AQwyz8LjZETYTnK42
65lQtNqxTbA8iSVLQa6bLwJVdC8hyfQFSzs8tm3YwWs0g9nPLvTwbILjWiuGkIVaDAPRFzvrEa4+
k1D0Gj+QYGSRkpj7nK5bnbJNZFtQlO2JGUCnE/Bou6vTt8FOSGy2b/Y2mf7s9MQ7Gq3P8WRT1cLh
9lZzBULEapQQqw7Ezt2XRMEtZgEDDMHTbtxlgKtWDOysloy4G2tKPBrVFLZZfur/T9guhqHDcI3q
Y4RPvKFPf7N4ilO4uqz7jLEsjANDjNx5ijdXB8JOnCeMieoqh+Y2qp0nksB5mnc8ls8ULxfPyN76
PY3hWvVvq381BXxFAy2MIOzoUQ+/GrlCtlMwgPWGucWc2n9y0NIryipoiRIjIP4BVQpLcecJGmhg
mYYWv8uhpjiuFZ5e0W4jl+VrYZGGJY3Y5x8yFmPcmAokrNpsdOVOqzKZc9gbdEklbkuvTsxFqrg6
vPTO5nZ1jfOLRiXxOJlWcqVbZMx0t+L9+W/5FEv/mGJ3gXOFqHop+pjmKA86p/dGH7vQzmGGf+o9
Utd8xi6eEyLNuuVJ/2cjSigqYDPFR2E+qfncLx6jd8C4wDqffqKQr+whMXWYqrVWwRMEvVTNtsYt
7DkIPvtCt4pNANTQjzS+zJwupZgWeNoHci4t2qTOi2md10vHNOASyTFF5u568oZW9aA5GMbtbPSj
F3ZOF6sxPoO2b2Kb1puRN1F6OGhxvmXUSJtXEcG+/5hxPgcVXWKs/eQ/8oRCSLengyRkUOXelRyM
wfduE4yXYvDqsGD5TUPZf3TaWWP9nIDeJMnIOC4RLDe3XFFEMs8rEh8h5i6SEdLair997ZAEMnH/
LdUhHOZaFiw+dtHawYdCOe0wY/MhDxtC7+zuN1ArcxJAfFxQdZeOXwnLd75Jl4jD8jJKDwuwde+Y
DDFijwcgrWtPrtJBdJZvumyU+knBTXgTSBoTciaPnVPfXDpXhERtM+L6reWgjR6Y90eXlhnkId0H
IZUJIHBvbJesOu5r4csG56v9Zk+AprkfkG4agSvKlbJmy0aP+N3gkDyUzsuOg93uDL8OKmVN+uve
hDH/VX2xSPexmZ606n1Cf4Ku4i2m7SjS+YO4XKSF2W8aoXn3++FtSJ8g522+62fmLbLCpTO8uB0l
Lwc3XjxYhioUHGi9EC3mOjtIP/XDh7rLzhNToI8OLn6rA7IxZbTt2cfORfh5T6KC356GB6y6ma4H
xnrWpiSwcDdbML1N3CRj+N3piX2RaUlLo0hJo6cEXN34XiX4TEvrtwhtlsl+t66HFeziy3pckB8c
3YVNRv4NYh+rQtj0Lua4CjJR75KuCIvPGKZ/3nXI3NUU0Fu4DTNgpKXJqfRIToBQijozCtNzXFL5
g+LWRGfomnu2enRFOgAvR5JHFEC39xdExjM/TeTrB8uO4rC2cw6rKr7qn+1gM5jAmbGQBEOEUThp
Rvgiy+0FWA15HpTPpEGrUyufV6errwpMlSigCaIPrlbb7XgjCzN5SYSxpKwYGkJOFcPf8zS2YYzA
hezn75uG3Xjf0Tqq0sV+cTJ7NNq9Ov9L02fFvoe+rQG2yVFfFOjG1xmg61lqghQh01aMWUEeAdfh
4u4515ZarK+d6WMclhlV8eiNNIUT9ksuGPKY4v9NKapdGJv97lcK/Osg7oxT0WZs8L4UoiGQHATC
M/9BFGjnIyQMzOE3Pp1jatKw2ObqxIf53+n4QIobiJbjL2HI+4hOePG5pB2C1QJ9T+pzwUwdsb6A
exLFwfQD7o5gM5ZrMcDSrYfn5cgDdJjuEKGhSaNIzKDn3ewjaHkB5s3SUFU8hiqOOsjTn/Q3pOsG
LDEpO40nvSuuhmJLe3E6vMCJ02wKZOT287Gj98vWgP4hVrqeaLDVI+PtpbXjQ7AmOItp6mtFl5bi
mSBtUazAgwSTa485yAzvC6RfP8ZToB1ntqnqxY4uBWSYGSp9YauzHzphTvHYdrLjrrEKFxnLQZXC
fi+1xly1DBmZIByPpAqrAyGvWwxw1tipULlQcpX1+B5gs3vfdRkPtSrTKuwwZhcLBAD9mBE8PQmS
3NtuLRx3KJC1gls3fzS3PwogYleeJ2zmKtEM7YtqtF+KWFWvmVpu+i7QruZ1W1HjT14pMvv/WHAA
FcsdXNE2VFnydAXPO3/c8dD3oJsCzQ6u9Ron+5F2y/WAWK88WxZCG5cNGBLdpEQnamhYsltWXI1C
dXS/rGul2NEBPAPSY5Ozj3osQpyZa/DPhYsWE2qJo2pexeMR5OxcsArmxDQaEAOIJoAK4TZMazRJ
5Ap0rYmtiN1LlYQCsrvp88NDB5p2PCwJfx0uOH1pSdbCaqBJIuktf+2G5IvZXpDzG57PvKEI0wJe
qtSVvFqyTbl3eoQBWzN3TNxvmYt1P8NupMr3xAoElSIJ0HgXoQzNMSRw5qYzMIZ7hmEM3WuIyEvG
a6zUNMvDqoM7Wpsq5eIEVHphSRrm9urH9qALGamieUeboYtZHPrDmRuDQP9p58qFOTHXHH/M2SOx
FftfGMnktV3ZTYGDdis+Uzq7VOI3Jcw3cg4oo+zew87zgjbO7QcPoFIP05A2JNRoIUuG8wwzl2+3
ER7vQ2JDivzXuEKEHn0zfG0F3wLAtV03QiqedLIkxdGdlj3Vftys0iG3pUm9x27NkWvT7ILlCa8B
QtS2vBo90dLn810tSXRs+tnJn6/jdhXuIiWxWBZvfKa8T55AyZ4llJAILznq/omMFZ0tNIIkTjr8
wIwjJGudqwfRNrp34SIuxT/fVjFh0I9rAESz4sxmiTPwxRc+Ew/aVDwEFLquna3ryzu56ko0DFM+
uMwGWyxIZUlCQYQ43pfgRZ4tmGsNP73a3O1yFZW7D9Ctt2QMZSsqj+xF09SMqPmTxXTZztTzF/Gf
lvt7UHs+Lq545bB4lkQXNrx2Otb6djID30ql1j1STfI3BZDPFjkJP6Wo6+yTW7coLvUsyhV2Dzg9
X5fGogY30kbSCeeif3sK1hZjuDpYTQWrjmL1hUxFEebhTWoVxjow/M/G8RbBwNRQBbcEcxIJDWk9
0C2WkOBO2JEU0xoWFuLT8JReYGQLM9TaR6xF8dbs2nV4tcStkCT7Otw3aRMGeaVSvxZwIvCINEsG
kGysV5f4pGZYUXUA08Sw58BaF4wblTaS1jLn4eiMw8B0g0pTpQ1axUBPT+qGAEkKgpKZSmRycIfp
gaGMhQ8aMZR4hag3NcAHWFPUYO2AtuxCD1scgo9ii0R8v+EZz6hoZG8jvM0YYne1iv4yZPXBpdmu
ueceILq0Gu0ztl+txMCnANYzyvz2qDWwyTb16pnRJfI7me7235+FzIwfwTuqBnTkqcU7FsH6kirD
9mn7zx2jFC5mZ5gPjLtPszo5mEETd+gXvYKpTSBJPyrnWExHjzYik+ir/xyEAJeNUGTqiG/BngL1
1Dy4Fecjm+iZBCYYAZji+P8qQ7Mp4ReQn1PWoaZ0mhfQTKb5DOERdXklSp9xPYGaaaYjIPhNw22s
KkA7p91O200rsRqeEm4kOawBCMKihZxZe62z6YfGVhWbf0AD0oVzT9JutjwE6FEIQ/k0h9+BS/Dk
PboPUZyXfyaSn2E2V9798gfFc+jHBbN9Pc9Lsi09k+PCJfWLG089PfjtFWijHyqZIJfkBCa2VQ7O
LDaLmMo+dm4DZ2enR1t66aRoWuWNueA3v/Og/gSVwv5kXsUFblvx0OXKfpRfPR9LBIIgzSdfipaG
2Afgry4IBidSMRtROFS6V6tnpgRIFppcRMO7kADosID2XAGL/qKnJNKdeWYX0cpeB4wB21+2nPNr
P+H0i44KXMAeCLeRe+s9nEDH0b2JJAOYSwT+LTHsQxL5BKeIh9BXp/YWlOUY1A42MecsSwabLSHe
aelBP0njHDAwA9lIdDTns79GPa62h+m+60WvVPowYQBXTLvlhanWh7oOeFkz+OKnjxzkBNKXkSlm
BxJjG6va94CPrAg1Iiub35tZtyPNliaJhaNukH59qMS+rkjylpfgwzupVp5LU492fFO9AsW9QZCv
QDPzdCqQe07UVU20hz2/IFKNfGy3+rmatotJ3vPtXTFj8REkwkcQeFo2EKkyxKrZTFTbTx0nfzEj
UFRCJ9TecndprrkszZB4qqYJmpoJXxgToFllsbXzVRbaT7Ddek0Zh8COpA5xHpeG/deZMMATD84a
oXrJ2Gc8a/3iocZ9wC+ctLt9QpsFmbd8c7kiyKuxrryBY8icy57a3xf9nJdBIvglF84awGmkAcyL
LvAIs6KzeUkfQ8GQF7XHitW2dnco00H7BqYbz3sgCSGHzNZkdsBWL24pzht5A73gjIhiMJTAQpZ3
f5M6EiQ/GKGBdRpL1+bqMEee6b8zRRiGzV72RvBk8FimpoRrZa1/DlclM0Rdn4U7HVGN4/Vjnney
SgUrtrL7fM6SjTSs8Rmf9uELTbvvcqNWzvlJsizyrxC4VJbxEEG1/jqDUvrbpwu9GbBK43utnt0c
d1PyOBLVuokh2tl8wvT2AXvVhJbaFl2pZFWO3YR8Dv+AGDze4F4z/GUyuQ8bmL8hPh1tr2zikAS5
lGcNemISBb96Kkt4rK+bqJe2jHHs1FOLhbzjFPcOTfOtkmwsyUj3AK4mmQ86QTSdgOUQC1oyOOq+
H4YZ6QFHU/to9JzCuP+DlPDliNMQ4dGELAlGo3rSkN3R9UF2RgtY0Fd2b18yjpIodLQCCN0S0Zmx
eurers84o1X/Zu4y5goc5cFfOcLlDiIgNzUkz5KxSpi+PKoYMavTubnAwhhTpLfL6AHpq56j8U49
gaDgxw5QkY6Utok7a3z5P+rsZ+0RJa8RJYHv51qwiOYB+XIJ+dHTNzfUej8+n2G2rvQ5NlOZbAGc
y4z8U6evVMKxIrQVzP/IWKbdmXX4J1IzE4GtlcXPf99V+t9HcnlPVVtJzv1WYds+vF/roMqdEqYq
imJL8cNCTSCQxZr/i9oimbsofHroUbHi8/+wlP0k5FnJDFGibSB41STJ4cg5jkD0U6Nm7vNFdVRy
6owY2qcaCYBnT9kq/YtxFShajCmZuLwfubCH6TaVCH773T+2Csqvx+BmzeJNhY86ZTO482bvpS8f
4TPRgF+yTMOoMPvB6GXNj+Zpb7Sqsn9lyB++tm/TsSwjpFQiU8bm3s1A/neny8YYP8kx+zGIh8Bv
ApsKpJeWon1PStml2LE/TQaRY3ufEg2pTZGjfhgkWK5GP8ahOjyeVftcSGgBtYnlKVKyM405yiBb
QmzyWu8lS7ab51GJmN2f2mqOfyfH1NNZrbvGm6E6Qk36nSp0rHfGGCngLZHUjXxnnSSiF5ofe8vN
4Y7VzbAU1Zsk1O7PSV0zA++YAj2ILfU9LHyyJxMnKrwVjYcf2aN1jcsRHbEYtphnrZFFvd8XIBZt
y1Ed1CYDRm/WoEQXASa6RPjvaHK/PkMCZ+TT/K7cd7m9vLGt6bqhwbRXr0s6x8DlR6zLjLuxfCvW
75f1MPZYa0T1AB7L2oAO57MjeK30CE+yPUFZmHt1ARVvF0zPISiGBkg6gxtmThEZS2T/W1SADEsA
K4PI+23pPwZrLWVgYu6OqvHDUFgSQg5aId3qEKb8isG62rtOsoX+X87uiw27fV/kTnpym7R03pPI
0J8gs7UtPH5Rk56Pl0MtwhG2x8RC1I7bl23LNDpsNDA0g1j/vuJb7B7WdCoAfgg61AWUZtwbOyT0
ka5Wr4qI3dMJE86U/w4n+IhckZoeP3Oea9CjM5beu23e3k/of4pZaBSPTqxLxAs5n2cHaH6tvfKy
ksCU86mS7zU53tbaLqGosGx+BeMJ2JcbCOCDXPXt0zYtjDkwHzU3ikwm190rTDaQYhcz/F6x2R4z
lWR4Y+enkPjw59W5zeGf1/y5dBuYeSqrVgSnujvm1wcKLQCR7nImTTllUgrdbBANq4X76td/HM6d
8RhCAcTri7QWQ1IgDOfuGW0amvdoxDqzA0cjaQpnLk4GB2b4dKLpaoa67JgjIIaRKhPFpDY3Qjqu
ab7/5njSishuyZHvYazGFBS46Bmv+KApwlvD/Ssv8cLYIThVlAWuXTC5xtq6cryh5MAMdE+uDy4o
PHPLJf2a4sjjNNdKb3cISnb+JBvKBJXPvvka8x2QA0wpw4fnKNcN3NYmpyhK6TNdUNr5UAQUT3M6
ph7nHqmmQPxKNVbeNJiGSmf3joi3yLupWJjEoAGl4tMf5G1gDwLhRX0yRRxY5p9ACaWslSlll32E
txLttfkntuhNdG81B5EcIgxCda1z8OQTt16/LMv8v0ZOezobzK1a08dvXxpISvZjYljZm7v8ZNKS
1iUtyKE+T3ki4wxiIsy0V8EXZWoE8E34Qo/gBgkGY9ZNzOJUcMHntCMG6YNqWh8Oq7Ub7xtSW3DN
H3AwMZHE2JI70K2frjqp/5uZn4ohjEj2ZNYOoZ6U6Hsd9Nr/AbZF7rK6t8tCenPxhqs/yd2PS+6+
xj/aAT2FN698GoF7EWegglOnZL7GqcU+VZqeu4GvfsP50sk9bsIgIiA4VIJu3pY+FxeX94/dRyfR
atE6uk9N9m4S8yYMosJP05aIFw9mFKtLYkkpaxERcGH/grzsv60MA+eBElQY6+fmSClaG9IMXciv
iTAtyNFJPcaW6uDYwuLi0uh+9/hwCUgmlz9mcrtOt9+jRMiepm1Abd2rDEEUt7BY2AcWlIV4ht7w
s+eM+G5i85Tp/8nFAZctQIYee+6xblToO+gWI4Ug8+HyVW2xlRoGjevuokTXqUtA9MfDb71v+K/D
bt7sfZts1mSa0t93DQ04VwAhWSsAiUSB9vqEXk4Ma1xS0P+GD59fF936N9SKuBW8jnGbZSSely1M
PPrQpx6P7UxaNhsZ1LNm8leIhv8i0Lltu8LL6PSQ3eeBgk+PSLvYI1LQLBG1gbT63a6Vry8hXT/q
YBmqcXceAc2C4/4vsbJaqHQjqg/g82dO86CNv9FChRUh3CdTmbekCFpDxE3yC9rCrw9sp9YsqOUr
qR9rD9jq0Aqo4/stluC4jiPwvt3WLAmMT3/G71lWc3mf7HdxueUoSfmr8gAG7RUwHd8GdvkwSp/s
ZJxrmGda6edUfhXBT6QDXGoloX68DcJLHjOrUfpzFLF6R5Q3ErlMZSTK3kwbZvT84XHY0UYRnGGD
VH564Xnf7ovWa9hIu7bdA9sNBPnk5FPhaDGAvHEnirOl4swiCAimdwyT7nDzdYB3FQnMyu/R6sq5
9jlLCSkVD3jRb9Zr3wUkskQ/tPHorcfmSTTZyEiH95jo9tF8dvM58dSA14+l9NKefN3SgrESUukz
KZRIkY7zSGkpi5befY3aPD9uGntWDcFDuyYDgY9OrZLt2Of/ZtgBUGjJMc5ibsLX+5sMqqppLYVe
QTHVd4hxfblDdscFoz9V6HHirVlmOQGcWn8ORKt86LwePKeDtxGW/Yld9UW3XhWH+iHTVhmtY2Tl
ml2C5ekBE7mwTmRYZ/yYeLORZgCSUVFS9jmDQCECddzvDSf45eruixd4PlRIq/mDIr2Yo0LyXDIC
XxVmueNRD/6L5op/YpUA/EOJ6aMA57wq0SUPjU+NHVCLU1boiZ/eH/23DL4PBqzeeP0wHGtQplgi
na541TgKsQVs79ohLvGH1kY14ouAYOeVNkPCuPKwigGXjw1qW7TCheNvfK9I4JrIf0pgcSJDXVOF
smDsoQoT4ypEwlQYS+dtMuvjjiY/wL3n8S4cOqU71Bwl1K+TL7d4QXW7MxV4IZaTnFjTf0pp47LS
OHQ0t+DyYjQUjpGU7sl3xG6Xu3wfF5zDaLkFQfIXx1oDad2RdkYQCVy+H7GNeQp8Fz0Hn7AfpKWb
GUL8YCXgNwbY+EGUwB28U88VFgDjzs1CKj3TUMD48uOktMpfyF4On/UVnzjY00943YuqeXhvy1OG
z1qqRHtsA9R4IfKRP7f2QaCTsy3uXVjdjg/R4RIvZWorncwlxEUtZV83k/7/MUZBrN+U3Zah88Sb
qkhBYDiRrDxRPLi6iSvckP4Nqcz3yiCkg434tHY7PsjkT7zC5OEIxLzxwivuK7X2XEpEmIfY31z7
WzHTAC0Ik1v9d8geoAk1pHtMgCFBn/bkG6q7iuZBeoVFq8WmnGIZMOUYKO65QwwcpyMrVKmDo5cK
6i9YHjzzSEMSt11hPn+Uo1iTnDRli1nbLYXuV/08HSakU78XLyzY9SscEiRpQC7XcgnyAtofJsY1
xw94R1ncSuIr6EWNKwKojC5Fs6zEPwG7WXHxlBdZ4mxqyejkW2/OqEIzUuTT9khTnZwAChxQFl6r
ZYBtvWDhP1Z8lhaoAocYsmFm3e5Ge8EzTZRxwy0DVVZdSOkkfnAx/VNAyADtniMXo8fOdmsElF6u
AOJM3XvkDh+MGowDyuThH42fdXctVT8LA+1Y7wxkJCEruzAJ6g9UUVjMF2Hro4+8fuvRgEUpoFAb
JCRM7OZtKubriArB4PSwo8wO9WwCM5DGd1XfK3Qlu8MnOPKfgA2lGz2dte64FuqVeMMpGbq9xuo2
IQBA2U2rMk8Qzjj5vOS4TC6NsH7gKv0F0vTgvH4ml6jKfazn7DeYOFpVpoK7OS3Bl+srnXoTzpZM
L/MbOcJuxMrgpMhPPcIbbn+jx2VEXqT5QOQl/0dPU4U4Zj3rNtu/AGhMePnbXVhx/NaDzsDWRk4C
KKGBNbCQu/hi4FgKpEAAbL29MHX/qL3Ut0NnQZLwXno/pEv5dSp8TCsy7W3Svwt6ei4oj2vUGLue
nN/5+v5S4zJU69SkgPUq+qI+A/oWPyIvGKmPA+nVNcJmQNRkRNsYZ/CMklPGWisUG0vECsOxNWnL
UkDHCQIEZwR4AtSiu3i0nfu5mJnljIeBJezebuw6Ubpg9PSlQZC3Ud2yHrmMDxdf2LYL5lEa6EX0
9CFQKC25bXl/hJODdZN5z4Yg5D/qPBdtbvNeARoUAGW5/ulsyxsxlgOZMDULeLm0FCyCpVeXJK9Z
Kc+IeYSdwc3M0J93gvPxK8BG2P3OMRaEQbesbtEi2yPkvmjWZnqASOMekFaai8uCm8eU6YAt7TN+
k9q4U08M117jBTIo9tlbOmxq3XZiQ1HUCYOQ4mnNXkWbRp/Sr91peIGC7KOYKlbicyUEVf9u8Q20
nVrLCkD8pGUHBNF3bsYXI59LFH8W/Abhd0PVcnv73NXFurxEcBDeafulVltQND1+LjF05pu8D6iZ
Q9ely/Pp+nsZ/1UsWEAyCk4ORXSEl5/nEBG0n8Adi4t9omjvhTd76DwVXhp6wFJljoTWVp33EULP
uuKCyVFonkbyy89xlY2v/vES9F2FBSvb9MpkRNqPaeR4hUKPLJSK7zhoS28DJnu4OduKmDs7fpQL
tVl14MV3Vd3q7YIB3mHPgAwu+g4/foi0slmBsMdfdZ13FFoJnUnC/gla9vogEecfKRFhSdh5xPPs
TF0rqshy2Pp9BwrFByqIVrFFzw6/vnJ6xXgvAsBI+wdw1Q99opwV0L5jPK+A/Qdhn6acIY46htaf
n4KPbddT7+Rh7yNXOWcWXreCb0vMuzJPVp7VQNyAMwnvXyp+lj3qwZPoeDNu+4BXiHyUtoA9MJ3l
NmrfR2Kal7tNjWd6ShV7flylBrEeA2DKZ3UBmROBKXURd/EG2kZTtf9dcJtwg5T6rDoalU5Ge5NI
KiNxO6YF1GqU00l/5GGGkj9UrVnNOpfj6I3rnUu42rko70b/lmRuQjA3Z3ZHhynyHypQIlHHh2G9
pSKjvZFTeyT+kiHw3qFheeShihKSftKxtdg2YL0LEg8tubuILR7KV/Q6WcXlFGUfc0IZj8xp+OLy
oK7nNGy8scA0zz4hg9ls6TTh9VmhVkq8kqKhZHCW3jVGiSAN/S+fT7QZR1Zg27BppdZm3ByFmwmT
tuJNNanviMjMH4IHTgLWpZopwJ75aniBPgUqyVHW1ej9VGsEVjAQnWybCfnWR9onvUzFLzlNKZQL
alhN6ZkTb195GC6d/LkEQ2GtJF6+YWEO/0mIVhv6NScwZKe1UrPX3wD5V2X8jPp8KCdAachKwnbf
2NJsDrWS5r7Uqa5/w4WeeuvolX1OvkpJ7cdR1vCg/V8/bjLQjYWZxOMVRdQFWwq5hjIrciqP+md0
oFYHbjnTUvJ9kwrTwnbqv3wJBo217Jw4uKEquOryP5cN6//2R9Ba7c9nax+KWec1QnSNCSKMEpT7
aL5rRcOUjmZQnHKgHMxLJ32gWyItScQl3cU2CqedzrrLMaayD/KxgxIfu0tMzWPJ02+NYVJhQ2vc
SgccEryeEfOnGZ7HHKqMogSdtrkS+ngKnbxbqpuzQxmKQ1xu9tVldmQtl2u5yZrAiu9YhUfO9ccX
+ywuLfVmDnUeAUfjUL8Bkd6SBsJlWZ//2TFsnYa+b8dWdyJMMlZPi8KnCC6ociI30KRUBAr6rt5e
ycXt/ES9v309WRDOKQsODwvqSnFgJkpGwVaRyS8gRe7+mbuBoqlBxiws15LPr1I0nG45umsKzT+p
3la/lvfmW1Cy+MhYyUHSC3KrN2m0iO30efwVD6o6me1h2UvYSbL6HmUrfUNYq/551tDJxpqv9E6b
0tKPCMj5ZlbnXTupw/X8L9ImvWCYjnoO14k46FzGJaA/uekWQp4RGw4uMa2Wc12bsD4lT3WsFCy7
HtpqbieeB1kILqspeGxksDC2sWyrdxjTY4ZpwwP9j3v4RqHrnLrJs8TxvQraULNTuCIb3gWqnJaT
qFpXclCDNRyEKKe2ntvml8IVlSyt0TWYzV3LubfGN3/+L6b62i40uPqwOQVenDnBbuzea6TkdbzK
QUqUIysYI3mehCStJIWhjTdYtQgLx1WoCt53MCYqfkbWlnZp8RDsCHnCQXijArWIcFrv665nlUdO
exM8X/e6q5IoPIhQc4kZG0grd3OjyJoUo5v2RpdZatV7r6qW3d2wJMWzNoTb5ers/VeGIQS3njuk
fMzAs7kCt+UgfSMzgZPtJyD9wGGG97tOAW+9djfmz5glhP6PTpia5rLUTfcgS86Zeg2/369YlsAf
OhAQfQDFB17oO2C5sc+kHEWeS+tuO1jCxoFZ7fDw0ZppHJBKdxdjLBLKmDk9OeuBZWTGYOmZ/qyj
veOg14lK44v+KT0ohsAwPWPszg5C5eeRmYg4Ve3fZMIGalaOvcTzeg0fomFWE5aRoi6/A+DoH9CX
xMH7PjAPQQJbGFXr6bEzXHhQ4Rn3tMWKdPtVtcARwfDYRHBLb2lKCf6uDLQlwMQCO667WXeYAZd5
SYKvKE6Ag9WcugltQAX3cPh6WMQsnxvuRELNKuIuAUXCG/jC+ENFkGu8xjCvq3NO5I+QcbzhO28k
U3EWE6VC/YE0Du+ds/3ZNajiaBPlhV65Qy3C9oJOesdBT3i1qm6O/8TBVga4cHhaarddfN7dTpA6
MZL+3yoKQS43bMKcGnfFxiKmFCKp3FQLxecGGwAUJcTf+K9CVEipWTmHagfB6V5XQWyYIJSl8uR+
MKPqKXdD7o8XMQaiI7qH8IByp1gsDiBohtVL9uhML9iHM/E1C1fQ8q2B8TqpQQrLSWcjAnrtmwPf
JCBaUV3GcDjBlgXXeCgDOLEHFomg8LlVaRA/95gUzV2zqukSm6VB3gX8SWI7CQJZoNsBgjtUe3FC
7y7nGNZDr04q7rxL/1Sa26qFtg67QGVeBWaFiQxzt7U1L1JEgp30+rQD4lWR4oeqpWuweSy5OJWm
f7dBj+IuwEQs9K5oN1rvmMU0Vj0x0+ik/lMet29zSZYYLURGfERMDFUqYcZOCzPjK82a3EDgG3Tw
W1mz3BrAjqX5UNUDiTvk35NFxA0dAsaTW8eLx5U3ZYZYXklZ+Rt3z0Nio8Uf/d2plSi8u4St4YnR
+zg7r5ZeYfTR+GdUMFyZkVxHPLc+RUvSzx0BmKLAnJKZ6II/DBFSShG9fYw8PuC/hQr3NWXfzi6/
tguaCr/gxgKHiPr9CW1vzshnI6Y67I80BjYZgPa9jkImczu5v1OLK+S+plVUE4P9PRM5fYUyrNfu
sxIEIoMXfFT12ljYaqp/ovVindjoQtMJzGfiS7+Rm2Ru+qsVaRV/E40aqX4tMc4IiI7ZE525Thrj
wx9wzzMfTMg21XEOqFZiSLDRGDEnW8AYMTnJXaSb4e3YgF11D/hs8qj51YWDb4t/ozg9AkYJ0Skg
JF3THCsO3eoa4kMn6UHD6HcC2eaAHRftKAUxPciniZ1fd2sEnVNFIVO8U1lGFueNgEBtr08FEko7
jXUB5F4Ro3MOJZBztYhR/ub7b0d+SSzYeU0d7sVOz0mT2JC7YCqtQEVCaQR9xSfO4KApskeerUqu
Q9EVF2Yz58uRGFCYgnrG6gMSCUh9QtYsYFgmdcqU6oWEf0ZRejHU42Ab3dKjTpNpy6Dwj7SZU2ct
VVi3HaHS0sDSJfA+Plgsjw/l1vljQCK9ZWnxsXd1/P5PsLWwSrgC9ul+lYn7dmzYm7nwhBkdpQjG
1o5aT99VIh16beOElk8t41X2G0KkemIVC23V6xhyph6ROYAcE2JDa6DUJwDGtyFcIOMif5za8JxN
H7JbkGFRb/mk9EodiHixojDXz3IGUz+MIPjVUVvv6HmmLVL48fYhn+6Cg+Ae7oXWhqrXgS3UgQ8s
iLQoPVbHoN56gUm9f16sgHm+1DydPg2NAvxN4eQASwcQN+Y4FyrHRmzIz82whaIEkO/LS6RY4pxN
xpORamP6wBh6MAcXrJdUk5iznkXNkfPDh6lQd14jlDy2KvZC5XK/sxEO1dIfOuIT2IAQuh8sh6L3
+LkSNEoaly3wrSJA1YT0xWw/+r0J8BsLVEKJ2RRuEoww/x+Mbq4zCkXXuafjQ5vSnKdve6oAUmcC
LiWWCehn9O4JyAkTgizkzc5YOZNWrdP2mSohC7w0+b3e8u8Fobo6VyvbDGgz1tZJ2q9zcCoFTW2g
YovvkmKyhwpY9zld8LeFSnZe9uwLpA/1MeL5aVyxKjPVsDsbAvJ3KvYz1/bQ6JfsGQfD2XCPtjaa
0fxjeR4xB454rOIzwBXhl5zX0vu37W1BWsxBhPTw5oOR+yp2PFtxn2puaJvMsDIuYIffBkpypRh8
33bwxT/Q1oYEsjgp4VEVarLsmcrtwRvXQCPRrpeSXPSKsVFLnYxbbb9Ly5y2lO05lICfMtzyeUqV
aGxxwKnonKkebcJgD99oeHipPzW4jkU7IvY4RherxEkwU775pE9hR/isIa9dbHcWnjKaIh0syBn6
si5k2VeBUmBEU2mBrMNuUMGbVbif4mw3I35+AB8D3grK+8/+BQ2cCVEFv0I9KUXQBgxcbveoCk6V
h5o3DYMJ/JWgSB7O7LxPtw/6TtGRgGc4nuWYMCo1rrBnnuEZyjaR9kJ4Di/AV+dKuQFNneSNqOmz
0cmDHMyysoh5kkwgTi3JImGk/rlp8AGx4YqmO5vYGXYjRWNba/DBo/8EA1Fmq3CeqXRmKFfjeHTG
/wnW8isiiB+FJLM6a4r/MFSPZJC1MTQ3JP5M1FPnRnC8zt5Nne/XFnsZQBc2NM/nWk8jxrgjU+Gv
9HgAOb7eg7H0fDzbN1uDa1rdleSG+orE9hiBrkK/OO0xcbcYfZTlpADixKnnnOxC5xOAoj+xl4oW
fO8Vc0KH8BrxKkZTDnNmgXMEYIUF0QnwkMjXIIX6BZLvGbe1VM8GTLz+6HYydvfhvTgVPKDWADqa
+GZqMtNJuXF2VxMWviw81nzVDBqUEUeOQbHNhERj6e58gXISbq8IMJ+ivsFJi4nt/muMrdohVf96
//luV02TMeeYA+NNQGV91rnxkxfxBY4to1icP2s8DTo6IxnLKc9sqUabnaX97F2nM+/QuPGQg5gJ
L9tt/7Tvc2r8/iDoL4TIeZnfUcyjNsYsfVt8GPY1QYcDyAX6oNbdeTmarqxHBxJ7ZHUKEqEM1x0M
uD+qZ6pD6hp0XkBYxcyVhVNUfQlyjeV5/WKCv6UjVfqnFjGsN8eX16ZV3pBgVQveFpfPO7POBvIp
+GKNKmb/f8tZ6C4LJCWeMtJBJdzJn1ZQITAzxvgkCYVZ6AIFmTMtR7S2Bt2kmjEagYo8jcca7Nla
nRhTQZYJ/06JoVCZVzuaRUxqV/aSevK2vQnQj6c9NRN0M1LQ9tlDcVw6hqick4LHKu13fxh00xcT
3HWXpzc1+PuwbUG8YHg3CC+esd2hpvlef7qyYXq5Fxh42daNiKFtn13tSIqA0kxYLrM5Ff6s9xhw
9j3EMlmkxdjSfeIH8IdU7WG7z1fUbCNmhqgiz0u1g0W4KJa1hGFmRbsJF7QEx7iT7y5uQSzxDhP8
JIWn2Sews4CkQSFW7a2HHQeiTzvK/FNrhLgRrH9ZsOUXHayw3kSXkE4GZgOPgAaF6oFoVMEJAjOU
gNMH6dknxWVkQ4mp+kLxSeRxJ/nrWEskseLruY9EdPAw2WCJugw5f85/IOwX7l1CSADkiS6kvD8c
3MIUOp5yQM0SZDegEMpPUwIO3rB0AjKThrH2obRZs/UUbJnUKs/TB4SQ+euTKG4LWBBkRg1t1LhV
e+CD4VovYV5Byi+mqTzYdqrhtl26Cmstki6WGznoU3NM8gjclTNDUJfuoxgEBTXgxuyHAhuTrR8A
cWV6DcEFRNdfPLNkInARFZH+xVlNPiQHu4OglM5Xxqu1xGr0ScC5obR5qx/1tdcAL4KFDf+1+aTC
2cR+C5lh2Qlwll8vdPkG4ROu+7alB9IP5vaT7W2/wp4kSnsy+fIlLwfFU3U//GA1K7RaNuotXs7F
xW16sv9gXeJwP0zWF8kItcuB/1Ds9MvnZ2DgCvagOiR9NmKBCsWxnt7mI2vCWR9jIpKUBsO7v+AM
uRp4dA4oIiTtRNwC4+3qb+jIxSomxhSelxUoUClI9wPXysY3ACgC+nlDPnuPfYgDNRcq85uIFBu5
4pRhGeWwFJRuC8kaIhC6s8mB+eR2mi5zcFseaefGGCbvbvedzgpFuAntps7rPOQvj7Fmn3IpjU+V
p46Qezb22U9vUQCy7vXHbPoIWZt+NROHfi31UTqkKORIHFnmdM7+oLDfh6/h/5Y+diEcGITG9WDx
kxor+7lW2ezp8/Z4dRbVmD10mgK0uIGp8v1WpWWs+VgP96oaxm4oKoz6hNgzzDazzh+Hk/nDJBRN
tNUOXJZaNxx3g5yYzy/OqIxdIlHGMOl8/RH8VR5+SR35C+J9787pLzpbu/xNnjXvgEgIUkcZ2XDN
Gt1erksv7m/7KGVhDLS2vg/a2jUtHgMg2V8DbzfEjpMLRBYZINnwb1yB/WJ/2/FQbxXUfV9mOSYF
deB85K7bkKcvw5OZK+TvKTslwr21vNxlCf0koIUrJGWhRjfAwnFn2aXMhNp1Vb59S+IaJ/KAUqz6
ATWf6twovxVE3oH6X/7SRYxnDzIq5D/btQb06hUYTkvuOw+dMQ42ZeBP/RiOqh3aBrcYswr8BJnR
QUXbJx0GqgFnEBpWKxDLAKiJQ/Yst5cnbE09s8mT39Pty8IiPSiKwbO1sYBZl7ZusU4LQxKtl5Tw
rM0TdSQVEhnpwWMUzHtJseschBKzui5maGohItU/gSqu5CX+ahaJxVWYssRYqUhdpJY3DCOvDUVT
j7TmfXPr2aussU3WQcwIz0NJd+c7aDPbd+3ZSEwmnoa0vOCya1vltcoZzF8DTDn1QWkr8cD19Fq5
Rs6ifA8beI56tiB3Z0W6jbLidj3WD+GTQ6W1MXUG0HDDVwuheWK6v55V689CjqtrjbFoObcW4e4g
YidCGEnt4HhorVf66WJm4rwxmxuoIeQHol7YNFpiC7FpB7INPCSAnEXhoNur8Dxzlma3paZMXXmO
4o5aWyS182g4hZhyGDztyyOApdcyiXaDADek4n6YGRajn1hand9yn5FJaszlSa/Y91hEjW072UwV
sjqsxXQHOuxoG2X+QnPxLozpAlOi8SOwsi6e4Uz0RJLazPnOPpj3MSug9kaXARVxkICwyRXFF6Hp
qbFg7SbwhzuhV+GNZkkhtl/RPLA2xUTV2w7oS3UWRLuIv7a3uIfcsHxQaQHERVA8nHvoPYKdt3gs
NKQA9CVj3G6zP2G3vaJA6BcGoTn7LainO6kfpYfugK9SkdsuehVfLsTh5jzGBJF6WZ3rLcG7Yt05
kPPGYb4Fhn1OMYEMhO3HvCLd4LHkgO5G2B31RV9oBLqr+Dp/cUO1EnDURht0B/tmsIXUTLK9PC+x
IvHTS9UCFTImp722i/TtpJcqO79G3JKffrqGTrQDQ2n9F3xePb0nh9NcpGIGYiL42mP2aoiYJKRA
8yjncsLDcFXljoNfPCKGNTLh8ntmX3Fctj+EsPFSV0NOzr/uMPUATghyLsjBHhqpB4oPmfDjvV1t
xiG83e8f3kBUinafr67nQVdfjL8JmBSOBtrX/jlAzFt7GEOTT10Zs7+JaOxBQoL6xDzDdC1nbAz3
//wX51bHKYu0Z7tJBLT8XR0I0JDU5+OWyqVxfzZjMghKhTPDzVxsXVMxVKfw0sKYriGz9Z3j1Po+
FpqTaJDBDTxfYL6V07Bt/jYrxhAHGnOqb+aOMQNq6Fe0FvpNfpZYkZFgZcfqiEvVacM4v+VCrETt
2/GhQLa8Yp92CtutA5Mwpt4FyGoVtRxs5QUw/8tv0EYEFsVe3NPTXSbcx7EnMgB8eyftCRSXriEg
Y7sTN/+dwzTIvQyuV8ysK9h4VgecEK726n9+/hGyN/k/I+3Vv8NgbB4Hjk1YxzYifJ3XFOs5KObm
fl1DI1QI/KvO6UXmqspVKCUaEtHBJoCnR3rzfNGGFjSD2NlmvgWvnd7sHBybS78RSQvU+uHoLjZq
PA4dCzIVIkkRx++wXws5q4qwGWTcwA1Cf45ZldEVnlPbaiEqM+lF0aZNCamdf/FlbCWSmRY9nu0L
McS6Bh0aNz/yOtDnL8Cq/p6OhB2DQBBskLz687HWxf130taQbCkcZZ7YYTl8IdGdigFLDCeqlXS7
k3bAmv6CsPdlgMZNUhktgYFYmFPnl42RevE3bnqRueZxq8VSL37IG5aeEy3UIDY9usbCwZVTqQE2
YJYadNxXn1d3nxfy3rmdNnMQq1WJXS8Tdn35or4uB1HGu5EnNP5XmqxYZeVRx2atu8d6udzoVGRG
oIajT2oU20y1LS+0Rdx8wsNNUJIfZjh9ruJFExz/w744hxrps8wS18ykKP0KuQptnDV1CoMBfQPz
ubakolWGceUI7lqaFdF6Ll5aIWRTSxAd23ciz+ICZVDOuTkpMP99ms+vyjcRq2mBBdYA4Kg+Ho+z
DWhAfEx4q/jqBoigZ2fXrsI0ioluhgzKocnr1qahIzET19gC+z/zM99Od554BHRsgarT1Z1NCC1m
UiaPsJaDzJ1u+iqy96O6mjhPUxrDsvpgbFpKvufdbgKBfwktTJYlJSM9WoOjxHToLOQGw6fivVnI
MReFtRW+BRNjzuMJBCp83mrkRoIGeRAAfu2xXA5h/zODfx3elDVHyMxC47rc9yo5YMtxDfkQB2te
IncBbzwhLGRDyMj0acmucrHK8jctbkM0+GHdmYyHkGLQbHBmmBjRTg2J5rxxEJmU+roh6tmrSyBe
rP1ktvJ+yoKOfz7kwwzaAOYbPJBqI6ysUPRTNKiC7XAogEACUO4SUckqb2KV6WoN28BWsvXzzqfn
37+L1fOELi0Mn6dO9fUDkQg+lyuExx/pFBCMxSU/2xxby5n/XS+xh82EBcwUe9lHryP/A4oFvMxE
puDMeam00ueFFB4QuvTXIpyITQG0v14jiZd8zQhA4D+SLcr9kp+I2OtfUS8HQLNfZwL37Gun/flR
mNrhyuD32y35PatJsMVbfOQm8kR7aMubrUH5qDaoCHpT4Adgmdft9YGr2BlDWIonJB3fP1U14hhI
rfNNOul5gZ54JqtQE4lE9F1YqCle7s5sC3ZD+jYPFqrLa7EipJVqOqsnwBcYWnwt3jpUwIA7iUte
DeKeHlVOIWz0L8olM0B/rGrYTgUJ3TKO+Is23ATrcbGnTjZnrUYsg/V7iw7EGOE2sbMuAT7u2mKo
TpIw/9n6OltSjUxCU5tkaYjoeq/GcyMPAaU8SlFfv0dcaAOdIGeoG50hxROtkElhvgoAveo8ooXP
D9SShdsFYa3dVkyuA6co5pSCwMCbb7Bb/VDxiOIgfkRkv0G/ED8BE69kGeO6PJmqCcxwFKJ9Xc82
mTG/Xd3bsEk53FvkMXXBth+QJd9DaT3MExiZKXjhXDkO97zLgSqlbVEPC1LRni87Pz93uwTMt5Sk
q0WbGtw2OYOFUWcrCIX0l21Hw5VdX+2hj+SW7ZLksgx9lHteq+qYNRQZHWy3FetaIkijIdFjipwS
TXEoTAKYB8+uE9+CwhuuD3n+7Xem2aSgkIMBRiGzpDOxRxA6MFaoA/hplBCt1tdHyUAgUb+lMFe2
gWF0cKDtAgCFrVGjaAvHejD7g1ITvUaz4aAr0VNvYu7X3wmkD50+THbbfPBS62+1O/k/aM7ykWT9
9LONVLgiPcogmu0758KezfqlWhq17TP+zQEmaio8GJPBLmENkxZ56imN+tH+C4Ozh1fzQcDUq4go
dUtrlQfngXXyvReC+R5mRGupSJ/Y1t3E0FBShJ0yk2G1mX0vpl1YDUDkLjX7mNacP8f+88yhh6vI
EXCPOwe+9Y+zY/WQi1WTUFU9sMSP+E8/6GGjsMz+oLtcicGwEqKpJYWzPJvQ8KlONuSCdNguoIjS
GS88KaIjvahwAXdKZNXUyTAaGitT9lqzcIO5fuOB77P/PCv8PpCrKu8bJFFPUX0LmXqfbv7r0yRs
eSt9q2dHNfMzXgVoQd/SbE3+enDuL9/HAcwg1NlgsBIoxCA/pIuAtQiPssvK6rF2iWoCfuuO2/CU
PjT6G9QGlvsyaP1ub2csnDAKOE524dqjvCi2AQ4dQV2XKh6TE+ys0BMZdg+GEQSFP+SK64Med1oz
rtJtmyJtFjdoPoNkUPw7MS7R9l0YT7pIdBQAe6rG6qoTWOSakFiLweWpT4JnK/TAwr6fUIFTX/9i
AyAV8WwREMrVyak691xtOEwl9gAHSgI+CQFpuks17pEcmUqhFo72/fEJnYEUPpnqjslmQ3t7J0Ft
bg2HPBTF41eZhKSG+8tW5R5oOvMh4BbVuhRjkZHwkgP4QLSx+QHjTKyRlPNs7/VSuDnSbNnCxMba
9VMGM+RouneQzVyCKvtzDDp7bKZ6k5kVkMWJSnUq8fdWw0Bka2F20NCbzMFE02mMfC8jWAPWxfVq
JqwnVbf+bdf0BeUtHvyfgo5oEA4XfbSZimE33x6ajLnaMzLe/7Xf4thttiiVGzXFgFSPwKcFQq22
d2dvTocC24isx0D0tjG6lT7j284VFQp5GVowwYigHjxCVfWm0sOdbel0fcvIs6mI1lmVUCSXmkcK
r4l5H//jWSFUaTvFjWvq/Ok9bJu83TLIZYZjAlDEHkBAnY0WpNsSgy3OpOCkrWdk+An60rCNSWq/
FS00YraidFXHRsGFHQJLHCWga71oIj/6teBx9oIeiod2tjtLKwLa8Ixb0Y+gncddI8V/f+1hbP4z
O2vs/J3YxB8rGDuJnEj5UGn58qBEPHn0pbbEJDw1xwHgEA7/HQXO7yn+OKOWgYUlc3xloBz3YKli
kgcFkIcGU/UC0rULL8ZtozUqqZaqwCK+8+YTl+TZtJps0J2jzfcNEueDfX8vQrAL3UQlByAyqcY4
ckJyoZaHdiqe3W9SkCotGemS/VOySOD2kBt3ML01KBmz4BPCyTSUgl8oLKUOrw63CpQ0BNm8M4Qn
J/EOX0KWceu3N7PBFLG4/2BAbn4T3rKJcIt96Jl+yIVUIfX/dDntltUsJZ6uwjZLTTSzOqAggEF9
XW066h9NGKSvx3CCNHsMV6s8WwgR4nPn5C7KsQGQg5+QXCRQDEymQhpu3h5RKd14qoWpj9qk2Ycz
vrh9QtcACA8rGPQisArBepY8DrdBBbg8P4NeRBbMfcZG6CpquZQVdmfi+cTBUZ7bsZqfusia57gB
1NhNYstaACHB/ekgJhuQ2JjnhkNsGsOoQMLaO9HQFesMbQMllKPtBwi4OPA91RT448SY36Pei4OB
iOu435Vejpt1oWNFk8mgCZpMPNFF54bqHYODMj4ObCDmkRxtRUlFaJyWU6aVjYLcGRWaTWx0Np6z
0AKv/BrcVTV3GtjZEtvguuHiwP2FJTNznKzh+q+8MhCqXl/ITRAMocGwgOqFLL9ABlzvJAmvPe2f
8842xvS/ke5S1Wz2HcDsJvpLiPUA5yrX6NMqvk0+TzHqcseA9YDfKC/ytw4xHglw30pW8rt5fsRo
V9UuY1Ye6xzXqgHBgkA1mleCYvSlG/uHZnXUl+F7s//FseB7gu+xjaulJu1eV3cTr8Kinv//Irzj
Z/6RMIGUUqeW8HRJy0JPQt+RijgljMeHMcXjflOqU0ClkPiUIeFF5aD9D4GCGtPgZB8YxA0Yu+r+
7gE15XXcRAYqgnqgGoCSmkPiZ30aNheR22Hrbtn6qAqVNdmC7kWZTq1as2/o+CbivhRgeGZWGtct
h85L87CihJiRHnKuLyzqk01fyoRyssRx7bHfJD7GwHoxeBPCX/Ldl4kXdyZCbSTOlfn8ucZyAyCa
K3sBhDnjKvrbFPYp9YtrOye7rgKykAeJdJWoKoBWFW5uG7MYbgH7mgaJgDyzcnLpcJengDi5QGEL
NYnEHc3PNbLj51fWKwjDHzJxCUUKggmC0HHAY5Zd/NPKss6OW0xU7IBmfgfxo73uZC/KxkOeZ2gk
/xPpaufUeULGj5CqbzzIrAVtlQKYY1lpSfjo5yzanWJAC3fuaGkLdyZJAeZN6x3OGlM9917A+Gtl
KryAHvZj7N+Av966DsoFQpTtYGkFxvlA2AbgMC8j7r9t/M3Sx4UJDzzO27wvDiwnWX+TcedJgWYp
3czHzk0uy/pyqOt04Dx9n68jsxgPWufq8zjf0KOtork81/vc9qe+RafK5CselU6vSVvW9PEhZqUA
/7Lhm3AsEdNIgetOm9sF8gXNrNZ1a01/GoZiqd2Mmmw/vcROj4Rfm4vTgkFwzJ/9PiMWgLACu7sB
+zf5Mo0Iui1/5KXizplu/O3JsH2LI/YJeWH9ivJiFtjQ/YZ9nuNt+1UR/cVqdHc8UpSkruhFiFCQ
DCRNEx/pnIa8U4HILy14LilyitbuzWMUWlUL3kjygq4RzTjEaN69S1vmIrRcH7PvRKFxOCbw9Xeo
wD6DNXUurxMCIxZe3nWuODR1S6hxbqlf82d1ClalANdXLeXa6QP9ylFRuJkF9l2fWB5QfqYhRN6Q
E4ZCbYKHFrXRbPAl3lqwa6qMGxnybfF0X9HP3K+9iPlWCq05SM5oXn8bxVm+1ugzC/Y3Tjnzid3m
BWjb2+3I5RtLgF6FtZ1LzQcHTouSBaWa6NF9YV5ySn27FJXxYwcRTFTN+v4nsWasMo06aHTIy4Eb
lqhhNpE6aLx8d4eyird/7iXNlY5JqMtEsmsJ/tLDfdUO8HEt84eFsU7zq4C6Y70a/OkIxvorBtfI
ohCcIwTFGOZle4W9LF0FxbTjGry6k58HdK55VB8KL12tpF0P9+1xNO3VImk+HDGj0h8Paj7QCZHt
xg7c7VZj/8w+1l4rNQ1GYbOSIkm0ZvaSQ9bgUXPntAKBu9YfQrthmiF0sGZ+GjQhFySE++fKR3Bs
P7llREbGGvLOJqwxRfCKP+lKiLhVoV1aVK3rj/MT85+Z7knIDhuq9x/v9JQiho5ZZnZS01jtQyRe
Im9mq+yOvfqTuB+o2sE9ru4eMBJZpd2cEAvKKay6QTmLE77p4cxk5UH39xuP7XO0go8+Ph1JAb4C
DqW/ObAe9AMzGxbYzWagV1Nsmb88E5UchQOvkZCA0Y8yCiZgeE3sNwd9eTvVUD/uxm731xLFTkAx
rfy410KodTx0qN+gADOcMXiRB77JtstM62tnNruzgcLU2+tmKHJOes3nCZqjIlZTdzDenHtg1+My
tyRk25fPJuWoijxmhuJOjIHtNW3R7ZMfdWAEq7M3NjmTtSWHt6BKjUxbxDYjJEcSELcnjhaOzIP7
boRv33g/zs/kuBJjAR3AoQGOeZZFnvo0BHJcEjh03pITnTTVfRIk5zk7X19fAh7zDUCNEo3kz3hB
TzMq3Kh7WAxxg3Hg9Z70MAR2AQD6DX/+5B/E8c/S6ZyLTl+iLX135Hny3efptIzAE70Ir7g/48bv
d/0zwGW7x8Y0kbBCbkxNwai7msyu6uzUSUcGZlK6f26atARym0aeQnNqF6PLu82dme7NsbthCr6a
spB5WpYRhNOsDCYOfgZVmeFp8TlcukPmp9f/hYST0DnXfNJvW3Hhb+8ci0cMPV048Fk3b9oQ+XGs
phiGAVZg0gdKVuiTs+OY11+6hjhg1VtoZYN2KYIQcDHsikf+bhZCqjMSL/XUfcUJTT8k37n0eZCK
FiBmI95IHX/Q2eEROin5fxRByhsv2asz5ZbR+ANhwkZAAnA8IiRj39feFmeu7Ol23ouPF9FvUNfn
DBzXfQzeX2VcjFySQ/LNT763Jt+WF7qeygmVWJaDKYY7D4l/gvSqlHEQ0Kn3/I9cdiDJqttUAC3A
gIJi+2oepeqSgulkxi2w5747hrDlpFsI4lgN143hu9tDHLovPxeckcxlAp3X++v7VV9ECP26Mv2f
IVMZhsdKAN8b6Op1spN3Qyn3lnrPWXJuZryOzAFI/hfz0UnkTpO53Uu1VRvEeVG37VurgW84uE6C
5RiVoOtuuhtiHe18kbikF4X8T5qpe0cgJCLFizC6J7klxdfbTdPl5KdIAz9685dAZ6uh2SNPT1tw
G4mPPykofuLPcg4j/H3/SNq0SlbQngRlwtW0DHB7rvwiKRYxi4mYX+esEFdUEkMPb+V26LoHIUL1
dG8bnqjY/gScbQldBqcbKJlu6CXOvBMxPUdT+VUTJXgQPVfqppJyMLCSOJRlO+FntZGFxjUlG7LM
0iXnlxuxNata5sa+0RUvz+YHCgpqFfaIOh5Vuf42pIuJOdYYdZ7Gq2Kr/EITQhH9S2q7ZTJp3miZ
HDQ/oM6Gy3AOQlGn+boI4gWntgDvi7AtyotXPKVsy97kYC4uIC3TrctV2C5+buAKX8N4kCwJ3YHI
CVOCDjSDaMtw4t0HCNEvjsGLFkyAu9elpoayFK7XyeT1NQlhxLOkkMKa1Mrj6GAQEU/tvtg7ICPa
QpLadCFmVTkdOUcumzohrRUjBzL6oup9CQUu8BAanwY54v2qc7Q6Q/++vIG2j1wKODT0C4YXY2v5
93kcRTteHrj7SlZkijzLsRm2FBi1j6y4raGeHWF/bsjg4GSh1BQuUZ2K8EbYKKdlmHJjvQUgaiB8
oONq9tiowLd8OXLXYi5Rz5uTCddjr+0XxS7Uo2/mKI72h8yRAOV0GftOZmK0lh9hytoUxwXbCQhd
FFZaWU+oJeKtX+KW6uuQkwJgWujotpzu9Jl232YjYAPLLE6OS9RxtkMtMc51MF4wRTFl3aFeXWkJ
ibND4RIguRda+Achs3llDoozgJqfuPWXRmupocr3G1lwgM5ldg8qtR/bCANO8vuQpMtbhI4Z/L6q
SWS9PRkQD9trVmUzCZhy0xTXIRiQZCIltNsWv4nZLlhVD2XooL66ehoxpbU2UvgiLO+C/hk24KEm
hZJnbiQV07MCKf2UaWcgsQo7aDbRzo1hzNHvoWBeE6bJrvsTlx4sdvfzTZM8jChbML62KtQZIMRI
UT7lf7PxliCm8RdgCZtkN2WedMapMvkdBy1pYWddiE60q1jey8/0a8B8bo1W5g8EtLEgwmdxugpW
4Q+wOLhJuD92h8fXmJUSOEpzc4IYGpufkV1vyYEpRqGDeAKRhnLl9kuhHUL72yWyLIJnqvj2m/Lg
r82vkSJl2WNBqJZnWvn4OhVusBWVAMYnWSB68RyZA37ei9R92X8LGtyXEvK/jFeZNJ1e2zoQHAzz
xMK5YVkbEAl3C+GgwxcXtCmItnFN3LvXCUbfvAXE2949lPzgzI2DKI8olVV1/tM1FYHlP15/ONYQ
yLXMbS5DjyfjzIremqJZaFO6LxkqWPJcl4Qf5jlDuasWZu63M2zvEHzzluQfyvMyiOuaZiRLymfB
NGNnqqytdYaNaDrz2ydyhO9Uo44C4EVVHok0tS7y2a3xXhJUSg0xtQvS0owtoxxkT/k2cEBBk04y
WV/WBFtHSWDNyow6J3SOmcfK9h0K+8sCMV6j4Hq4JKx1gqh4/h44Ls++YI8EnUdBZ2Dj/2PI3fob
2Qjr1gU0rkbfcvmcld1F1hSWSNKcOIUop/BkIOSiHiW65LX49tW6WjbAmSJv8sx2SvMgxYyZOSjd
AEM5J9zT6G9Ukxl+ytg3hjKcacTHIkjxxPPC3DqO23zaya80NNLGh2PIc1NkOPkjyK/1MJxmPWLi
j2NBFThRL1HzgGM4DJBIHHnhWLrAz6AjNEPAyRTW+pQQa5uGX4piZYMl6dvmpnwEtNLSxoqaLRKp
54Kt+9Zu6VoMTnOnFL2cRYDZIBaBFcwrsFuVHfGHmoX4c2D9G6GVtY8WhBX1hhIUw6T23SwPEVvY
jncvufvlydlD+IBKjaYifFnbNU4Tz22WLtjq3R+5CGCz+LKeGsR9HA1MLKIe6McOhfwV5ySBT7d4
/QJoLOTCzp9SbUQAfZ6tZU3U+7PXuzZxKcFnlcTCDhNt5NiBT7l+c6MXgSSq1vFI3jz4yGUBwWC1
hAcCwQYp+j907K+vj3/6bQCG8Y5q74r+dMdi3ld+V5mJHkLEY0z+6k9K+fREzZEYm/7FjuTLlPQU
c3bSJAhCgy5oH2wIkx+H5pCA/eSIiLTNRpOrcOJTNDWXZkn5w+BZOECppuxrQ0lxpPukFP9vMd5v
gKTtJj6AjIunAMNWN5GlgPGG+dDR64N4D6I7BAqGJn/CKPJSB6jYh6gCVA8ukaTHbkFgTGOGw7nC
4geIyX5FBAcX5I4XvCSZHONlnVbyAHAiHEj53gZLBHDHPFvk1o65gSrGSYd4kpk4hlelpe72D4R9
hiHr6QjkFQDPFiuINCVgyhYV2a0cRHN+tr/9FTtnFlI9PMfrgr0EE8mzPMcaNUiBv/2reRgmlmLq
psN95F3GceRm3+NvQEwnw1hY7C4Qrrisx9PoRKR3On30PYZiv2ztsOaOO7XRvNScLuvSddOG12IR
Tlmsan3zlWPr3IpkOmHwLXtvGDSQVTk8dFi1ePM8mZkkKwGrAg//fG61bWWEefvLbyqdPKfYEnxa
gLmeIj0Yz8gfUCAibH1sbe1SbMaDKyri2qHOCxPHppN5jntOTvQ5OfPP5/3JuDQ2Fr4xU8OhfBp6
e2y0vUMX7xJ2hIxXY0KpGaBcc9MQFAZ6xyuFEaoql1YDXmmn51Koib8aUb2TPxsHY/QsU4IuuPpr
8GcgL5U8MFz98qsM7GzJ5NXclq5BNu99Dk68WjeXt8wU4EG2EETGAA55lx96tTimsj2qqa7+nhEe
M2mpZVfbc8it5Dmi0YwtsKLyJYOatbynhx6Wm+IsEz0isDHggftXdEi2nPUWiPukjwSkRhApBqNP
Lsk/P5ao1ncN5+p3o6LdpeiCD0MRXQH6e0nF5rjDJfnzTnjL+sSqat7SmjzAuUDXBdnttQaSa29T
NdrttZZt+b1/byE7/zsWZ+nX1VE7VbRf93CvBj3SwnETPImUs4w8YlCcUEeGTT+mR/xeUXjNuZpZ
OxAhBAa2c10uiAhPkN7C+lj5KhE4hFCKYNRElTFLGHjGLu2Ig+yNz89CDKztgeKvqhPBb1DYlWrV
Uuuq9T7ckJrrmhKcFIYQJrj6Ec4rqAkIsZYudn2K5H0Q3cswsoUZ/vbQMGhY5gHgAQIA/DhO064A
UMI/Y093nxFC6jjxV6Ddl1P5pYrLzC8f3ORo3VZKTj/vLV0PUN1LO0Bk+7iITVMFNykAgFFUpGCT
Ftl80T5cpXjuNtMmVe0CEJly/LeJurB8xyn9IhNMP1ngJpL2hKmuiSwmK2pS8tvG1Oq2vHX6ADR7
MyzId1S0nHxzLEcob6KrWlG+cz6FAdDAGQJtYHlm2NlkaOqb+kJMcgoiqvOa1apT5MKYEWLcX9MX
owYyi5GlbkHUTa+UnDQSNu7y5+QYzRjDizmbiCoUOrXA7Z53L5l6+2bHNquhFkuFORB2vvhRFWWv
OiP71JTQtbLhvKZIDBWIXsffiq0JA+6qadHN78neOdAal1hoU7sjdg3lwyjrfbIYDKmmDZFFhATp
sRcixyUDKtoGwVBq5EKeI8207KfGvKAL/Tuw/1q00HkFSB1Rs4DIfdpx9EYEGnq8HokL/wmJT+VO
zCg9b8mkvSTzCagTzx/SKqKP6Sq/ISQDBsXS0N3SgkWvZVArUrzIlcC0wSqL2dQz7KWXyf+Mz8Bj
78owlvMvImqnmeg6jcIehkUVxcC94alP9ZUlbiJDhnwwhm50rcSeRePtnhauU3nq7ogSxwMPshAw
3AEfj+LQ5DEtUtimKKIqBvPeuXGhGiO8YWyZveKraRFzA68/4UVsduaKLlrcT9zwc6VceYtiSwqB
eM/dv9HQLPRGyjJOovGCHN1z9Pkw3xQunrxs7H4wxyW9AA40YfboVG4sDfZrEWnU0kx/gsOTi78N
DAHZ9HZDqiC4OTU18xIPlX931BOuq4Gp8yV14tFkmNzoq+4mP3cASNvpnPZwcryLVNlMWuJvFgGQ
YSt0WOPpi+fXJH2KPvt4iRAq1dxtOuBySVsqjpM8aavP0oDdQYGMvUARGDlyoSzQJoiH1TPgmEDB
Rq4uGN7+bHJWrMeg/0ql/NGgHcDTRxW4fMkumu5Cadr5Dv4CD6FilFsrUSwH5dSErspH+JlCNK8M
XjrkUWc5rynEp4E1pbPaUwB+FVfIz/QGjd1WYJEkWhmFPNosS4aMjYcdiyKzQYwoVuCvMeaOUKxG
iTHlTIzwl5s9nNXV/gMra0EJ9rIRG/1W7cFbzdKgaf2HN1h22gfWhHKjRP9iwMl1lMQTowochQi/
XNVYwR+zjkpnPzumpwKb6zUBdlXDcDhvu/tXX1G6ajoR/iymsX38dgtFRThaNmdW8J8bjF6yPVf8
teZ9+f84I9mGuzsuhcIzGJPm/KpyTYnYQl0fd4scwP4qyLAI0htwL7t576v7CkRJlx+JAGaEiU+o
TZKCmbguH7zmUOrxVZo2qGCBrwIPKoqHFnN81bM0XXVzCnPOBbR7g0Pc95P+pNqonNpgYhxh6gkX
vKm+dhaGfsUIRr/z6pw9qoj0iNpi6emJt4VqsoQeTa825ljjy+vN1jYyydcXcmMw/7BclzPe3DD9
QwRPh1rH+2aDcTBBceYiUFFN33Joneusmee4OD5cdcLMwSr92g6Z6EMDLpTcB6PMyCzXKjA3dJuo
3XQrdO+4BYMByd4DJI19LRu4uCZ++fCS6WVon6nooEBYFp23BgCFA8iZCYh1JWQpVlNlhKiLSonS
oXWOm64EYpQGK6ZCjzEdKMnKO9LYWJSJa8KV5Xu5SbnXN+P0CVRaI1i/4z2fTWkrejHtYxqI7u/R
F7CeCgBHcJhBgmdBT/ACMPxKW3kf54Ru2JXkl9xznxs9CJAsJ6Z50nedUkqsXzS0Aonh+/Z8KJPf
Dum/4aftv4Pot1CBIg2/K9s94GAhzkg+TQViiLATgFge05mlAn3fepwlv8QYnWPHutDHV5YMmLyK
gn7cdqUZJZpTD6Wb6wjX8S8z4srtVaLgYojMlZ/L3JJIDR0o3NJehLRM1z+M3Z3/Ww5keQHvUTZD
fnlVHay9Hm6wgi3sL6FHDyYDTWVYyzRMoyhCU/fTByidyERq5W705P4kzMnpfwAjWKr3IKfoSN0f
ud3Zhf2gCvVqkc+sVU5rXRiETRWnWEDndexpfIcnXjToIJuHChUbtYnA3rPxIB+kN8HWkI20pBl+
wn0Q2lTmBmCD2/9vmZLhnueQCqs3QLpu3mCiX8g/mbgL9/s/Zvs04FiyuJ3J1eA1kmx4tLf5iH4F
yv35rljM/Pjw3hrx7fkQEECpGEx4CM98iJqLpcf3F6oFUB0ZYbNl+GukVQctH7ZuOnMNsr0RIyFl
EvAjlnMPMakh2JyIg3Di8XHfDg0dtlk55qkCbeNSKl4UyksCL9iKu8geo6XhON6yvh5s4izlmWuH
X78ct7ixTiDN7oUoJXBUuOrhj6/cD0LWQyPKEGIcwUHsD8b3y1OpbeVexZ5eZ+6RLRHyDYrZXGZ3
1RxelGK9lpBKF6wxSVbGHjC4WA6llCF/5jsKivLVTH+pFXLLe/uLwWV8JRovLTBkXeYrtLmGSTJc
yjPH3Pyzf8mHpPDqo2e1NH4LX43mScEZ1g+9Xt3yFxd5Qps+5RWwTACgEWCWsQLgfOM2AqGmMel1
JaMdqOYct8HGdFVwvuDtF8BbGFasYhqyM5bKyiVOzQaRa5UVBPP8BapIngDMta9pgQM7G3EME78T
YuB179+HRQeyqW/f7g0xL+v2tHOAxfqE2po5DM9DivgqadYND4IYbGGTH9lgGpqzgGCYLgm+CxCv
4QRgPUiqejYfTtQJDxc2lRB/UEBjEqjlNCZPLevEyKMJcm72OcaApU5xLQsh66BiwbbMUnolA37i
DwALsQvM2vcYNDnGkR8/0Kvvd3wKQbwkqoMmfb1UsGne7qWA2wjYnTMI9F95oY45QdcoaG0+Osvr
3aQ+tY7UoIROdsCkxeLQrIhChnOl1hAKbJ+IlsdOzydSQ1vuWuNyCjvQWNWA9/y1Az+mDlPG2R3A
CLGv+8vdUzfgMSOgTO1Las1RWNvEHPA5HfaB8E6cvuG1SlCyf9OeYTy6zgCa4QCLxty4DZp1ZbVk
FSUcpmCo5hwQFhASvycIGLst2lO4HmUQjZUKNrUqlygijzpRwaaa4kyejRjnXOReXJ1OQaBMiE6V
fIvn6JxST1bVtfLlBH/Uy9pjMqWL02VG5yC5rh+IB+BRIUpynFqtWbm5gvZLuuYdLW9tCOGTyGFa
gdYqkOQqLh8cjQJ3UekGww+8dAlFQ+A1dtIo2uqidOGI6O1qrzYpySLrZc8Pvoykza3UASTz3P0p
42Ls4s0VyrPOxmxHY98ffcBA0OSmPhuBKN8cQ070nFATc86kDAl8frhpnKegHLUTVyH6kWmpRUKK
e7mOg0LbBFGtlifqIlZILrGr1josmEJnYsJ9c9Rab0TZbtnIYwCO8CbYKuqcSvNUz1FhGqnX6AfJ
BhcoiEJO6pH95/lGsUkDW1D+Ybw4YavDleupmU9nNytpfIxnjJHWfT2LsWQe/We7Z5nty7lzrY0N
ernHNu310lrhVQ97G9rw1z2u2fVaYqQjj9xLEUu2zF8IeSeU+rIeoJqymF+uTdMMrcQZEfrSXNqk
VV61QgryFqGFnusnx39zQUCFlvxSCT2QeHDbThearuL5vQtko6mylUxMreni5onLcL5E4JlCHzJm
afxBIYL7A63d/i30zaMzlv053gli4Ic2ykHSaAYw56OQWD8/SmzW7azMt0hDHcZqnHTiTHjTkNhI
uKon1Ho1Vpi4EhmG2T1dfG0Zcl/QQixzW/bBbuHHWek9WW8ag0vwXgMdjqblhC5tkosNY7FhVDYd
LcbTFiXbXAaParw+/wBrhG0ChYCe/EjYsRkl8wstQM+RLVrRaGI8LBJ/6VPPsMZJ9bKV2cMcKEBD
Ij6B2PlUX7Wi1B13uI8wDXQbm+Yf8UQR7RYOYAMDP9iwBAVhqXmQSCTtYcb/5uy7LiJcqsU+e/QR
+Lf+2MM5uvHxNHD58wxwA/j/Hk8TNexEV14CzCSBezBWGsGWoDwR3JoCjKO/rXJEAptwLEQ3skUd
F3/Sof42Bqig3ygUirTCRXzerbhf9BjR/w4USZn+VczZ4urGpNL5b/kTO/GhRv/0MDw5iv7rAI9D
rQ1uFVunsR9/nXa6PNrOxrsql3wuLwTqf6okD89XWT1VzLwbkpFNjlo5hwdCQsfP3yPCZSPSusHv
l6v/Qn8UgkXJKAXVSO4cnOV9X6vBzab0cZHTHOgFsemrtgmmUQwo3mbdIC3LjlxewJR9R5AWzs/d
+OEdFbG55JwDp7tCWizcjC/Lc4w4xqOPu9sVQkCZea6IApTbH6qljLY5SKOWZEWSVWGRQZ9t+Jxo
BbSYBBC+xOQgpZRxPP57jx218oCEOlKgJ+XfhfZY2g+JZyVv9f+Dd1TkPklhXB5a2snzKt2BNzFG
f0IHx+pSVfElM8iy4Hv+sByT12pLaHZAQPuKRTvX3dAQn2EgEXz4/Ng8aVrVaX56/37hjIjYorbn
hCn2bFU3L/6AvlGu308MxFSO6lRuiuOALrppURwgjG1dUNoXamN+gJvoQzMMizkNrycYdRbQ46gB
OA19NqAEGUxwnmVwDlhSU+ENe/ib75WQWdH1FWICZGWccLSU6ZpAXC8PETWr479J111koQ6eZXza
rt7UA4QAgmm0ihbQ1Qmu+3ACsJEjBMUf4THV3S+6m6mYGhpFRj4i4vMMucW5W3TdQsROT/pnJVA/
FSmbUEAnGfkp7varvLfvIqUa+Tt1y70/l8o4yeeOI4yQkC35n3CQYAWkngzu7NPJZm4AjcBYuWQK
H7IEwDtL7HLoM8r/D35NVAMbIE1sBhMhhUK01O1+0p/eqe/Tt29itdV8Xg9/Eq10Zh0SCRMMzHwd
ZMkk0rYoUD5vMLHB3hGbewEu8rAxxmCxwGiD7VL1UpJ5jdKY5H+UHpEwm2rVJZSm+87UE75FpaYD
s2TptIYoMbiqE2jQYeiJekzIlSwyTb3/PuY0He8D0tp35f/qSwkJJnw4Fskc9tYruNR05vmAqfvg
ZFQhSd06yWZaQDKnwAjouSyEcKQLz3IzSm8TI0skgvPuMOwy1Bb5FwtedtGpcm+HU4cYpQNBKYy1
EKYEHxDnoRcsyB9tZAvFeA+s6prLKktlH17NHG3qk+dYQEQ2hFCs35jy1arbv4tDEemSeyGwTgyS
0xXm7HQqIEOEE67cDbDbrAq9WugIxdZ6S/IS7X8n2sp87rJ43cL7H1KuwvohVluuI3QBEppD1UpK
wC/hAZyuO6KBTnH8bHkOZfixBrY4BraQ7Bc/PkxdR8ECtZgFQNZfLuhwoGkoIRkv425osc9CRW0E
WTgiixM42Bn8FuL58GSd7RKEXQA7jjJeykoI9EU0JuXfZRyo0EvSedMKB9loz9JN22+q9jGW+nCh
scaqrO5qA+Ul0V1HIkLE6uQ8/EH3EaQ7DmuQGMwlm+DWZQiV4j85kX55KA/0tMioMyFL/og9mIyK
DxL4qFz8VI/6SSi2NmmoU/I6KuTHccnDkpL+zx56JPJGfA6b4jo/lURvtIepVM00RZURd7g9P8VW
IvJINf9z2VuQbQsHgNdgeY37QPOwoE0OmDopWFv16eMy5TF7lYY1nsWYQ2U9Ua+Z+QIkQAW5C4jf
oim9haBkKc/xtzxUtegNG+5f3+QCQvTZsBEOxEg+S37wFdDlQe6mivUicoQbEdiGMMod8V1/lulz
TTL28Mz7VqZJvko9K0FAmOQADCk3ZHvm42ocnED7gURbi6JORePfK6CcTVPD/sHy7uy/iTCJUyEi
PJHMp/vSk0birS6+cx/u5Oe8Kygu9AK1k2gpB8Zjj+zAOYa1o8+CBbagRlRmTSDOxq2GwSiMxqR0
b4kUHdAMuOtTv1erybylTMuEVNxBmQzfmB7V3Bjzu0R7xmpyiAIjQthGm48AOHN9aWPz1FqXivCG
OPoftz0VVIAKiCDm25wgKuGWlqYnubuXQAadpIjicoGrPSUrYcMMcHIXtHRKeYRj1+Db2ooHgmSb
YlivhL3e19ormt0JS41U/vsoYBbjpmEQG3x8GeQLCn4MclJN+/X7lLJNy/go/A7lSI6l4qi4uyjt
nW9wKmsZU55bdeUtIMN1Hnx1fcj17TDBSidDW2db7TaH52fB8vZI2mUBJenPM9XJVc5onlItzUp9
EGLcqFdNnSD+gph93ebBN77jIeFP20nISjei05/f4uTAfsga/csJdI9hIMGCPTw5utBdofLb4YCh
ozGIgUCI4WCzqM68HSY5a4Wmf95FPAOFfHmskcVtdORuH7/u5Xsqp+gDbLkxnriuKvH1nw433azr
wf//d+Hhk8Zi5AzLlmr0hGgafc0Hz92RMiAAzCQf+KOmF1sZsDN/pXHuvRS2Eqwz9G3XIyj/4NUW
JgAcMgx8gY/7KWF2FaUo87CWmeIBe//NHABQjYk1IX3eOyo7uNcjaIIJZZGFU23k098qYMBuX1w+
wFyH73p+J1VgbFb/vudGF0zgfZX+dqqKOtm0cD7zRgRwpHMEBT2JAWznGZc081Jpfm+0pId0heFB
Qh2IIYxDoUqRH7jf5jfxX0cz/PslAWO7g5DuLxN/QwH3TKsGSR7430p1ngTTYXLjspm9uByW2CX7
gI/mLl/wTrUL29VkUC6YaKYH5kQwLLY+Yc3CiFYUjQ7d6i/RhYBie1e9JvlT9QoD1EYjODZA+U7Z
QC8x/wDQLk815fvqt5HWYpjcUTeldx3f1RtlV0W9S1pylZRAz0iJbAO6+l9xULMt6Suc9K3Ewx+m
ALo5JFLVng/PhCIXnWB4usFabcvZSYOmIp41gs1o9i+yoTohXv1L/CtXY99pqCkKFp/CjMBDh4ab
PNWGe3YI3y6KG7haRto3PI8DLV5qRcJs9iiLDwNY4W/Hfj16ukottC1aUmTHPtKCwYbk37dWrtQf
ebFNueQc/5taYxmOBIAmbl5pm0ojHYRgZKRsBBgXD+WwXB9uEXKxdKSwVPvdU5R9jT0kHWDd2UgV
Ja3wzzfa7IjH71X1xHiqwdxRANaaSlZuihL1aVuShlAuYO2cv5r36gxyrc3f2GP4iPOyelZCTiRs
lfmWjtDFB0gFOo6J9/iARh6DJOA+BAVwisr6sGqZaYnqQOnk4t8A8V+wbtP8zyIC9Kpg/rpN+LdG
8KckSZyC/aMey9/suoqbmR06zjpbe+agH2mZ9lh06LxHarJDabaf4NyuMjbHncQPmGFLERf+KTbu
IDaLhtXPN2LKDr6A1JHPOUq7CdFFvK4qjjRuBhbZLbD1ZkQRosuKx/DN26AM+xKTpW6YaT9DgzUQ
tRiKunGIZx3q6wDzPPi9Kuwtzg3WkLZslkC5jzl5Uw+csUU/4QFaBth/VPzyFWbS+mrkmW54gHsC
FuUiAf8C4DVacBTuT4gGjRk0Geco9FFQ7ujExA4vwmhiHzDuWsrPUqG1KY1BJ3L/Q2ao3Th0EPK9
6IlzDDWWAmEsiddO2GuzGtlZX3erntME/gLyGLBbJ2XniObEHJDrvBVHa3kOAg7t6gf5uGeDN2zU
6QlSPMoPcTcL3mqenhSjUf7Wzi7HKYCaHkGX8+9bmfVwG6imlpjcTHdGZMErJA4sdsJjgM0d6lIp
FSuEMwlDLS941bb0qVgmpCIoGuerWc8ECXfz81uMowF9bDnpldi6Ww6rAKBxfCcHOPuJtIXE6U+A
mzaovQBIgcYFOGtkJDtXqfzvL4aWzOLj7H4Pbt+t3ebCamgNkE1SUUI6jDOm0/Cy+TXk4riDMbKz
l9SWHxyYos8JAGuCDhT30jIsrzN08R7DwO+FMZDdLZPzi2e2HxZ3dTcJ7vMAUQcREVevk9mIptGQ
Gqv0In7EvaymKQId1YPLVQWyd0rxryCs4T9sK51eeNNsLKftLng9H/0Q7HdeGnljXmNFr0Lya6+/
hTQHmbxljSiMYuPFajM0O5WCb/UreZK9PT15080wpqqcWPsv+LSxosBCbJrBD2vDUkvvHDtHrvXS
DbCm5smI4fve/+FDDPpR7gdKpCHnQTyfxt25NtIQR+Oxhj1434Xsks6EliUP/Ui5IFfjWlzsmr20
PNfbrl81KigxT5oD1GiOF57BtyL17OEZVYNk8zwYmJd2Kx90l7GuaPW4cZM5vATUXTUEjxUE0SY2
7MQjJiWQn8rt0U+fvTqR/YepgzQxFF97yd3u7MIY17WaZqNj/t9pktci0OlGnXW/Zn1SPkS7TXFB
plCFjQkbZD0n1HyXN6M/IJg7rtwCsvdUytX9s5dX32PgkqOdbh6C3YCpumOCDzlYrNlg9YZzp88W
jyWidg9v5OAnWrSMnoRVQOekMBoC7C5kq3qeIkM6Nn/xcyqoSAM48pI7fKmXRfq1/aU6GRckk4Kj
QW6Jmy8a81ePzYuUTs+JcUNB2s/NAV+P0mr13n80uthXksXBFXEqik7sq9ENofIDNw+hXvtT+wi8
IvXAzdfOK10o3ZnVd7wna3PCD1XLv6ruS/hxyAeZAc6ChVBgq2IZ7A0b26pGKKuv0CZbmSoR/bvc
SmzzRfBMTVTaQH0CrPHoIfKCy+885d2dYSKbUsP9qsleSPpj/pc6racLTo08vxdNH9Qs69CZ3X/9
31WZjzahG0fmrU8oC9p/coxtXCB15zcEZNju5vOjWLIrbp8bHSoxabmsz9c+tfKFXaB8KYh5+L0o
YZ5TgK0dA1qnCwroCW4uRTcPDBrj7yVUkls+SG1d3TvXgRWs30okKownND+b5/bIecpV4kZB8A5r
TodclHTRk3bfOSE3mG73FL52a5VKmwhz3rFedGKrGxqy3+HAq44jovRxoH665PBIrGPHiANHHC3k
Ar1g4fRqSho95fyvMEOLapzWyZcd4JDH7MB/RWWcyOXuF340jvZHNKfvvdL7VpB/zP5y0SzCvKEy
CJaw6/PaOvaaSOd5PbpKdMLE7lINHQfLIqsm3Wd+GaA7D5+PGvlAVTn2V8q8WnIMu+5h7Pe8eyk5
2Q/QGoOFyBxaYkjIphDqv9KE3Z0qZ8t5NO/HKEV7GkGgWuKU3GDUIfKMQ2p3I1VrlO0wrUEvJvzI
er/2aOxHo7tU3BJgWHoylOzEjZ4bOjfRV7o2o1fzZvdOCPn/zXKSwsy9ix2ATX8Tz2ogLELHb4a9
S75fBwSwe053QlQuHRRF0u+4iEiNNnUHsZy4jh1tNvZnfXBQPnIrKyWqKHeEPhtF6v9cjwnkRG3s
7TMMIl8VserBSptEW3RIZoEEtGk3CkMLqjSOnwJ6Q/AFb3eOod+Q5chYfUGHQ3/ut0myOFHpet7Q
FugBlW+9n6CuMWQxQANKPavGbyLOclrWKoGSqDMGNaxzQ+tZT1JQaSOsOZvcYMePD2BPC2EVQiEp
JcsalPfvw2r+MvX7XYbbPkQwx2L9XCOFjxEJnz5sqiae06mB9/VeJaJlU1KqCQLbpsJ1j/xPdwFr
Z76uom4HGN1kbs4XAlv68A3CDlcwh3gKdz6yJFn93+peatd/czVl9KBZQeTDMVNaal7XmSNgwGP2
lZdE9n8WsMMj6tNJhvhcCrICAk4LEzPTbjhzF5zRxpbMUB6/jwK8JqfX12bPspiLBhtwOn0ILbQ6
z0pVSp6a5iDiUFyakolFqnBqDKaD80FFC1bcwxJEldtkpY37YLbFZnCmjqpATQElBoLGfzqYSuKe
KxLG+KRJ760kDh4LyYCt2E+B+fnSNbKz+3dWSgXWQmiFRWDd+d9QdQCNmWp7aa4S6HvSolazAx3H
XPhwV/Gn1AemUTKt+bDLA1LxE3Ua3lfIKbR0npE9bjLgWgs5+wk7FyUrZ6vaVgjBb6ZZx7/QDnWR
nreRhxpNY516jEDB4IxFCtitlqT7B6eCYWV3AMu3MzBMJKzwz276kvYs9Co3hcTm098LNb+x8uy6
MIjwgcxsjFEEcPpoCmJ1yesTAAdLYcMC08TlpzRFgJcqI1WgWLPvGh/p4bRjS1Bfs9Q6gbUc/u5M
+fegGZzkH1/ai5HKEg0Mxq5Q0TLgTKhXhJahUbUl1WD9T6Hr+rQCdeVpQqR2gTRbBxOG35vMy03o
M6zyAuwRf0vFNU4ZlYOVZqNpGlctIQnGEGrEN0qqP4ArPysZlU7X2M9rK/KYHZnwCFlGe9mzxjMZ
D/90JlhCKa+f/+dd5DaaUX0SWviBOtmPNPSSPzfQZQori3HW73QpjXRjOTANstvgqTXPWrNujbIS
7MgLkSzBwTRFSBfzDv49HtNRINdSXrROysAD6zdDYOEL4/0L9439TzeaQ/cQlW7P55z6tjG6E4mn
bjUEGXpbqZa59w/bzqFZDrk9Q8mKbmp3UUkTXcqA29zOeJEDABpfcBGiO2rvRgkV37Rsi62eeFkh
yr5oskVb0h8BbG+RSgYhj+CO0dw0en4ZD1cAg0c0LJhQSKSqr6nKYeJg0O/TNpqoR4TOMUCC/tfv
tt2dj3/34BBBEA1/ud/5ogMo7wlc8tu0BATDWqpJThw0ypcQ0Ks5oJo8q0cFUZ98MS14vkDtrg2N
1Ct9SaNWYNCG0RkbAE7EyHvsmwmj8nk/WT+kbL8KrkcrExqe9ZCBHWIh1xdvJcZrdqz6yX86ENDJ
p2XyLcCEPijyZmfgL0pdiP5vNpuZHMzDg/WV+phx82Us+lHK0hUBKeywBGbx+Y+Rh/UKFCdZcXrD
7b/r8ENnReA7OSY1oE9hN+9X6XA4+GB5Z0ldswAOp87YjSuL/wJ7pcQg8hHx52Q3zqas8H7rM3Sl
qISo4zgzQcQw8pETCS7Xlxqs1OWsPT4jfWbQZpQLLiLhD21Mj4kJazhv+PQ7FXsXsmiOk6z7wB0D
8829w0cO+lb+mq1+W1cnNYyXoZtp6hXFza2rmqfbE+CzWbbdY9sr+c0vF0LNOBMJYDBT371nQB+b
8tjGt0X8zdM+L5ttL6432/ZfIWbPYdb+CmcxjH062AKj74W035FueT9RrR+P9O1Com3QcqKhcznR
CTT2WHLCWr8LwBHIrUGVn1r0OjQjydOaujQjLtklphQ/DcQ97WSSJP6LaKwMs4qvS8ZfrFfBUc2O
VLp13uJokUwHxWuREGPP2S8JICAkSg1eu5wlrfq0pkJMhtpCEdm8eEjv76LWe/2z2//+k8CkqG0N
XzaW+u40mlfQTS72o3IslZ4MvP/7wXKhUUQX90mmRTXIGznS3P2SFaqzP+Qxqqhe5yaKmwMFwrfy
jSy9cdXGewOVG9oOBTGmtFnskx8OKN0+hYwG+igwm+avKgD8gKUL58mJoboK24OPo3qxxv8lCsus
DI4a96q6HQUGpmJKPnKZj5gxcir3s1WjvEJZs0T+TK4Af5TXehbRoMi3Q/atfOh2mdUAY2vRmsxC
e47wxcPhX+KzdtEdyDC+3ltyBEfhjmjrmpfH96eTj3oBu7WV+9Njl5Bs8eAKUjBUwzUwadjhLZyk
uvF73vmFRojnEB1JZEFbDedEeyRCx638P52PJtKbPkPz/oAW+qmr1Y0XKGkBWjh8R9AolKs39ObL
jsCnzSEyoIQitup1/QQHXC9mZ4TqSXWSOWc+gW6uWMnKYc2WwuV9LINuz+IswwmOL2Qtw3bX60h3
4jAw9yJbbMjL29tc0oPFkyEUnwKUb+RBGA7hMN5o7L6ACBs7AsG5UuHMtdgnITKNhGvjmJ5bfC4D
poxWIHo/oBEhjLdr3AMzTVHssXHgfHAKcG6kzwqFSQ1GtxgMBt2TtXA7sz31bEnWy/bsC7DFSX9t
N2vej87s2TLFRuwB6/ZKTwrx2YuKSvTI0KwET6Dw75cn5PFOatpTiFXPJSVJuOdNwd0RvHbW/kZU
vM+6y4lNSA/8qT3N7chTRhUtT367JiKkyE21YY9eNy+fe/F9igOOab7AUQMPhzF7WjaD5NfN0B8V
2LS8ef2Sx3eUcnltEfc0h10pysBfhKB7QfSY9uROriRyUAHg4oI9xe47554iI8SwRFYYLNWKTaQs
h/C8gj2ARGGS8Zw5yIQRuc637xg/t5hDqYC76hZcJG+KwjHnG1wyvsiaaDBxUAheW01EQ39ia96s
GHFEpfQb7lHxzq4gShBSFU/2N3UAY/7Oae+Y7QFpwiWafjG8LTlq3HmdDr9eQA925uCu/L28bPx+
heRY1u6tORxpVTvafFlzfwtujFXCWhYlNfprZHsVybnS8l0zX6YqQGEXpcY+Nejn7gK9iqWNtTBj
AgjEfBcHqX2kJS+NGT7ko7sQ10f4pZRnXyHW7byNC5B9YhPAqpRurQCt3XJneyFXOifxhoLLQ1be
QGqP7NHQZUfAkcbUDZJ96cXfrY9xiPPMtO5pw405BwtaBonE0MTbPeLWFVzhlQW6uyhrxMj7fTt/
H7SmxLAedy8W0TeS5CVyxpNvPR+PGBhmjn8iOvi99/Vn+gk52s6FkTrPVCYZ1IJNKFQ57PydcYmk
88UI7zxyyG97vSJ5qH9J4Nc3lHSYeH8Zn3+hGs8oJRKlQB7iLRr9uJEOchiLbl/MHfHfYNAXSuZs
KNN9TPV1c8fpsEt8ypsoZ9yzMo2iIiYKNm14K7p6wyR50iv1n6shp6tu3bFCgw+Wba+AncV7kSzo
Ue3J3MwLB0MiEikv/NRpaX7kb3XJp2/i3w5J+WDXVn2u/QDT4S8VtNI+AtALKmSWn0/IxdDdUPrY
2R+iIfwAGN3oB5nhRG9Vkg0p+dgBrZxczsXS1JqwnVetuxPqD/zFR6CLIeEJW6cKrRYL0SMO/A8z
8O9hR0ngfG75d33vQ28D9vzO0Jf793vbLR2ThTJtdeycmv8fWoMVfveLjuQry1KzL1Npe/U58piG
gDs03mnEn2uSGV591N1E1JQXlW//dkxChHVD2+kI/m8Gz0gbuOe8iOYO2ZW/OhFI7j3mA5KaFQD/
QN5eAaxJag+MzYBYpL0wjm9GWxAdum8j7guqGeJI5fVqVkDWlVO/jSZzuuf0ChCeYBw1tI99+btC
rMfJC0bScCMZiwhodIejZrZH1mEcGwldePwJezwxSr24whrUggcNvWCmflx9/xre66IR1ZeIGnMy
qGyYkCD+lzzyCB7y5thbp14KgeDl+3e5nyyf1aKmAittWT/UHRW/9WQ4+haFDpF4wPVWEChib8pl
5T8f8iGB8ThsomMDPji9qlMA05D9jbC1l/n2z8jWQ98jyY4NOfITFe086DazYJvP1YsUH5QMUHbG
vcVr/28+L/ZUCwk/XehLPBfo6S/WsIgP0xxrM2ugWQN28yTJB1NI2KcwuRfkQSL6twIVXD27CeDt
V+3TCT6sRZkQyqBzvmIgbzVbDL9nAmT3/km2g2QkI6Zyvh424F+HaHXVMwu9R+Fhp8LVI/TJnG1M
0Yj585tnhMAmTW57M9k3wnlszwvEz3do3CdsJNrlkuUjyD6GwQ3SKK2VdFrygQ86snD3I5xin2bv
zRxS+97NirogZHuy4PmdQyLnG/57IoBxS6AXDsjB8d+JnA8vLZ52RHX3aYC1d4Wy9GUAhKXy+qnk
zGCFqcpSUVCaHLgez7XNN1BiWR7cNJVvi+JJfguXimuWV9SDnIXblkCUJcFMyzuqDuba47RmL6xI
SguXPNTtzLUwwr3LjQyV6y5Qfa3HbYllEU+TDSKcWbgY3y6T+4j6XLJR/hoTegwaoHjSRDsXcJO7
57XUxTaMJMYMmsbJcjnIwwtmJpa4zjIKCop9wQH2W+4z5K2NDpVk2YoZ2iNvySaYkN42rLAfXQpV
h75WFr9zeSkkDs8ltpgUmkj0P+iJc6dXDowTzgBViYzArhOTiQyMMcF7sJ4S2Lupd5wOlnOeDK4d
uGmsxb/mEgf+/Z6tajSCr2Op/Z3jOFkOHumk5egBA5bI1T1kc646JZp9cBBkZxEXRwx9KRHG/50G
cWdJ5gGFptGgO5+dJpL87yhkYQjtAQ43cQPt4raj5EzSb2+cLKSrQvpIWM7Qn+vp/rvoxCuvP2s1
4059Z1HV9e+AU25uivBkWn+6Rrmw/pg4J+UfattzHxqGiZIBVbuFt1hxpAdSv54niWYjm4+1265s
1+sAZo1/s+NcFWCuK66qJ0Hz1swdFTCKF4zag4i63O1Uy7t+vS//45QmALc7FtO8XMmBO3WwRnhi
Rd+zdamCyQS49eHvB22ToLz2KgiXaQ+wHPb8w/OC+y1m3SIJJsHrBlwjzmnkG52O/+jbOQl3QVI6
tPJBy91HmaoVf6NTMlRzwcghtnblDXad2vqmNunbW/uiqIrqnrRCM3nrjFXqGcbP+IXd17gwurpv
eXr9xhT8XsA0ugRpIl1wTMo0cCuP5cWHlE3i6pkeRfv1qp0Lz4pyxoD8sLk57OHCq4mvM7DIOv/M
/6gvb9euwwJMrZVXlWPFCcmratxXuuFjLgaZaq1AxtfgatqPbQn2/JFBqbMla7aT9vwxVywFIZ0w
793ByYAGuWawGYFKBcUBWqr7dJYzxSWT9oifhZBrZEBZMX753Jf8FeUHGtI2mc6oE9cWKKVquzCw
bJR9Wjxk5QdwCNNiAr803+tEz+btmDWDk/m/nSQGkHe6j5aNkSWaPHxV/cwK9p3c/ySwGw3MDYsP
quTMBoCeQ2SLCGpDXa/KaV7GhuWBw7izDZtPKClDdUSZQY4f8l4KxP+9kmnfk7zzZv98eGigdaQA
xAKK8GRf0lsY1sDyMh2x0ctC3/jvIFWmAvNzLiWnxc/ERPo6wNYRIdiaboTh2QiGydYP7LMANqIq
lZdxY41zCiND1Iuk0GEUuk9qpNLtSi54D6Op+IIjNbmqry3C4r/dmovPkT4zlvmF6xFUtsGidwxF
S7KqBKrUsG7z979oyqaQzvj74Zz5xx+v8cfGp/q0A8qoMRUpzgOrHKUzBbvIOPQwlDELKtlUIIJ8
is2JpJ7FXld3Coz6S2cXuG4Mr+jugut0pik3G6MwVTxjHrC1GG813VwYCbvv2YzWR8d4IA4s1g4/
IRC4jQ4m0e23VFamHIegyqCEM+AtW+OdydNFCypF4v2owUqP+muY6vPNQw+ae9nRZgv43aTeqLqo
F5Ay48xdcoYie0fp4/X3zscd1ACNuEbg/isXsiSSAzDbmKkb5X+Vklk9RPvqqCp6hECx66aUwzww
ZuDrR1Wp61Oz9hyeWAfGfl971ldo1+/DiOskMrgpdcKPX3cohnguzgyWc98UqVE1bGyszrMTF3Eb
HxDhFdTDfo1ZnrPqyEqcf/MStfjp7Ao0bXtREVYcHhBLOOjwzsDv84dCuyp0V1FRirg7XqeUp8xD
wBcP0ojjPM0QIY01sHffYsOob1oW/S6JRqgTFk5o6yS+aSuvMNwDY4tS95lPJ/4YEZf+CUHnZVCq
oHZ00/7KJG5+EAGxdDEyPGyEixx9FIz/NJ2HTs52tudyNQYn0UUV5dUhQnPfccFgSV1qjr4k/+bl
Ug7vIz0UCmDBSRql2idbplfuVYcVqdc6cF4XqSeSKSirMQaq2B068P0JW3MHj5xyaY4zmfgwaF2h
a8viJ6pOk8y2CMgavknqw94gy2d57Ah+eqqxpBg/1ZOwOJTFChrW3uzodeydL95nfpYfU8r+bEQr
Qx3Vul/tvPSve4hPXbQiVPoFS1FQb43gGlLR439vU7558n6j9p6sORjUcsm2/PmnfijsqS1X0BbF
G2Ez0m/VVuHrfnCFrcWPbc2d1jvGHiI67fvjYbVvxeLQdz7WL7biiNOX5CXfMMlsZMQXdmIjKsMQ
9Dm5MJ5L0CizBzBsryD9ZF8qrWz9z+lgA7Fumw6Nqg2R2fG18F7CmkFGcjNuPRP61REgQDdpLTgb
P/2dODr2g/YIZEFcKj6MXKmp9jsVde05Pgy0xeBViYsFBmuo4KfKJAyZYLZK/9d/SglNk585MdLo
D8vrW2UITum92Src7xS93azJnqEpBI5fsOtQgwoqrEDksEoP6MraSnYrZNbW5F7OIz5rv6oOSJZs
B2UkZO5jY+wJVszIhOyC4Hz0AAQCT4Ga6h6n4TCxW07sokU8nskKUZXtx15iC500G2XS2ByMGF0F
dfDDzxDHSzwJUfx2arBdp6rBxaIh58qgcAsVgNMwHIJsygaPSoeNLK8Gz8cK3K15wZcYrSXYUv5s
zsb9xMHiPmdnCAxkX7ULb9Csn4smnCVLe5i1GrniNb4bDhoHJXHa9R2wNE41KE/Uhgd68Enm6IrL
VZ0N/iPXpEiY18E+EUc44Tm/Ks4gUk81lED3tvToympxJvxfLuW0OXVT6rWLFTW4EvW79zzBmoZM
UdUe2rA+f/uTjcJKrCDszcqy0EjRIsffWVJTsa/IjOnshVEDUH/W3btS5Or6YC78zOR+p48IczLH
mmaMs0V68fKJ0RkEW3WDDGd+kbk7hzn0Dmp+64ba5xeVBqU6LfrMPOo4LSGncRqryNxSWln2Daww
vSenhxDxSgppBaiYLn7m5O76FZsyjzWyhQRZsKOzj0YlPxz+Ca2RcxwydbuQL2GQyPrgHOp/Gv8r
mvuvcGT5b7muxz6xxzwht4YPq9PnYbOzDhkU9/mfGzjR/DHA3TZZxq3BamEttWdosv5w3qyKN+b3
BAwmOjhX3p/w7m6JayfCGXdl1GlUNSXGqufZqK+FOUD3Llnkhb7b+pLjbiPm4Iidr2oSBP6/jN6O
1bdZEgPqVaihoFCbXyxrvm7aHTlim4QLp54RL1XFRaSdPch+2fxC+/sdazVRy1GjElPBZxHe9Isz
IG99CkkuevViEJCRkLFnRFztl8wFeEqSkUfbMRFK1P4wAMWml59po7okN5QhWJ+p9phEuwbv5O9A
CyLD4CaNVYeLKHtkrMwT6oGA4yo9Eo58grHYMLQO9vpAwujSycsiAr6UCFxUsuH0oHrAt3JifbQK
OV4q23hx27dxATk8UTL9qbRxu9zomtnRmhd4tia0GeNTbv+OX3GIzIui/5lMB8aMsKSN7XCVif6Y
uGCPF3fCuPvAld8KZxokX3e6Ls0n1ac0X8bKke6tZWiyMBh+kVoEv4xha4nFAe8DdFz7S0XA1ZwZ
BAWRfau3l0yX/SOMDbIX9CS+1mDwWXm6tEQgwBUt2xhjM5NZq640GznOeYh6ahRiAcBLQfRzyGTB
bsvafAZzArKkiYXJ/XfuIkk4NPkrUhbFjcmMhLzvpVCtm5yr3vcVQfx0ChfIPtLfxbthjDJTRndG
2GjWn0AHxghjk5x8/wWw59idtdxJp53adm7E2XDFXfGjx137U5wOVD6fDqdzQFeTJhh1TUgp0SCb
rZA21cRyvG3ntBK1rx8TNCSCN2P+YoZXGQbwL9vuA/M2x3B9P4gFNTuTRJquBPwqCeIWgfwNsTFw
ITdHeUn9s/bbelfuflI/l09rEqhdieFzRaUeZMcdOEe0aQHJE2oev4+DChKHHQRxHt04I0lciwAQ
wC9VRB5FQkq4UXqaEZJojy1HnKWwMhMAa1Nz1qk/xNTmdFlp06vMA3H+YAYMjgx/sdSzg+1+2jGg
3uE1jg7a4IdTMphaXf4LhEFexqQCCcy5sPp/BTBvKV7iTOmu9FTD9VoRf2VkLbV1/p+aoFyZoMtF
Pd0IvYx0K7PHzSgaZvseVh5+8oLRvixLgAQ0jzZXu2RFfUGOKD0QNeiX6ZwTsTK6O7/HnLLmrXq6
cyTSxQ9zfup6URgZmtgQbwdq7X/ZosBZwKARYWzGG/FbGFyfTAfSLhuv1IMWDTQRqKsOhrYnnCJW
tThhI/ARfRp8tobslH6iVsUYHjmiXVE8men4Y5N9saueH1HNBIaB8Ce2muLoNqz7dA3a2V9Ju2s0
8kJ7ULkuOLMoJgxdTAGm+vf8hMMWOo8pnkbpC0jKYUJywN+uqBeFdY6SgizgNi/APeS5MIwvdvm5
G27zH+mfyucb5SH0nVn1/pcmFiphFFrCrLYKPcuRXSG25G247aq0IThOoYFWkLwCVWoDK/D4okWv
zgjFpC6kzBfY0KamMfYSUT6exYNfTlRWsmnAIWRkVD2gVdnIXjW80sKR7Zcy0J1PjU4kd41tlTrN
qHkjR2mL9YUmB6iVfaPX+gBhGmZ2IGZNMaqNtUE6XRgS2HmPjk7D2McClBpWlcbihDg4sYznpZwt
cnl00y/6lNjN1mj2FpFZkwcmDrqidt05WDiTwltXnJdfkMiYQnKeOiFVLwZFD68s23gKJDQkiXHg
PcF/KIuTHqJSv1AxH33q1mI41KSdnTfSXNOjlJjDUPNgb/mGVdXeI0LjNeqYzaTE99s1qTZOtDFN
arSOlqUDjixfunYlzWp9YuX9WK3rNkhsPfh5g7sIFr/DENTci4cNuc9HMsTDZE7hIAHKYmksYmfm
h3hdWDgAtRWAqwL9rXtMLYwxh3C7+EqN0nWNfW3GxhBxOt/inql2bS6HdRjPsa0ovJc5Y2Cutp5h
ObDOEGj0qUw35vS7jIfV+6/myaO8Y0rQtONcwr30RWMGq2cobsRWEdTAKF8y9TnA3wNCNoVkLhyR
vLc0YJCvMy86nHo3+/dCHLo5wqN7Z/R25a7pdtT3qzkJh/BdwlEpUO6LegPgWsuq88/0q4I6+fyl
O79qryzpP951T8vHKf0d/e37jX+Xs5NTlUrnW4iHdgRag9X0DzOWvqAedxxfZo2s6Qo4xGzcfMZl
haMPLfnROs+t9hvdSnbDK5IjsYUElRqv2pBM47ngQls0kgGNFMy9LOXJtAHkd2c48lQC6bAY3jsA
mcX6UmU7MVvccGXACP5S1iI4ZNcdd4s6H/Q1PjZ9JMwHzdLFWMI2TJ8dUvjTu2DcxWX4DG8j3JhQ
AVP39et12/9B0wgMxPyVPHR3+jiRuISBiNRWxDgQMStzVjtGWaIBP/iuGZ/M3IR5M0bqjbz0FoU7
eU6Agtj6YVDsUkZqmrvUdLGk/4xucgCLECVDg1GLuWKrslMeULD8PvimOGhFK+rx+vhqXcwNG0yA
eMR4sjjcJIQz6BEn8AqmoHPhnS6kLkeh6GsCv4hrwlkNtjkpWRRgQd/Y3NcfT51YDEeDFSUPp3xu
dQvMlk//OBcs3XtpamEEFS0H89EVlsTjkPjC6tTW6gJP5QsjG365F1BosKYHD7iT+mszWCgSah+A
vu7F+mLEQFGlKT72AtSIJFM5/9YeJzoBb2gDnK33FArcREm9PZ1AUUQZB2QlCAjsRvd08iRLe8J4
BQJ1Vskr2EqS4pBfVGQeDM9nf+vczFOYOzVPRCvo4ddqIpcMXatt6ej9CHjKUUUuSjIixx8Y0hiX
ghADykGCeRcLfDQrJQR1lJd6NaRMcSKBx5qJ63PFUVX9HuUQ3yWFaW8Cb+3S++VuT6kNjZhWcWtC
ZP0j98W6jcMgbwf83OiWAD9cGukU4iOS4N3e1b7WMnLDKx0cTghNoTlslP0St1lWxsef8YYHXyHM
iwL9p4/L5qLQzSy0tehLDaYaUm3Eq8C4HFGw3GSl1zligcA5r0iZDxd8frRpcQeKEKtAj80UBHLS
CaALXh8oLIQp+bws7VutT18OOXoBOu4nigeDYCzwtswq1sn+49lM9rt2h/N38Oi4lWYTqU9AKP3R
4B7fItneXl9H77KhZYldOvRIXiYLNBZrRlygsC3BXnyfCfaylFioC36Txgw96RR/9wmWyMLwDpnL
puZwijFZpYZAzKYWEn5NdYYm9dcRtawaZ5VdRSZnY6utxJGAdLSHyJoh6rj3xtjkunE+eoYS6Y4Q
26/xCYpJoCj94Zs9++qPGvZtfCxyDarVBxGmBFGLlcXEknqCWVMKBg0XCbkijI37+Ska76EeSPIw
bEAY5yYNpRHY+1q8dkKRkGSX/6r8w2+L8dEErF5JDYYz+diWMXP68IL9eQkbAvGdAOzuIQOHyk2J
W3xvI4BcCyQRV2hTCGlrGcxK71+WtIXd+lWUqZSg3aGSTsm6nH9CsVMuIKjmYZxONDss4lkzUUTr
cIVSuyEt0weyL5p9vb7sPh4yBvPXlPWM/H0MAtwKqH8PcAbizIlaKfrvHr3y+XU7XBwfic35p2Hs
m01vlnAbfQBFU4e0mMB0ZZVpjwzV3ivpgwWrobTiwUnmqCoD8DzpuUQgI8AEvn82uOBA7hyp/ank
DzssH0QoXchd6fJt9ykR9fQ/5aeoI3QINYhguEMKvCCve7zkEgzxFc1JiBgK2//rMnGyGWBsVisx
e8aVJGk69yES80dMp1XVOIhPlh7QJ/uRvjThJhslMO0XbYVQE/VRskhYPZL5m6tQci8+yow/+Ws/
MmDTYJKIR1gHed67TmDdoitsN7TJaMjPvFobViXLQQ2QzrzO9BpXYBFZeY8PfCyrhPYDr+54WD82
9UhMebpN5BbIwlFxBIYCYY6MVp2ci5EDrObM5U2+ohnQcROvSUlGWI0j6DPjMK8MkVGNo5ALG9Y9
FSBT4i+7oAqJMAabFg+9Z1uyLOSjcrxcN8GF3glToC1hmGFEJGcRCa1SZXOpXlluXQeCFeWTJhLP
QC+FUAlLEUlOYqn2pHe2E4IasX4z2J3HfQlrb+RSgpLSC3RtiY/lZ9NL6Ns4OfbwhTi4aZZ191CP
8jzvHDXctHRrOv0TsiZcw+M0m7jQOli3iGBIQBYSigZe/TqIMcCvfP8whA+mb8pVOInctFgATydL
Bmzz1xgl6I7vqoy3WGK2ChiTkMmkOOXw3OcaqwaahcZoHL/wTWGRbjeg0cKDjmQrkQGr+3ssb3oH
R6cwOPp3zvvraGkPVyRK8b/wdDONT97H8YvUWUyqSpcoQ6c+NknOpz257YvnGfE0EkfvUWu2pMdu
a5J1q7TCsZNdqf21UjALy4dBRDB0PqaaVPYfYQrwiVYfneHoYeaFdTBg7OCQaySBVYnUb67BOgt+
VvprvZV8wQVTirpb+EC4wd8leinyy2rT6SJy4LO3CrQbQkNLwRYQgkdT9AQNcT6m7m3wxN4anVMG
IlbG+hPoFIzpUnmWRwN5VoL5Q5RiGNJhxu90wWKk/3smM+VX6/iWRTWF4hXztCfM62RPz+uGC3y6
eCRkL8v0Diz1yAIu894AvQtVXLD+lh3V+0hi6m9Bj4BIrgpcpx/zaWCqbx9H02YCjlQ3Tbztc4P9
Z5fxwSgs3ZBTxp5jld6VK5OOEkKRHWIi5yMHNkHA99s45lsJrkzh96YEZiJUZHR8NFxSP+hgxSgq
eZ/Ppoa3LTb9GfeKSVn4yWzo7W3Pexnl+OhUKFiqqRjqHfHpX6RFlNMwHE1Z5CgnVwZNDZSp8CtI
Y0bj6s313Vm0xn61znJQGee1Vp7Y2hMl7ZTzyOFVPbAyHBvQw2HNBLJL5EJ/PAXkBxkaGtDbCE7X
bprfSvz79+HxGHdKcKPE0u76N6fJhR1hloN+tuu0e549dxYxOV+5h3mfusOOd9DR9ZJt5fq0zFV9
hAvxf2eY73YJhIQMRkHi2n90ADSTfNj98XLQ+9psRV0zJnHFGkz4Xt6F82ccIxNx8fQLy7JfO62G
X081uVr+qQK4dzfn9fZYigCv9Z1+7ptiklsRw6WGZkkbmMAAZn/mih253kS2qTX2JnV6chSkF0na
C4GL6enBudvaYUAa6tjaz3ClOgh1b16KRQZ9m3i3H7UezuqLyhnBb0ortfSmnVc6d9Th4gUeqbhF
05Zj9Srtx/RjxuujSG4Itf3PNqQ3lH1oNgDhh0usDREF0lWtPOj7e46BKquBK1aovbbnrCrDESNJ
2vacp9cu4gdcFVqqYAin6eZcQi2AO299Ql/9Wd5WTpJyegytk4ljCButpNqAOwAN1BxfZ/1Z2tyI
iCmjoumTNZcS9l8ZKViewbQdyE5RaTJDgCMgIpWkypRs/PaqJ9kkBCeXfhlQK5SMRXw4AjkI6Ld+
lHArf1FRSuSfXJ3WVeiWpvpecDJ6AIe2OeXMcTtFQlv/Zt8L2MqIqCyMPjgtw9Mcc3spmQVAZhGK
BY58IVnDD5rlbu98RrFPdCNLJ14gR0XV6ETiwOC2ulBrB1kyyLcOspnpjOc6i9gJ2qsgmsFyVJWf
9tSmjsMAafOHrj+nF9CnpOvF5wiyWCxW1g1uefMZV5tolz8GxLw2VC8kxbtjWl1oyyQkUuJl2wpD
Tu+bu6eci8BY6V8AIRb2wLyFkdjPXSkrNEC8MwbfU+gzJ7172DAjN/UVbwSKr0AhakkxGUC5KdmE
YoBOOguMcKFXSPkr8xgHnhymyXWjeWNCDEyP3aZ/H+9EPsfVYcbtJpQcylnB7jC212UWQc7+ey0P
8FanaF0UdmKureq2HmEWzGwUUDPq1PxJaOI/twRHGntIkX5QKFMyhZs9ACkoD97JnXku10k1zj71
Ixjn3YMjwHxUS8r7JDrBd3vfc/Mlz5dxq/hyiPru63YGYeDhhq+X/SuqO91P1GjNQc91cNrNmPap
Om9brQoHTehOs+yWy43XY4BX6eYHGbukEcnMo0fNDJEHb1xSD9tW1M2KnUfErP2JDDohVCbfYPbe
kEmKkH9yiGcEWKBGV/L+eqS75VTLd3YK2RDgtNjXI/6a62yiA84I2v2qmhoLpqAaxbruj5ahQsh/
SlmTmZ3VjT/8OnsQh2caDwEVPoIsXg0Dp95OdUbuBHzo5fxio4bY5wLy9sh9V7y7o9D6Gq0HdmeP
mBmCRG1UWUsC4AVh8mprpsuYssKw4PaD2Hl2gWK0X+4gYZ6XlkRny16D+fk946I13P0uIZph5SvB
hxh5+DYLaILbqBGR82uykNaqDwGldzbUrclmK4vbinEC9PV32WOLYEky+tkm9Z0aT5bLY6QVo8Uu
IeGVSATnye31Q935AWO+t2q5QbrJiPFbMdvyjehXAfWms4YgPHinEev2zUB5gsE6UZTTSSxgq21A
WdxOIcp/7xh6VgMyTpb15SWP29dJqHwQLf3XcD2Q+qQo/7+maZr+OkbWGfUd4ov8EwkRmOVjJIpw
ea5F6tt9SU6wbn0jxGX4EKFmRyxUITV12irCsM7I9SkdOrfU79wEBhEhkCUg8110a840/y2My/o4
O+zWTU1Sp2eO4fxYkKGkEicpxFy7uS183C2oMb3k4+j8t0xb37n/xtehpwhRFknWqWVCk8Ltypcq
dgeOD1vJvj6FNrG7x4M4/RjzdfbTZBWDobMxY5wdcvJkcijz+OusWCeIdpLRvpY8NBP2rF36mQzp
oq7I4QrYFdpu4izurTbLnw8mJPMCenIDxhL/WhmxqtbMSGyr7nD4BYTtEBn3g4f/3EyEX2wzqBXI
JBvwogNbZj+SeFiJENGWDysQukh11hRvH2y4y2qhY80MQG+fHSWLX4DDOxQzfqu7uIm2Tg3CXokL
ojnTyXH8yiOzQ644TtDauzBoT/0a1j5fXrfBksXB58ft75YTC8wA0FvyxloZy2S37kc6U9+UHCyQ
amQsALdyswTlwJ/ZJwWgQgjV0wvuFG7Pf7/fLqdAxncocFD3GRtRD30J3d0BQGA5utLmU3FHkCvb
NJF9Af6PcmqQ2ioFtFffRsoPdofMqP6hN68D5kMKupZ3sktEgXS4K115dth1QnV7hBzOKscx6zq8
04xOOCcS6mjX4Prch54C/2m5g1Ql6fHSJ4LiNu94p7z/kOM+8tou4QhX4wJPhcGZoLQEOJATwFpo
uDWtLKwQlpz7mjxzYpZIjX55jO1c/zNWC9408sW1D0DomTOBWTsc21c0KzghJKnhHsFQLbOim+vn
ahcEQ4qcBpjq/afjcwTVE37wIDA/FxQ2l430jNpVLCoeTFENdfDC2cgRoWKh2rlX6FuBWiqIt9LQ
sXWgAsu/5yjYUHYz851zQS/xWwacu6F8EUGFxkpIK8/mSrvzDqvNN3DpgUNLGnHgWsT4mT21tWm1
rJ4Zdrwh11QjnWRbllZfdPaJoG0Hhd/iW3roKJQYqzPStlJlwm/HFF9KKI5kkdSo8QbOCtOWjpvA
cIdJ5PrRwVAkbf32ljVyp2B8+5lUclQVVIlTR6aZhhS5P5c1F7Z6rdiA38gLnOvc2WToCGpoY9xV
vwA6YwfOeQeFup3ym8ThRHon9euX90Xnv/4g9s+V2Dg3FQJYE+bxmDO2ySWQa0s6q8QawkSfBM2o
/6C0yzKZjOn4ll/lmef7oD6cLIlo8VjqUsMmv+t53uy7nxnIEe7p+ZDS+xJld/Q8IyQ0Vn//GOYp
0oUL6zZfheLVCT4wzL22GgDItgTgYZavnUjUbNUdOr6ys6h00DCG50rfat9MjjsanwaMewKQEGdt
r2UTeEqPTIBAh6WXQ3bNumN7mSCHeBPKol1g8VpaJr57pvLUy3RZ0UX41Ufyxlb1i74QKJ1MxiLU
8iLKDZ+8xjJcGyUHhPgz5+D+weeriygF9qh6HPC15whMqsNkFFl5VywgVKelMQJOJFtpnq/mgF66
z+4N6hU/Rpa7z47teS/tLRNG7tcB0G56hX6vhUHVwERW59Wx53M5ZR3KqcUrpjJdBYV8Vb6BOw9N
iVdCfbSrXbswM27tQdIhd9wl0IsijboUCerH0DaTtaiQQg5dP3+/vFHgYikzRErWSL9z3BaBiPAb
EbpN7R2q3/nBSXmb2rJhqxATNY+Jypvir4PJa7PsQRbTqNxtNXotetF/OSER7QSULlfwWnnOgr/f
cUlDgt3uMhCKmA0PV3kHc9TkICKz2sJlAj+8hz7w5YxJEc7vS3hyGDjULWojkfty2GU3FIYq5YiP
6ykYtQUqYG4f6mEdqrWFQ82Xrif/p2gRUblAa/HRa8MaMbKXozAtfN5Ou/0WFXukWeNOfsdT+VMM
SQCjcHAS4SdneQ3Dmo8JJC/Avg1g6qaBrPWeWXnec4UbwFo+dCtoHrsobZuBEj9ZbJWLLzED4vFh
EEAzYHMvnIZ2plfSDXT5zZJZEt2vqVb2aMWl+2WC2gOtBXfhX0IFAxPrk1ci5AQDfuLVjhJ1FKMM
EkBEsFMqSYLoFBwhcmghwrVVYhf4Lx91M6VAA2R+IGgCvn0rr1AoLxI8DMK0yO+jNznZBmsvGFGr
867QWov+zQ1ReOj6eVp/Cd8Gw6H7nFAp2Ij3s0zNSrXO9J70Eq6gakkesl+wQf/eof1+858WoqcB
AaO2A6l+fff6dMbbzcxLP4XmcynxknVrlezUXSWwETtjc1JTl+wCxKmusFb94Cmy1jVbI4nZUcAM
0nyHyWDRRK47NGrZrM7SVxgRZoK6AgFe9Sj+FWpg1rO9ien8MMkqJn3p1OdNwZ7aeyehAnvaEf0u
GNXDt8rOKkQUt5zTv3E/DrsioK20DfFDKe8Kk1Z51bTGkLez5p+jQ7rwoVQmKB7oXdiBwPkWj0CP
5YOnEgjONcMTXlXVjPI0i21lyC/ky6Cpsb7DAen/94EoVQ/GY7LVCUlY1CxAqwUClK21mQKPzk5F
BsTDvDKOobz5FO2eaQqZl3DifM1TK6tnFsxQz6f57IR0jWuTXuO4R//pP3H5uAnIkR9LCugC6PM8
9eZGlUXQ5kkFC6o68/nnfe3//hLr3uFrE/jXp6vSV7FfSwW1oycNJyDBrpRW+b2OwziB9u85X13H
O2DKwlgj9ev9RLWz0h3I+HxXMfZ8OgPAwSwaGvUv7FI0ssqA4EvlCIDxAz2F6kqZ4AKIIT7n6j3+
fBYftFDcAvcEg9jPVoCFbm6STHEzA8iAXJFhCVu0PkagaPoLSsjD8B39vJKBCGLnKw5i2ja3UExJ
UjZ5AR+CSLopdDWbIVWAfgAzRvUklQNWHZSiNjc5BUqRPxVjeCx7cEoDP5+Jy+nzTyLadR5Jmk9F
5zfFcVRNRNfSCmxrZhaRfLS1MYQgHJlrA07atKHvRGz4Jc8YNXOYLyI7pO1b/ba+icGgUUcSSBnT
5FzECgEoxhrcZ3RqUqYbLl3tCVuJ10iQzl/iO1DlBBpTK3boQJUG/JeTyE3jbM40vtjJmiQNPRq6
EIVlFz6EQLlWexSC2QDq9IazxK+oDEUKe8LAnS2lXK8L3ngkqcQg39PKDuF3zFh+2XvYB1XhPqHI
UiSZYgon27VES0SDa9PcWpkRPhIcys2f3+ekyN6nltTUQW4dSznYaQOE7WbfRIWHi1rc5UMD1Fdo
QinWFBO4GzS/mgt2DAfrvPDYeBHdMUhWJAURY+nFGG57sRzUPY6XxTYK4etWaNgUwZzZM5WQKcaF
qzsDQtlugzUk+f+ss/qpMtuizxLgbAIcxDxrNklLrd9l1l/VBuZtW8rHtXDZN1Kvp8vYR7sakfXV
4t25ktVUtX1XcrTGppisz7DADrKjQFM9MPjuFpnqoXEperDpxR+zSx4cohmu7F++SMUr53SRMJmQ
BenI8VfyFYT5cyqDVFBlsL6BR94Mb8av7F/nCHjYB2rONm7nNAK/oESv4XM5jzosWTdKuUPIsmAI
zGdSiOHJwEXOCLCsEitmbGx8AgPn7qgGQ0VrucpVUl5fJ9XHRGQTc1Z8ID/b9KylR2AtKZs28cnv
wWmRA1C7tVCM6XmAui4RaczM1cra33HVEA1kPNsz6Lt/cZmAFaOebDYLMSZFFsqAxSQ4vFqAJDQd
nMQdpSfLEnlqN/2/KAWPHxYaFIsFY+Sd4Wdqlt3FB9QIkaKlCKcenlwWHqua3Gsus0GCqARvc2/h
6cQRFjymtCB5xWb4GA60/YUKt1oLqKWbpqOFJ7NIAw1RPcV8e6nc8bqxcEIJKN3YH3wd1QbfL5ll
JbwKV16rujruy8wgzR5gXNr7t3dZZ0I+hbDdkJXV7PGVD7gdI0tc3rwJQo+6uFcjD9Pr1p6Xl5+K
c41ufSNj8h227xVLDoEFfAnpLSRxw+K7gcMLwLYQKN3QYGCzs1OtyzLA+ksqjOyHkf5Ru5b/pdWa
6wkW8CJUCQUx2jksTzFL2m4D4KbxKNqm7otWPqf+L+MkKXJP6RoD+7icRM92fw8QrLb8jfAZIY6+
GIcPR4cqstPNsnNAcQXgfsJz5du3aRWNsaQM+rFTdUmnJaBIrZfkHyZrL3uIJAh2nU2D3ulfLA4V
80snPIA6qfvrDm5q+ukDLL+8Ghfj4toJKSMrWEk7d9cJ5LtEvFQfa+NJ0d5b8KgwRa15IcA37rHq
mAyGu5F61QAkQpBxZsSIJVba1rGc8uzyGSlOcuocmo+dejLftekrZlpygD4JtLqYPfKfQmt3gGQS
UNqwEro3jZ4a+edZpk1uyizhsVceKD8rW73X0SxZ/9SfXI+Lt4YT7xIe+4lzXzD3c8PLwxD/Rfjn
IPD7/ERzLluCqciDrdkWuDon/ZUbywJozsvCEIins/Gj27iy9CYmluGUaPxLyXhj4Z5jpNThGa6Z
h0uLlY6g82CF1H5tFW/ID6ueQg/o7Plk9GY8EiLGJYzRvUx/TlUmALxEnVKY3JGBQBTQ6pn+1CJU
Kl0ckTHV7pYVS/yjZYhr+DHtOW2LfhEoHpS1AZFyQgxAF6vgFAhrI5YqajUR8686IIhVSKEJIzqD
G80GNyMyagQoPqMwdw8Ol6QuZVanbC7ENV9AqYATMvk5/+hs6McWTq0SiRbelSmj2eanaHtB4Sqh
u1WLPtbCwU8M4HQiq0Dt1XK0enZM2i8gLIKPZgsKPyh9PUmvO7u2nYGkyBpeqx7KNdfijANt7B4c
IYr1gMXrAfX4UtzBUxyWglskKrry96aHccnUHdpQsu9FJ8UC/ZpZHOHeWHvqjftNtZlRth/2/HNH
RG2U2oGTUAD9zCZ2uewS7E4yVCczrJl1I/mPz6MGB7FbL6mCTssY1/IfBVx4vXUzK26/pHstVTp/
m5KXQiKNfckN+QaF8gTfPpg1FErbb1zzBUFqP8irgM51JS/fUL03Vz+K88n5HMqeGaxdHbv+0aQo
OH68pV3A3iwd554sWOppqdEhu7n/wOlVj7zOLvCPoYM4Z/DJvAPpxDQLDpPdo4n0SbZ2i0Iv6ahJ
/OuL23mbvbqDacFpOazIFW/8tHqLPHtzo1+Sbwl7Qx5KmAt1TJQqpZOzMx+12trACCNRSpC+SrKA
/RqaucghSyk1C89Zu0m2saR6gAtjO+nWnGMhFRXRL7+auH77bjVfh2U7GUsz9KX8/1O8ZxteDqRC
XMB+sGxRQoJMy6jr8VZw6V9NTTlFw/F1Ipn/jlTTwYr+FhkE5Qiw66YoS6yu0QnpIZPeYBVM1Pnn
L4pZMLGekQWDMB60MwDjMHNW83PatATFE7aDOvN7uYPkFt+51OZKiG+EjJhe9eUZoXXFQwv1kxwi
jx7gGax46UQsIj24fz7uAlW45gV4nwz+orlfm/DFqve2PB6H4/XIPy+C689g8f9WWeNFAot51j2s
WKbIEQLhLEqgh3/SkfX7at0j2Lzxv3Go66YzdlK95968hee0UIZtrv+mA09C0NG2evrhI1ZFui6L
aGBgwuamSdihNf1u2Xb80UwyDJoXWnEycKPws+Y9qmev1dcoWVjdMz4hmVpWwTC7zMd/1gGOKGPt
TjyvrXiWfrM6P7YddnZ/FjJbgtF1MYFN7UyGaM+CSOl/WAtkQCoEI0dGN6w7EcfsdzJwEvIMGI5M
Cntjeym1D5yMXKcQa8P3Ra7Ugv4i3c9B6BwajoxUr7yy+FiPkeTMglxzAXTgPGzK+VprpxkC/Zc+
dCgNBak+3HYwk+SupxrukxmY/C0KAgXphtEoett5/iVHm3qhFkNLT22TsXZnMIv0ac354Z5JDUWV
RV6aoNtCIaHNwFCIBvtJPlL736m1a72KrA4JbvfLlObd4xJadiklULC8U8BCIp1JZBFNqzt8aLH5
j0iGxRM3MEJYfTVvqPkb3Q/LTey4pQ/R/wJRzeogP5wC8FH+g35+Mo/PsjA781PcGZi/JHrOG5bb
EmfXos9MgwHXncs4NWWEYGn85EUJu1GInDGAHEeDxJYYXxGmag4XgOQ+AaCSHvKnOSF5mk7yKn8E
mJyp4Nr6zFmuEmSY/njWLWXFmbBj3HY7WwZoXEbiR1d56Hs1daXphfyiUfkf7mR8cLK1dmwhzYHw
XiHEwGxKOItjhxXFTGXxdL1FsZmb/SP4FfeJ1U754pSg/IfBIuhNckZ0Zw3QhQ2h1c4Pgf/B0j/R
IFW+69LyMW1F3rAYO9mIa5wPYDxoeCAjreJDcGPwPHbT03/dRVEJeFKymJVzUvp+oGd3TOwkmUM9
CMhugbxfkSvX0OpHPjnap2tgzBACYU4rbtLDaQ3H9wmWzleBIaJlgxKFYHQsojuhIRVgMwkUs34l
ylXVJ5hLXmYTCUxixp7/D14bCqpJS5xIW+7Bj9JOIGd/VH5FIfp/YXxpySw1IiNynPSHZpezjEwj
hIgI73emq1p7Dl3C0YJrq4k+lVsIFfE90eez4fJ6LCLKv+QUrGnGQhZ73zP/do+GjZibNNZsCSF9
Rh0F8iP2QLkxH8gJxuKbnByH+dU+kgJZpK23GsrZKHHoxF/2iZBvW+caiTSTJO2L31VFQFq4hJLA
a562aJNzYe+8HqO1bzwzAk16JhgGrSINSoI84fzz7eVtbw/7rc+kRboOO8vov5mo+yGuZusbcsrr
yVQ+gjYRGHqd6oh2CXSjqnWk5NWiY0DRdsFyXujUcI1O4pNXpIXnTVZ1jwG150qOv6yZDdTByept
LoTt69AjpdwyD5TPh62DLMC9m32wlz/yBwlh6MzMpaVzLAf0YCaH5X9OnGjY7y/eVV3+07UDqGU8
vGZKXwksf127KRQURJGgHukAphOffa8UmxU8YWcFfppDmbJFExTptAHjngABwq9ZRZ3Jf/mE+Uuj
AF96e0f9eBhIR9Ru7K0L+bMV8icU0ZtNzLzEZiKsbV7/fqCBl2Jn4x5jCMnsadobAbXPtyE41bvj
p5oWLGcE2uzyyTGfzqZNOlsO0+UEcPofMmcUVae38mdOwKRhfr9phpLJKYWXpoaO7edq0DoWKF9X
7K4Udie3Woqlo9XP58YUTRj9sWpaS6mxyz1SZDNWcinJWsxeSNElEgmNk+OzlfuhXSMLTNAElbl2
zecHMCiMikKiXBs57ngF1DNmRyIB/6cOod/l7buxcOTiK6xXRVbQj0iMm3ZLR7MjnLHsoho42ImW
g0ECykQl9Ukn+4wS9vkyLGVSPYk8iscKMQ3QIUGWJEjcQzq7TtlW0tLM/IRXEX3zfX34QD+F1vzI
s1B8ykzKHRwssPj3bKbob6dwz8o+agfU5W2CzwgQv7jONqDBRm0XTc6hbawukuLvtvFxypfbDcAZ
iahZgqRWcUEARJcK4ALKF15bwSRdZ4QQDFRzyWj+4v0PTb9ASpHa0pZvkuCEh154e7TS9/F6hYJO
Vqarku6veXjo95HPQeUEFALLypUsLNe6HiBR6IZnkasfpJXsKYXmsiFIqswh+NkPcLB+jZUDx8NY
jeogTXAH6m8ercFkP8zpHnd3a7IbG2WzijyyjIIzb9WvDoVNMzcsKq5UoryVl4a5iJzscmPNpWep
IEHXfkLKtVeTphGad0pNa2o9kUI1oOkIJUAFpxKKuJkz3p7KGy+K710eAb999BCLwHMRmWUMjmoL
CrRWSFqfdtxKIC7yId39adRFAmdDRe4swEWiM4ZwB4YsE4rJ6mF7rdgbFOz/xry7L7yvBw1lD6/C
6SItfkHR8qLCyKPv/B+k2NfrPAkCuT29DFuEAyISGknCy+634tx5XoOJhEZGvRUNs1KT0Hr1Xs8V
ujybH9J0z4xwKBmTuN22ucBrtGtG/XtGXPnyQkSHLRbE7608mJ6XtBDtj6jZctv2C8Mn6bPga/M9
CNJVR497IRn/KWlTcPkUk1JPUlkl5SOlinjFWfvmDPVnaYMK0ipYTOg4WHay7i6RtEE5sAybjidC
rKIhHE0dibKD9ns2surmNNHic69Kf/+1Kre2UXNZd3mDhkGw/MFfQ/2Tq1fvzO5Uh5fw3C9ajdRv
HPEXWMBrNln5/h/r+cEsmY8CWP68bF/CN1k4Bf9t0XHU4+mc9vk1LjsM2r1VcLbFyX13tuB7IKAD
qUpaWbyFcg/54EbxMBLfZT5hNbfyI26xFb5dppgMGzPkp1b30/95WL+clLeOP147omn47RsVPwPB
mX1MsTPXZxvo5ZuD7yrmfItGO5qaQnGLYcZKy0hjKCSPCsZbVEFreqr7UoswQxZKJgffngdFbd0a
ndniOw/8RF4NgKlmMfclCngiBjBi7/1BsErLo9zVt67H8deLexMRonGVZldrb83eGS23YkgUg7T2
SSSEvMrqvRDogJgtc1Quw8L4s4AOyzq2Y1brXUDF0rRjRZo87ZqpIz1Gpo4u3PAo37J0X7rdpoF7
vcY6DzgD+IU0LZCLpc4d8jQjt09ZJeMjpVzBcsO/LXgiLu3cI3bxS+7Epi17Ef8yCj4QLdwSyohJ
a8SxIvcQBsGNWZYBJrUzjr6659dL2v38IHqs7jJHvEuC8iXE/zaHu8BvwpYgZ5bD6k7OgLsKN4NZ
0b57Be2oBY/xTapPPZ0x+x7UtCHl9B69hnDavIKMnPgoLdboIYkKlmKe3T4gBpFMBGfmi99xbvLB
npyfUTIvsUekkDITYIynFE2YcTrivxBfezrX3QmNXBKwWtry36BebErOzxJjm3vAFgwDfCpzIVYT
857qm4ArIxehjEIMalBsvVAlpPQdhwmwzu6azHKaeFiRZ1tWsroqPevyPdIp5n2wA/FONjZI9Oge
dRnCaZcpwyEAdshBBtXn5EDMbloIdeezBxzaC361ZpovVzOfs/nqWhwAzEky8pEjG6SWJfQeLByJ
EKaL7DFJxWWlUZalVbgCpQNKwNf99tgiP5B2l0duty7LxjmMLkEhIsKlfIQoU78SLn4YDNmbEy1N
OI/wyFls2WsYGUXNYkR1tDT287LlsHdrTsG1ZfuJeCgUVSpyLjDOacPWvonAg/pfc8Jq58gw4jdw
L5MaHob7NQKo9/Ored++uGzDpkzGK/LlMXtwzuk4j1t9pZPYXB+Vaqly0GsjUl4kT9XbORzmH/fD
5X91Y6oiSbPInZG2bZ75q1dMmQ8UXLCGPgQvMVDwx+h7D20knKxTT89AweS6PpJI1M0oq4QF3il5
Q4qBiPxaWvXX3m/9RxPB5Xi3HO1oj4O4vBKVf8mnQO4CO68Sh1MSKMbTdtIckIAMwT4ujlzVplSo
laINzkXbqXmoSuoZAuza0UkzOccLuaQOA9NyOsNIB6phDEk+wageco3AxlCWVV4Wx8JAcmfNd4Ds
f3vONenMgigFhkE6H59cyNMraZw5cBRBjLXr2oRqskCE0eEujjZ6kGrKINkhAlktbg0y+oHBvWVW
PTabFFfQrqLLv2deyRuyrXRNuExakOS+pg3Eq0QovbRX3boGxoR75Fck/wh9nbr/g6UZZT9SVOj1
fRxn1Ydmsi0ozntPmlcADw7DHo+HjWopWYusdZ5YQbBD/bG21WOP5+UXqZ/9IpplzmmsW3DWzvk8
swu3he3VjdfT2MqveUDYKjzxIyUnR1njRdTa9THyykZ/6ExYFQZr8MrFq9KYJSVT7cIcMMHGj9qC
CZotZen3T5lGhcIlGlooLOZQfu8k36hok4Aqt+gyMpb9bj+Dd/K4nSny+4TvLsM/y/W4SoqDt6p+
CFseYFy9mUNtr1BIvOT4V/eNeewuSho4ksMIGQKv/VfEzRG8eIePuhOlSV9cvaek6HMn+wbo6je4
cWKnCofLsszuyY0SXdEyu8Zb3dkS16vpwKqTGemJV1SyrKHLX25L2bt8IqHRQKv38+DnRgVT8Seg
rZLWwfwluhVeiGf+qc0sDoq1ZC6GZPraxYmqcsLkVVd088kWBlN3oeb/X546aQy80txBTbmYTXGP
4AhhYYlQavHiIHIizk0hDa7WUck0ldlL1lwsScrW8iMpoYmmwwbJVgoXKQMrPWvS9WgIaP1yMaQy
/y0L+Oz+OPIUG7y3SK+K+A4cCWrT7ejqeQY/k9Kmu9r+splqmsp+cICO8Q3LGdRX6C+faH/IXPbv
2carbp/Mb2o3zZYwXfVM0vkmKl3GjgdIqY7zrTJXwO1ZDZPwXLaZ8tpDF5VQHrdZuvTYWVrMMEAf
7+dxNJrwQxKQ6Tuq8HgTkbzay4psUa/DYpV1mxSXTIVPNg8AiozKj+XpHPXd06rvTxlp8yH9HvT2
PNWeXvt96H1/XtXLOkEGocGgTB349MiqdPSf66NscKHdRlBadCWw6WlOOxhWIZHdAPioOsQfaEb5
h1Kh2JOE1np4Qp0zX2s5jNBgno7W+80w2GRBNGPTcANIuRHMfoO/yPY60lFMrOaKoIaRlozKGPIy
uY/qebt6uaj9Zsm8tJbVpf1Mi5H5LFi5Vf6uMee9fwdzCrtKsMDUTqx38lTJscmWief+FfXkvqyx
qJYoNNw17xlxX9bVDVTWyMUiS6GnWcpUdvB7Yog9DGthlhtbEtObB1SFFReNJwRkqJuSaZAYZdWr
Km1ou43ofbbtPvXUN01rxsOJ7CCeXwjnIl5GlDF3WUYGUS6Gp2HP4ljeLq0HPlU3DTtlElSLg8Zv
2tiCoYqfj+h15sF/gn6HH3+jWpdeXxN4mKTNOE9fPWrYTX5LU8h5oXeaI5vZ8o3b4Dolu/mk1udE
i/jrrRSpdB//oZJ7+xubfRI57syy2RMRfJKZ4cQoZamsDENLQLM/7Ah3NUi3DR3jG4hUfcEHT7na
M/OOfbxFNXG5qy7TX+fBtXgZPhW9QugL/6cT7BTbOyzxZnQ+1V0VQAG1S05VRO/t0oMsImo2nqxz
9T6+gtQ7kf0xcHhNyxA6LnP2zoAQ6eH4zXB1bwqwfJL+9PQjyu1fuHehvj9mSMbk5G3LcjzTUnk0
8lWs7L+X4tW3UzadUJpyxQ02yVJ8K5BWDrHZ8hlOiKF+rLNKTumTwAyp78+v2c1u8QPDjugh0PRw
D5Ng7wWKoBjzpKDjRHzwhhdBkGkqfFhMSmg+qlgpA5LY7BLyiOaSklQHZD11DK97T7LEHHMhA7+L
zZ12E8Z1TxqDuqpsDoWioFMffWVzu8nPCqGobG3eWAEB7m3uICcAk/neBkW7+89Ijx3Rkhfbcwd4
KT9d9XAjIXL7gcxNIx2Z5bCJvBKnpG1bBIO8Cayfm3URHHPO5JYCyUqB45j37wX3PNDo0XNi2wII
NYLvmwc4kkdhIVwuoEo6SMwDK9SzEWXHGUafn5S/rtADqyf1jFxvx/7mThKzzlYGPCHNGQYXV3Be
tpbWEaRPDAGHFqRUGGU3FCdRaDudrUQtoHy1WSBL1Iv6hKqkQaNVoGsebQk/SBi55jGF+IxjKi8z
N/WuJTo0n4grtFfBU3Od/XXtY3Nkhnwiqu6OV4Zwcr2VmQ/esbkXpBDhSUvxkjqpFP2AdHHROipX
jfzGLApjLg33hJXczBGnKO1P9+AeznYA6fIrrp3YUDCTV/AFEwJXKmLXSTTsbc64+LykeTj8cmOc
+mYmQwSGj1bEac9/bHmDqgdr6mItYZRitO3q8OBXypmj3ORq3cYp+XFJbDw1YEfv/YSiWLmlNBRm
FpfvOHZ3E7u5C5QbeL9ZBv2lwLtbLNLSQN2KezEEaysLQsYB2QyI7UfSIlqi8Df0VBUI7QHCOW8U
CpkK1Hh0myZYSH77/A0Y15pHwr8fyi5BXwnlnVBwLfjM5PpSdlp/m/v7ZaPXFJXZ2u07Kus4DYuf
QTI4ZAPrCcmbSPStX3Q8GEYhzzErB/k89QBo84MHP9mUUF0NKEvXOL0iU1WfBLOezklMiom0MGwg
99A+AV8KY4cxaMHEHN9Rq4qj42MCPQJ5lesWBeMiOIrocbDINGNPEMSrQTxAlJyXQmFDcSFCZ9Dg
XIgLVNsYm8tJstpRKlQIY9zrbG1MRzhYkB116Yu+MSNIpz+QWdfzMgaqWaaMCkrThGShjux8mgmZ
0JXFBziW1h3tUYTpEXyRF/BQs9/eigXAHZPGsXPycQ+dz76g+bQ1mnuEZSHFUD9FubR+8HMEIslq
TWnFEI2rw5dMznr6pvpDwT8ACGZ0hiEG61hziRTSSXjg2Lj8Csjri8jSmXcTze5/36mwwVyIZeai
ul/V4Iw0/pTnNAYf4vAISyEE+0mwNHUfkigoInOUDU6rYz+9PUc+SXoYbNVTE/WF3LcnT473Y1QL
Tj6bc9ctievZVpD/L2B5VHebCZO7ofzJtZ7MAwZuzz9CCPJveEDvV3BRFkZ7uj5jZFYyTIMMRlKL
LO6vPYn6CIyTf1GLzQDrqoEDKtvIgt4bcW4tRk+PqWhW51T3wGiiVmfY22tfXzhI8ZfPmIljBUut
3nPDhvmWm1OFDlFAjhziKLMRpWTDdRk2qEVdAFL7ZRjX6RfRhOZNTnpL66ixDiwpz05lzLtUdzmn
d6HtCvN9vrsVYpIq3y1gN6PbhQTa6rYeReXFV7LkkTeToVOrirsMYp+9gXvuzU86f2I5mqp9YK3o
5/WQvw5bkNiXFUs2S135VQlfX/NK8sEh6KVp4DZysNB5XF79FHU9IHEC3IGBxYt9SXtbN9YyILuK
3FB/vVqkMgJRddPvgC9RYlE2l88C0XCNYHJxAvyP5Qkfb9h7vStk1s9Q1CX/YtUfCFfnat2lWi+2
sZEfVzvMcIarQwEazZwyzc+ufA1rWHBwH/lEIj0vzyfKqhD1r6rIYiUyWRrm5RqyDHgOb30yQF8F
uua+zyj19LtW7F+41VeJsw5RGwGgvlKJrIB4A5xH42T0PHkOj19Xsnlivbp2OeEfCuiBZVBLT4P8
tOvpx/MjvxPjSrXZCs9H1oM2eTvvj2EIHA85+yCbxDVQRhnoTTZZ784H2MZN7dz2bJTXisEdzwZR
YHzOEHR/qMB2Xnn8QiYybsG5zV3JNRVIq99DcC5et3HOmgA0E/agGEzltnH0CENWVEWlvqg44fun
uueaviqsj6PkQA1vFV2wvWVkVotwkE28ZoQ1XZKImNM0OZ3QEBswrJwfDsJ94//A/7iKsOIYmBMz
apYGkerA1Lra4u0v2YDR08+HaP0vvGAXYxq/P/zdQwQQ8f/IKwkXB245q6LUwvkRVAlm2VdB1Ptb
K2zC4iQGRl1ywUrMepd9rj9ohmZkhMG4gQgIh87DE8u39JE4TrtzYspPgB74pklXEZaHSM/3ghMF
b3vOgae0dcAHPv/+8eNYdzKHMce/tZF/gt33eYBZKRoemDm2zs1S+l+1M3auBWBvca2D0HIsPoIT
aWs+4DoFLO8eFv6ofp6lme7Yff9tN3iiR6DPHltwjJuGfdIgGrCmduIhK21ZMrwhmxHatSRtZpXk
Mh0xyeEQgvQ4OW3gy7ZCZZl7tLbd7Fzd8NUq1sKU0eBkQa2+vthSNv4aNhTheaPhdfSlItcMyr/p
NgpjvGRT7rrUr7GqXQWiW6gPjc163biSAjT69xaHtpa5Gq7p45Zp91Awew7niwWZgb7jH3mdeRBw
CRwx16nGjrRSTI7ItI6VwqO43yG/3ahofexTS4Vurn0MQ0Nrw4nrUvUN8aexev5KpIuSKHsKlbjb
mZuyF0prWLU6iw1ZOflDI4EHf6ftdacY7TQUZt19Pk1aJPX5WjKBzhWmycACOj6KCaarQX2VVvtU
GalQgxRd7pSb1VcybwjeKg13GqK+FaeEsUzcGc7aV8c7ySTmQMC8rQcnIZSsfhPRz27OT5F5yATS
SeEcxYjWzMGYMaCmrTsatg+CazOLepfMpISlDFEM+E00OU5kP2K4bRNJ3OsIyCFdtvxT/2CT+aiK
ozrKduVDc8cE13rUOCY7TNh3MHyE9lo251z55nST299VWw96adOp5S44Ss0CrBrymz0ZAFcyswhN
4eG23JQJ1i8Abwe30FBGmoPugXfGoayEAFEFFkGnEXExEadOqchrevj9s0KypjLtRFWNQgAH05YR
Xq5FGQrhoBGyrKt9plC1ZelBT9RUNCFeWMxhfFfgYq9KBJsGWL11eI0XBwaDMo1WeYWLwxhRLbxU
3hmPPO8E3XzaniroUocIKQXW36UNf+lvNNdF618eR9Zkq9G/oElwutcHkcoyvqlbx3NM3ZzOP1c1
N+qSHiJxHi4s3/EB9dnazAN+RmMkMq7ieJvHQOIAGRTz0Ach/wj8Fwve192dedvRxBeAO7i2SKgd
wCP5nyLSnak8CJJxoFnOggQ23zQNip/5Bjqj7HX4lkEb1DpwLEH3RQR59t5m3GB8sNPZU+tDvHjN
lVaV7Gkrl8EKecUBMgqzD5kNg1fniohxhq2oW91iHq0rCSlLczqsHW7srtx4mHzqgdJ0AuH/d95D
shT656meVZ6DzejSNRiY0aAPiJu1mFJNq+GolJe1m9tlmnam19/GuTVTIqtIcT7kHvSBckGC0roZ
8OaVpQ0JiNcGqLJh1Lh5XbPzQ80AIXHGj5/0hNi/uBiNFfmzhVTv+6NaFg9U+IR3iHZJuEq6NKp8
NHdqP1RzVHw/uAHbQ2hDYNXdgdESgH6JvaRAroaw0nMwLtkOGd/cZLOrNB3IN0jA5Ci5lJvATC0r
0gobbfBC4yKVlEJRjYYMulSugQG1HDhQWtA05TmxoKI4esV8kAp0teOZAjxMBFySQ8Y22TsHbRou
gUGSjzxc/1UDqfnpk4yBbl5THeK/xFWUYI+q+HWdmryXVqHIfGql9HVZyXkEKuUe3B94aON1ensS
Q0BsWJsUeDksWE/qiownoxPKmL7nw3pMidDXmfG0Uw7O150irJW8buU8XCYb2zA8eLPys4mfIzdP
YMqhpJwBP3axyFde/wXqbZWdNQ5D78p/Z/apVJa5gzc79QbheNVi3qbMN5QxNybU/0Fwsausm4hz
zJh2Ng/4daHy10sl13Udxoul3xvEhvI0UzTtnP922f/DG8C536ZBGBgpLiMuuN77CZ8/SakVGeOj
PTDXdXgOyNCuDhhNDLwFYNiRQT9zFbxUq7bKXo31lbDzwv0GWh+kqFWsjmmmETPppMSz2egF2iFM
5oz1q95lFH8207ziau8CjCM3Qndgg3M1PFMLeVNxUuS2is0wa+RqdgenPKXTrc5M9p0k+8bbc2+M
uAkR9YRAFj/CsBtQYmybFMj+YoPQIhylUb1fA3FbSYN0wUJqAA0uSD563r9tiQlhQM0rC6bYghQ+
ELZfSfKQX4ns7W31KPuJfgLUkm1qTIId26smE/zrhBYFbwExj8q0XZAEHL9Lt5D7ynw4ASUaCH2n
Hl+48x/ushvd7OvOi3ave0Eu4cQbUSQJeG87o+QEyEH2Jef5bgDOxYgcMNfF+7KfE6cFF4f5oqj4
cn4Ti9mfCZHE7wvVlJoVB2wmfVASEL8W7XbA+NYWtBOslRwzYMSfxhQHo2oRM7XE/QZe4aggl+hb
hVGTpAK8SVgW2rf7aX7QhsvQuOfolWNmXkeGwpoeyCKKUfcMKs4w+FxH16k220KnXroswglnQwuw
LqIIOQOPKi/R9PU/nmsD9F9N2sODdF81aoq6sS5w7vGQBKIJqziSM/WwzwVBPgmdrBi3wi1aGlzc
A28nfrALTsnObhs4GGLMzhpVmbAzHDrBpMUmtlYEi6z2voN03mZrsRjmOEL24QFnkL6udfn74yDN
cW3QboyGDxZqyesp/3TGLzsk8aKDfRjM1MFgYoYNqsvJxnLcnmOWmkXQ7xAZAh7KpngI8xWntaPD
0KMxc2BdBjhpRRmBAOYdCD/YMz2gumVfde90F1cZW5H6jWuq7Ecanekd79unlU4qUqspdCSsjqHT
SPqrlfhjdeCXkZrNHjCp0sjEy+S+7Etzf7+7wi24MiVRkpC0xP8Cwsbk95KUzqpITASIiNNpVtML
8K1hop5rb54a8G6at3F8KuDj7sMuCsNod60b923HmFIwLrFU/r+UjfGUujpdynX9Zz5N9epWhBqz
4+RAyqmw70T9pVgiLuwwqQFEtUL5JwurBNB5zC4vmCM1XxDTM5OMs7UkIxuLmNolbcANpPke6/qi
GrJd8pLTdFD5vb0DjJdmSCpXJIPcnwSqfgSpED4TMp/2OaeycKyWsheKZ8uh9wLdpQCw24n119kF
GkRfmmMGhYlzaT3lVQXOJrog02oDzsOBNa1P5WCvZf5Rd6vv4PqXyxrQV3GssD6GhVlMIGus0jH8
r5euG5lsSB/xTuruvnB4QKsmuBU2T4bQJthZSK1yVK0ccDjAys/LVp9IfXY44N9H5YUiPos8XvVJ
kybB9UQxWTEfl5gxGhSUMUDoRxT3cf/R652Gx6YZLnrKlZqGylt+PUL5WMMnpkCHcINkG1yypXBe
FJ9Y5i6r9kpOVlJ0VGcEzR7L1D6GuFGcPVa41wDGOtNRarRm66LRUYysRH45rNRD7NOtFgM45XhV
7/cuL8Yvj+QBfhARf0c9OU1SUfcJNi2lntYYwvGyVEZRP94hgd26bUJ6/6ae/LPraPk1rRjHRoLB
2WgCCxqzb+m7KieOrZx3TeD0iYFXi7p8JZe3o8JMJ5t4JxNwIrnhC0x+LzXFyZ6KDiuCJ9iGZiRk
L5+OVYSDSBxiAl2EeHYyFxgfZfctiA0M50VtdBpc0iO5WIWL1BYqVGSSOY2G+Bsemvn9mNR7HBdL
2k4MNeuh6D2UuORIm1FNYcqfSbVfFPpBIvG818nsQFevGXlxZBXytO2bMaFWdVuL4DmugL0NibDz
vfM4XUopL9uqvwvJA6EfXnm/FOoFe8+QmS3gu0NlivjulI/5j/gccMXJzSLQdd2jKeY6deQ0ZxOA
JQCpQCudnjYPORjdKa52ihdVUP+lNQgT3SbQXndZjXR4uZ/04MZAMZvjJmlK6wFK9/wqF0dvj+2S
WGtvMsPOZVKmCTutUzaATJMGuEZcGRoYj1h7RjCZcI8NpKJgH9GiNlzMcVveCB3nXQcGmVCa13LN
3VquiV1TMNuaxhCab2yQ9B42Iri77n0Nv6PESfDVIB1uCjYuCaKMQKoOoyL8QsyYmQlB9GPhEOuK
T302GWo2n/AvVyOkaBPs/EJxpP3paw5QUgPusTIHIyUokZq2NsC/6RcXiFcSreg9sDLsO84+DoiO
IEGDN1ysu/39BvcI8YdsFyFoJz7zOsp0NTyi/9wfSOKluy5vL6G5rZZ2xyLgh2JlZnchIHWbkLcA
jfyIwyGYGK5sPWDThu69HNWXvsXw3NlpC+GTT5BraRR/qBEK8SSAFXCANcx8xUf2JCDXtUvwmz5b
aLFhIZaru5hy2uHHF2hGXA6eCK1lhTxiX4HQzqkkBilhnQY9SVDtTY98LnTUjRmrPUfOEjN4Q0nA
T4sL35jBTKWqLYN/V53U5zBt1NEZbJBLrojB87HXLE2gV/y6tAW5PAwlwCXp5DjmKYmsp/q7f5BX
JqF8j8ZuZzVGihaWZ9/hhMDdwhOxmz09Vo5VLM2YM+kiplbK5BJM+kGcySmBqXGw/4yathYVnq3S
QifWXswwrGWhZaJhIU6qslES2Ay0Hv5MWVVDKl57Vv5+lKHIrVEbFc64wP4ZYV++za8hHoc6n9c/
lM6FiXjjSzHYY7+0Vowo/HphiZfG1bNEQs3waIvO6jE+SjhUeaCLeX4XD5tmGWy7KFwrjsYlP9xL
6uSrNnVx/FqcSD36eY6H0mt8o1YfnPPkRLdWp4rVqptezXx436He4GmDAxaMHPS4er9E3N4lvd9L
9ROV2ZFdc0qD4sPxqWY+MmaeFmI0VQpLHl45LBNVHQTzGakxwlJDgEVD6Wow6Lsptb5vrlj84PPF
hHRW83o5KcA+qULVcZHaY87MuXdvAhrwMQheYwZ2pEBq0WilL07Xh3vcwaNn/P2ZY0vUEfuQScHK
qtaWR4DDlKhLIRjS/Ux8pYTpIPbh7dYPlnlB+h6ufBZ33hpzaXkFihPIsCpCvt7nobri46duMCEo
l6kiA9ySJItX2PIUDWWNeQ5nQqcih5VU/bk+eZUd7Ah3PkRVM2VSoOBA8qP5klwCF2Tmyo745q0T
vvocGmpMzKLPveWUCGfoCutWEdw3GIu+9dsI18P+xdAburBFzDvutVOwTig5LyTvtovOQQ6onOF1
cwoFDiFHnhTjklUbiHja+1jSlvySLyQZUoXuEsgW8eeaG4GReoGHsLC6h8MndTg6KcYEmmLMkFf2
4PzWiNHMGxnAMhJRU9NshzzzSeL9Zu0vvYUr+HKa5J4kc1ffJ6YMoEH0K5LMNkfG//kAduEm5loJ
W/m5GC0qCy0U3Mxbttswsh0a0TfxCGPl0nwXs+6qwRbXhTfIYdCPzxLL0oRwHVlkRquD2ZwLKHP+
MfrhYZZMF+GNxim2219vcfJH+JcADL+sLdZRCPCKZNCnD5vBH33frfJFlsM20w8KO0BDmO3g1hao
7bCuGZImK+FeKLwC6MadErIlEIWdHiLDrDEIa9YHSMJiExhjhvVzo8c24qpH2R2ElDq9O9kbw1G2
ZWlI3pdsa2g8G/0t47MExaklMY67tcOYA3nha/BmWccASTGBGqv1V8SXhQEHWVO3/jBRp2GFYsSL
w06iLnIALzFnLe8TM1U+653yV9YxK122mpC+fIN/xOWnBcVKPsz2+rnJ5VTL2Q2dktfvpfDv591H
vcWlzOoAXzTumH2fV01lIayrTjMmKRNEQqrA90vEXz+RYGpUa4BPRAl9ey43ucXFiYUjU9lm95X6
9lVewmntugf+rNTBKwKbTbsFvoicEWS5rYPjzwkOoXU6LXUZ42f3e1kpU5JPCpqkHGBJsMsENPCu
i6L3S/6AS0lk4G+aHFTz14ZrFu6Ws9Kq257A6n0IKluQqP1B9hHzpAJf4HnmH/gO+bXwtqYIbF0i
WcCwrV+HDKphX/CyZmD+Kb2n+dRrk0r8hsCn7yyK+EM+5CPYkeDhOCrORsGjmpMRsFgdQkhe0qgc
V9UGM2GVsQFKWWxKim+r1BPHgqosowT7QJAPLwrNkFn2+LyJbqqyaYWi6jz/IpaPNZWlqBa3ZZd/
7nfrHIPXebphgX40NeNpjBF9pvUvrTfiGZRld3wzbg1JKZ7Mlrq4Qlcu6jAdnW8DSx8De2GFEyVB
Lf5MIfGnRJrceZxbdpZnndySZ/U4yQbjk5eoSoHxfVaaHDd5DOMwjYJO+N5uOmo1k2lOpO66EYSv
/+Pk3Qkv9GjGwhlEx9ph1Suex3b84ZYgTQpwXLssvDZMsknKXhrWcZpsse65zitRu16EkwvLlFVZ
tyIXsiniXQjLTN0aB+/7GADVzCy3wzFlISSSlRGarAMMBiyTDtDh/4YoMYjUmTJ9saql/X9YanHq
J9zyG3UOMmA16kPlysN8kSCHbLHZGWoDuIq7A+ow8U9TjP9mEUxS+ouc3CrCBm2VAlC4/oVHSVZU
D69TW+szyMuzWvXAiA855Sw3BRrzLl64YgaQBrE5GI9Ma1ZOhfJzwuZemCcTWd6ZJOjtlsTTGMb1
7S7XjPV/d6pR6anmrir5sYf3YhmFTb+33Jejl2gz6gXMHky2afZTJzUrXzXj91MAbBHRYJ1FmEyg
uJFCaQ2s0IMEdlWhvi72Lo2KbwI0APSpqFTt7Np318TpQooZDdVv7e74HhqFzO0JIiX2I0ZXN8oI
5QMpLgLaiJ4CK9pyC4uuKlxNeN9513piQg2oIxyKErqlLcQapLnGgNcoX5NvaJTa26vrxwXhUT4e
OJAxTsLhKBzwwigiaipB4NBx9zLcUQgrvFnrp37L00PeTb2ggIboS0gW9nK+T+58+UwrWRKt2mV4
f2mLrsU6xrx8sb4ni3m0Art1G7k00ZX4WkpDPvEJ1fSwY0EK5apwN/kqGEmUysZyfQJoGXT7ZfMm
l5Vvh+t6vVHAPKwg/ltA0tBYJxON5epQ9JdOXYdRtSD25qbL0BMqnhM+GvejnCZLyIx88NhN8vDM
fKwbX9i3Lx4INXK1akdMn+ZZ2Wie/YfV9RbxIK3ye79ZFCJAvjUMHlZ1m1JLkkAbZDICWdKNX2fD
1b/gdJ8fWa+YRECvAoivMMlxTpuPWbtnXi9uQULhUwwaeTjOjR91QUa5zMAuNYikijXLpZekjmTV
BfUDzWGY9rsnZvXVvj9r9kxJczfwe0a8cqPEYLSSR6Xl+U2JJHMzb/PNEOpegn0EQMau3VFfdG0j
2v7lTl/UuLaOdSUcmbK+G7DEvgeR/TcU/QUtccQkj7xtuGTc6f9k5j2DPU2sjk2C3cOxOPPVHCJJ
2T9JX3oQXWRxaGeBLvWGRBi+kBuOyOWB/hg4O8O9vH0brWVHuIjh2Xl4zR6NQ+kc+Y7cp1nY24zz
3ZTsghiOzfPXdNkwez+23mSPX4JFPZfHWo33PCEab0e4iNhtB41LUl+TEurPRooCempVXw7F7KkX
vxfU9YCtarVSbv0673YiqtwlKSWhm7BmJHGRRDKs6FGhFRx5Y0c7hJw2ljRxrPJIsSPnTmTL14OG
E/GjJ61PxayisLjqTDK/mVlT1sa29zmTu5xL8EZYNfuCWU+FJpK6p9oVp6v+Edg8FbxYmtY2hFTv
p89Iz6ySwcsMU67nnXocJWqUuk/A6sa4Arca7/neiYt9E0IwDF2n4X++0Q3vZf9pm+w5Tp6Rq/KW
QlbtfqgGg6qgeqHhvE5hdLhbRVVbWiEiCocxK7MCOgPEhqX0hD/l4vcUwo9NSLExKC2jWB3yNsqA
ECKq5OAoXaBOZYG9TaPR9EQcVgHfEJuedXpFxTg0gJMDbtK8iQOrtHexflUl5G8AaAhcTuTgkUHo
JcdWVnEsTa71x6UXB6aiiYJJt+aIgfoPp53FSzvlJqBY8k2xXh4d4fOCoJ8f45ImxtNCYne6uey4
q2L3O+UFFg6io2emlXMyqV8clZv5R755hev03rkO3+S9825f/RlOpLO8Y08WvnuXuEyCnZ4Pvq0h
dnFvOuEzNHiBGKlqeJfNUpR3ItEtWDPlZ1X7NyGowqdt32zyfcVTXY4GszzlVx3T+9/5l31nqk6W
ABE2P/gXzeAiAMLSxDpJXVOfDCtIEWqkTzr7Oto+gC4r7+wZRzzV7i5Ll4p/xQJl6XAtTaUbAOwo
N7XTolebt82yPYNhmkjZyxBpk/s2VaZQf2pxHtcG0H5mpOgt7JuTX8E+YbYN+8wwPgxHCTFU6rE5
KeyKbEpVu9TG2UneaiPEFQYISRcc33f0EOw982A0j20uagOs9BCmu5tcLK4SVaKkAXjermUMV07i
xPMtbWs14qGxAx/QKrIV4fkHX0CB3sUKA13hmPt3jSD4oYW+yeTWAWEO4vCMw79QIUTfsn8mgyEe
sk8+gAJAlr1Z96rq2CZfNVRSEl8nNCw8p1/OY4dsFxuqw4GKRLekfPi/1Kk1/umvHBQXZIk9JZAu
hfzAXRXv+2Z2K6avrPVNHlJscDOcqWy7Jn+YfY1j4DftPKRCEphlFqVqFUAzXV6jOiHcpByY+MLB
2JTt1PWPReAPrFMdidy5KR+vIXE6BMw0kU1Dcy4UlTuDYAYtl+xVbf4/6sqYCEA0WgLjdHP5Y8OO
LgVGicLhoUbUxEmxx7fvJiMexhSGHwPfDIgVK4eQJ/mXDH2Vl5QKkl4tx/0tezaWcwGfNJ4zFi9F
ajwS9jhgFQp+ED58WnXdUDlk0LkxIA6NfWnJXp9nac7dux+gNbE0vgTolAFRBuSekOMn+wfAQN6g
4garZXvpMapIRGtzrkzvwbORcgK+Le1EIFHO+0lR8+ZxSUh2dRhxzV6lgksFeB+udA0jMaEZfPRu
ePnvtZ+usQuDA67Nri+LAKK2otOqmZz8YL5UFkFuEaqB8xEdToGImAoANjQw1/dXIKCpFbi+dO/h
y8fIzrHomFFOHhKOmuXtYKWak2TnrU3lKJRE2b6O++fUUme6s1yZIHMKWzqyJA2ZY0KXDij2FceF
ajNL1YihJ7QyAt3N6sXYuX7R+wP4jJqXn6x7YK5MSZCQCWG3EWgiEMQfe2kWw1RX1OVT95WEiEF4
nUOVdf3ublf9kjP+bwNYpaX9zC+JJ0lCoGdYBQY8PdDdSlXDKHfxOIHwPZkLNTGhnm93nYm5lWbe
4v8IKYxYYCe/GD6UXOXy+KCmu71Lz+1mm/7od3Dwd8Ma0CAy0fNmj2tj/NP4fKxycpukII02c+no
5uFtdXy0oNx4MxUPmehZv2juyKyjczcHOImhGopq8DCBAbYKWT0J4tkq+qUXaI1txJW/2XqIRY8T
zcmQZy/GnsCSWkICD92i60bgoSZcZuFjiQsXFgNEI71q1uU+PwE+RWSEOdQryVOfMFwUJx88by7S
b2bKqcwHcLVohh/+wyK3iPCeaCmGkU+rGyd/zCg+/7Dwhakyq4gIUqQBgEDnlaH39rR5LrDuReRJ
U4PVSsrASfMBVjCLnyWf6THZ5v1HWC9J6kRukkZeahrnD8NTnC7tGbUyub3KTq4zXaZNzb7Tuhps
MVoUavq+n6X3q/lIu3AtIypuavy9RsR3vVKvQFMxBgUy6s74xMR1xeHkle5eBbX3zbq+8t60GJLQ
N9WADc19AQzorpatKTvbMhI7gq0uXpMiNRfA+AZug5uw7MA4Q29Yv79K6ty/tQyI1UIoprGwLiMU
crjiqk2TKzEBnZFqdiHbaZnrGcRebfgiObXkYKNV7mCBm9eUnqggBNsjsjOX+fcD1ZGKD2tG0/V5
Pi8/qSiyfZL2a3aAmaCZhi/1xrd7liu7dQS53G72sarSNnqDoKaTFgtPWUyh7WV5+QnFeIWXwFDK
u9hrpPyNVX01T968q45tE1huTffiqO8NXySP2SR7OodsH+sgQv7D9vHBphY3mDRLzuTMlx9mXLPE
xoBjJGQwg5FiClLuUuHJJCswSVMpyx1uiHaFKjyg0b4QpLAxCb9whEhU86t6oP99q4epdhFCuptU
xBicDJTNsFPmzZLnGTR4+WthH4cjsvGbO1QhktkU7tcCWMn59n6chyF6RxsifAj3LurWW9rzEpcR
j52ol3u5f9hx/6jtKS9G/2RXdB4y7WnLothE+CuadfDPNpCdo277zcYIgNG3QGmfIFs6AJs0x8ZT
so5/y7+i3kL5V763hFeY6GYGx3JTY57OPYa4c1y6IHbfNtTELdlGSqYJrjT0CfDo9x/BFld6X/bC
w91zMlKmhPDjcr8hoqeI5dqWLya6x8v4ehBDgjeEP5AjXhjgPYf2JEuodzmcs7VXdITe9lx1TbdU
m7LhCDygglGNF9iwOjVc7z7nLMOr+ex/B7WFRSyMpd55lZz6fo1Ply0fEVGt34sLqI5OvRPs1Avo
cGWzY1lr0jMm7Ukie65/wuA+z7/w/lxcw259mLp5Sj1vSQHbM6mWVOsSs1gTJYpjl8t3lIszmoZT
64Xqgc5hi2f96AxRo2OByQbUX7YpwCzq8Q6KsMeqfX3Go3IlPv5KM5OdWLWbpZDSA2/314PTMc4K
NgaBf5Wh1EDNLsEuYNtC9Y0BpZEIK1DqezJiLkhluzziWZTdSns5SpDbXqD0U9o+ilmU5D8EF3rq
UoDuR+M6HfC8sIr/Eeuf2RvvoHEZVgttEoF2pvFegU+sh+6Wc8uzsQqQ1aPAtEB/cPn5SZaoDHi/
SB5MQudUt2+uhuQmeLRH4qM1FDTb3Ikn8pANPnufssW1eN9Q0X/Q9xcVbTquWsTavveKX5ZcKcmk
5aVDa6cW1WcfHbV3CbXGndGOIlycxXjfBMifYu3M1SZgZgirn2l6Xyf5SAIs9g2cMcgF9mFVt96G
G2yu0Ou7w2t++v/bzl7NZNOpjMVCTpdl8IJMjHh9ogC7TvJDUCC3xtxOboEEN3h+pHiF815kNEeY
mjZ88KoqxGSoN28/TTiZwa/X+SJjukgE3ppTC235tRUdJyAVX/Z0lziMy/B7qHecZkzFRXLJiOFe
JfirC2nA0TEidHIaNwvOUM9UJAoTgKsod3l3MkoPvVzFvqCBjTCvlrbjuCo+fRp2+NWu5twH5g7d
g4K5Ijvd8LhEQ6//325UF8R6iEqkNjfMzLANo3CEvbcjuhc3dIAk/lKv7TcCYGAmRdAjiq1sYHBE
8Pb+Bt/QMTRyjsCuDmDc+hEJrQvDzzxKOhLdOCW53cWaB86rfsp0tWEKbg972Fcx7LYPtcQ7+YpJ
0H37PkU1C6L+YwxAnJWrfSYkB+DbHy1pLTCgJGMqhBANmSTrPNwdAItZnltOlBbdaYNiIfCmilp/
BSTYaKIWUFt+9n+AwoxbuFClyh6LLoavOfKM8IAfKtYLivKOr6TF0NmwEUu7sjw6nUYq4BFwhqvz
liqCvpClxxRQJajTOlPR0B0Q93aLEcNUqraqGMOQKDvMOIBiP238UAiuTjMHuODofc//N86y/cpR
UttoB917XRzLN2U8C7RFw7YaBfw0fEoj36cSigAwWsNt8jfC0k91l76ITazrTTupxpORV222VpaQ
iu6+86C+EC+ykP/d8Egy42keOMY14NgfYSfyubOzRYCwb/zHF8Ph8lsWWAY0uQ/VViW+eIhVDrw+
pJEQy9IyweMWScK00Rjr9Px04XwP8Zh/Emgl9Wr2an3fnW36zGQm2tv+9YgiwAQr6kzzYly8omef
jcSA/VnsPdFuN5eypk4hgd3t9C8wTgrKdPIU93OSsAeDReYiyjHkQ9JbHL4xCiPHvpvXouWHKAjx
AaQQDpuIxTDKpi+6SkPNdYHBvyUBPVULkwxAwD+JcePCrGzOrXZtqNNCuNULzJVKh6jYn/UNxq1y
X2H2Kuqt2fVTGxvM/icazP/EZhAJ9YRuXxEkbN56u8PzboE0EE3eWqKD2GZzunAKiRwWQdemUQbU
FYPcxe+MGsPSnw6/sHtfKeJ8rVtMuo5M5bkp8weLulqJ5MhSGztQJmrDE3nSsDLNRc/mMtxGpUxn
KGpqM779yscw5nddlpRJ9eXffIeaaP9iAzK30Nedt4Lu1TF0SN1oR7zUoqvkjUtHGjd9uzjshkoW
SFcc0w96C38zU9bu67HP1SOPPs2agMdZf7x2uS6sdlTrTy0YnNQjxTDDA5SHKU9P5pF9nAEp0MoX
SiEqJQDiIZ+6RxGV/2iIAT62tEbrksnSI09lLYOXzVJNy3ZKsbv5y13MfLxwKT2R5w3MNdSoVnvm
7ZDlsS67dm/fybBkV6dJ07zHCudeshGyVD9Z+vz2+qg17h9l8e8qcNLPO/gENuPKXBWvxoc2RNK1
3autXN9T3pDJsKV+CVUqBvFTBawhp4MS1gwWxKIOnYjI1ZmWMEpF5jWITFUZYDSiUE5KEmC9pNZd
OyZFLPX60WyVYeYw2lXtwmRFysNKG7lbbSBrB7MB97a3tyZmtt1h78kBX1mJiD/n7R50zjiryCSV
h9ziTQUVOgy5su3AJE/yVpHkG8O+EjXWAU+aLP1iqRbKpgUBc1PjaOejXBVrBY6RRimeiEdxYNcd
QsUyg5TQ+5T3QXJ3Dy+dn5FcyVwkdz7YvlWr+a5CSDGwEwth1oOkxB/ONXLw2FVpHXAwFdcjBpza
EZFtx6unUlZpJKyjz9UcA2T28OhB5blbgH3fPYv7DRUgPZGNNazdcMWEx9emrRsSYYFaphseFYC+
5YnS6OLdlSiuk0Jz3ADM2RkmB/CeBysTkPrvIAW1/KsIMQBmoci7SYZoGJKyAPvI3hdpQltYO+6x
KqinDPEya7UBgoOJDsKtLruRShwASb6B1kE9iyW+DyFnzj3/HSVNlfY3vw/5XfLS+6vGh1Tp+cFF
nA9Wa0IaK5VkkyQKhbt5urrjGvIWTTGYeGx2NdNuJtaM+IHcXzrmwfut790f3j+mXaDZ/B0dQjjB
x55yp87cgw/qkJXS22vJ2wPYgbyLj+uC/DwdiIYTrq01AlgXxeHpLrUlZ0/Qu8isDjaN9AoB4lIB
fSOFQh/iL1Zn/VWZ1CjDlPVUdeEK3YEhKeRytXM5VKRiP9Uo+OneCW0svsSOzBzNV+4lm7X67LwB
AqgROXBs/6IrGVEvgPN92rU9hU1UYvSq9RAKQ9vxC3zyx3GJgO6WTuXxS6uwOuWM1MPsuMEe3B3y
CJ5I5w80epQwqF93mx+piKsf90j6RQR1jLrOlZdv4t5lqCi+iEY6/Mq2kq67ohcn2gBCsiFx0+Oc
aGegnHbu72wNBCMFxz+DzFhutZo9zhWQNfiGxOhC7IYpb6hPF7+aw833UIckeG6Qc6FjHRm9zDWT
RdaPhHV2btq5TZ9Hnr8g++VU88TTYDsJ6q/Bvk9FYYvbiLddV36eTen44ZUbJPjO04QQklcGSHcw
/sT87iQs86t+2Q3ibAXvgL7Jb2jgYTiRx8QmGRdBV4D7MbfbBl0GlW9MkcTH8hHVA6oXxbR+VMj3
wW6+pMTQW+LxmYYZM41ygF+1N+Djz+zerUT+ECOePu5pO7iNG0/mJNLg7EFdggUXmQhDwK3v3eh1
jrxuppPBWJWtmea60/CdtNnNGhnU/uKSRYoBlebOLWOue2J1eo0CcEw1sG/cboS93+24nN+LRk1y
y3YKgGo3Nr1qfnPfnGVDhkuFmUw01zS56OYpNmx0BYtKijPFGkDSN8w5OS5WiUCCyjlOASwgHYeL
igX1UldpSkEsG8KXzxer1O26ErqCJS1l+P0UIdj3GvYwDGW8QoR4Cyhq5uap0DIbwinhVAAlbGlt
riT3mhfCTaUl8Vh06sCkW9McYTxslqSt+sRI7ZsOqhVll5l8Nbw9om6a7rjibthqrwbBmwgz9xdX
NfankoybWXrW22VlwpadalDT0qneYIeHXB3/MTybGJbN9VZF2y8qCMKQSqUqB8cmsQgcBVIfIVhR
PX2E2NpNP3MMgk11RTA1AV7k56oP1yISIBhEZUs7BkyFHA475AEsyKphwVCd0x2lkTnVgmVcCCVz
pSHuZl1/3EDm2D1keEFvnIBH0sOWfqGwIpF0SrGNWw3/zozcxRf4SMkQj5Euzj4Ev930hPudvEWW
e91VoHRGk4zsiVb2fGLT5hipDUx7s342G/m4STgAfQ2inYWYiuJsK9S6xoXp5s8rVEX7YzjBch0v
D+DG0y+CzVVaOvvDjxs103HfaeLTlymcwlW8X+hjWSZCHVaFvG9M6OGnNnRt1zcspFy3SrkOIoLE
2FcEZsnF1EwfDz2RkUaoYf+HriE9EFUg65l5QDgMyb5eh+Mwe7dnp0UnyrOAsxgNU8tz1Yi2xWyv
zFPeHkWn7NHk+omGwkSqKE23IBJae/N9+g+8OgmmRAAhsapaIGcMpAGdU8dDN0+iNDGpCVBQl8BY
7HO6wD0bT6b+eTYpyW2pQUOvGIK/d6ReZCBqTn7T9Kyq/WN20udWH7FVGW1CIFGRJWBXJ1MQ71fF
gp/sXQm1lbYxWJ0hJda4qkjrD/6KTsdTOkj4Y/W2q6vYygqQV3Ef7Wt3H0NDKafb4/3FeaO4s70/
SBt/97C59noHgoVt2eXLKAcEouBTdLqfnKd9wav+wikxk54FH92qw7o1VNqbWQbCSHK6f0g4kCMI
t565f3z39kmpDJvfKuxcbdoJr9TgjTg/N2G6GXsajyRRhcb6E0FyADjYjqKtetbS6Z6Htbd6wpMq
8zc55+iOjnZN25y9+NrjINdc3qm7cPdZXHzqn5KaH3HiRYaRmwnudqvjaeQDvdvOHaQ/G9NXiqPQ
RGTNm4sBa3EPfKYKL9UXwpfQtP91hUyA07U6b3Cb7/dlcF7clZ1QfPZqf4M2jChhCwUalL0/+RZ7
/xqpFRjEio0ejJQ6Me3Nk75OTlPs31a9TJvzA0AXCIeWbunaggMAk+mciErdmJTAQ937AEeYdiUs
oLuaO6BPEPVfhuhWAQWvyXnTMS2pVxUADKpNrdsENqPmw3N6+6puVj41NCP/7yiTYIxKAhFDLHOk
woAzj9vegmJhWlFRPieYOSUXA6mUug//9YE8UreJTMMWD7An4u1Y37vhjV+FRPM220dVd7sqx02s
OZ2hoAzzvxPKCeZfrn+jCoNI84LXJGpxszYFJuSG+Ah72SeDIAWFjv4v1ZMlrAHq0VfAg8uYt+SR
yfvePenihas2/w+qTiF1wqO0kb+Wf0OebecWu2bBQ3W5Pyu34fUAODIVBnedi3F0aLzeSlh6ehTc
7ZPTqaHy1GLmYmQG5hK54HEQLGcYrLLRBIqkZpYv5Rw/IE46PjsQ6Ow3ngMJeurdn09cOcrKRZTL
72qcyQHREZbRbk9gE4cw4W7lIf1fhlf6ooOquSpEN3poL1ly5rrzd1k1smBxy41xWB1fzqd+neaf
uqpYJHr/zc8vFkm2cZAxm8ZZZSGAhhdXqlhP81ZxVYCG2WWHBH5t18GYfjwR8i8fl26oMsdHKqow
BDh9dCbpKG0UPKkgIoYmjdcsam7A5f+rP0P/vwGlFCa4mnvGsuD+bCPjFixpb1Upn5IE+zq8H+64
rNZ1xb3gPdc5LyKyrRLHIzdKMsvfae984vrh+AQrWWRCol9IkC52bl8lrnSkqpBFUEiWIZL3lVTf
7wGtNpNwYpVZnJfMFA2DVIOVmnPIkw82bH1WaKGtVZ8g9u72/+yvCkqHwZLSg/7wYUe32CE3Wr3y
QiuD7Dokk7GJWpso5KEK4ABMJrLC8rehHFW3lREpP18ZWZfvanKp3wi4CE0+rY9Epax4093hoyeO
zDdDpd/2sHIGTL5GsYiuMjmWBYDgXZb7nC9INR8rywF48DCVkbpYu1q/W15V7GEwDPBAORgVTwtt
8bEmg0tJkAfQXj3n7i6n1JtHmVp22bvZeIDyF8lSgi5bfatndL9sOn/owCB2KvVRh71XvgzaShZK
gpvxHfJ+GnnnB+VJVylWtFs6FRcrt8CBMSShk+IH9ykJGZ8J/+GZODZVPgFlIkUTOqD627XSHRVZ
vxZCQrmbEwIxqnc4jdVO4fUkytfl9OgRkPW3u1+dtFcuEPWzYivKhbrw+MuD8vp8FETW7JsJ1c8C
UdgotwyYODc5GUDIweJrKIuQY6twpS77zcFQLRoYvPP3BySpRp/tuCA2WwAydgbZm4w9H+4KxoBO
/FD2mWte7i4x4MY+X3wfEMH1jOSa0WcfUs3JT1Shrf+JVJjxlUIebp30X/CeHy9t3cQ5WzbtalfU
pdkNY+NPtiEOjKNshXFDe+/PmHwL1tP5zpjZIvtJww2z6Pm47SDwEqaJyr6nEledTz1vNl1oDT0p
61/U1o8hcotnGv59ZAGSVgekXkEaBtt0gdLbycFURsgbQH6a1Y3gb6N9KscfFNeAevpQ5ifT+POh
uH5ug7WbHCPMvDKr5xtiQnp4mGHBLq8G+aKBtVat5WJ39Sfd/uSmB9dvK65BLTDzEpxI/gK0KsW3
MlxtQDjhhtm05d+gVrMjFvO90au2LMXDyq95v+WanY662Ov9nWshNr8bmpKTuB0tpcXEfN2GO9aF
As8s7QW9wA8796/pgmhdnqfZ0Tmw+YlUVPumXXdHxNQZWJ/wx4vHV8A5kffBVLPI0KeEzDA15G9I
HyhZokxfrEWoS7VoaTGQ+a3t/efiWWwlhr32i9U+bdtDJ1APVp1tZbR0P3DctNMPg53pGfrsJ8s7
088OEr3qJJ8j4fajTR+mpPlPBxFsl2LHzMjoPBpCmwo1wzDGMkUpH13BHUIjh0O4n+uC19IRUFEl
xtL2QPsGy4OncHLp1w/RbmTF+RoHZ+6VsomZOOz0zNXrXEVY//7Sb52np9k4yJDM9ZgYMipuW7h3
p6fGWP9PxOnMfSliKhA95zfGDILApzOUcd+/f2TTBSFjq6sDP5EgJ/BQbADBZa5Bfb0xvQ1QMg3e
BtXgO/Lf9tLTUwDKtQqUbOBkqtA2am/TJSydpcclT/qgc85VMGDxtIROoCPOTDMMk7MtflKO1hbO
6Q49r6zH1F6NpPX1oPtvJx8ML4ZvoKBTD4dLneGPWDgTYwW8SUdJv4VBQs/z9rUiRtWFLZrHnGzR
fl6A9YjEdI1+6iULDaD5B9TL13vm6bGpt0zudlm1mJcJwwBc0mZK4zVGEWcyYrJl3Ylnm420WtwE
WhoaqEXzgMWx8diTNYf1yRaxkyxZFr/2+81tNKTOVtjif8KTV9Wcwg3t2vqXasziHdwyFV0glmZ6
A7CWx2J7GgpQehPsgc1MI306dOUrGfi2dTW/Ex/cHpTDhbGCpcuxqpbZ/RXe3AiG0O5Fz93yfLVE
r0lVCVXQSqXpTQBESwOcouf11ZJ5KLErg0fPMNnklA31hFW0sQBuCPnLHX9BFSBxLc5frmUMFcCO
DEStpx5l/28pv9dkdo/GXU27L8R+DXwrLTnRIySbCzH6CSfqORltgLlUtEWnEBEf8wNaLXV4lrnO
JP+z2RrpFn8NfdClvBhSmaEtDMPwaMSDeefMP2uYwEDnkd7EKuOs6yDNmsCSqkwFyIez353Y89cX
FQUD3Wz28iY1JcK27wAAqWD1H6vi9S3UmXDzJyur8433hD33hsaXClxJhdS1jbUF3BNolwOScnsJ
dP/up7Mbr0VpnjjtbL2u7/tEQ5yI8GmCdcaEluGggaJilvTXXvigmzp7LW41euHXqAyw5SNeX5j2
NdrAt/o7MWJMNkXmei01zzhwzNOoK5aJSgHvTv/R00vKunUP6DjXSKWjNm8HfxOjKIMCnObq4/dX
3pxaurO42E3hfbWNv8FPAaGVcC0RIm+pZePto46YaoYqW6wtQ6X2Pnp5SnIlHVAie61LO9xOCW5Q
MPRQ/uZhyIt/dHSB4XNbqaoqkyTNeiivgL4mQ7JQCbcpzlj/jFZZ0pio9mgrnxzFDGDFsZt2d+ON
GUHV8Oo7svSeq+vwIm7gKMLLYr0xxJmKuFKZ2sof2Z3mAS5b6caTpickcEpceDhfteqYZgMQDRw3
iDLFTYwFPwlDvBtpNpIIfGCOLPGQuIukHClHiqvSyygO4O4a2w2qScfHA/GrC9hrYHB1VpTBPCBK
LB3OAl4ORYgcY/SedTE0FqC7Qxh9RfFEok9pEt38H/MrXll2S6aEUa47B9XtMuDWoA4a2pGYbVIp
9v+icJqDQgwXfXqYuzSQ+ErO/rwWMxox2hBcmToyJeiI4gpEeU/dH0mC14l0KiUG4tO4KEEEObem
VuIk8LzbKczVLvo7K1m1+QbPa1ePCl14ay/FlJ6l4EVlLfzo9y8qLlLZYuM5c4AAm8ortZZX3boL
PB+pOQsLJinPAChzIZ12CKtZxJwRM3asHH2Wikz4pkNtK5oUNznl05JmJTuFcbF9wIFLOxhomBIh
XPm+NriKIolyJl/cSlfvGeQ33Sz81R4itBcqeuuHVeqmpBTV08YeUsDrY8SAVIaW2t8wIIXoKxpC
mNLQxNL+aKJnJWDraG3Rzw5nwIHYfsBCYzJ4sM2ji49N4SbJnBRVbmKsyE1OUStDU5upwiqGMQjf
YbtqhRnPa+rRJYtz31VeAGy9x34i6v3Nh2jqLArMG76Jz6Jgc1LIrPSqjSwnjYgiml7x+ZR9h1r/
NS+YMNjFMh2c+AQiKIxgixOKHcR795Dp0EdjqGmStT/zc/eIa4Oa0WOLkre9M+jAPy36BM0GpAUh
8CKqGrpPgbKQvYmbgAmmY2r3RzFFUAfKR7i6FYiGifup15+3XHqNnjN1bZV/XWA3kqGMZD8KBIuO
z8i/PIem8eEo0NImq55NbpQRWbSodvsJdoATT4MZHv2akRJhb0GR10++fKGjHW9IS4MGOC+/0FWP
q2d4zcmQVWPTlEh4q7OPcTq8Pax2Y1hVuaJlggTAkRNdCLzofSpVrFGAOyXIQsSFGwL22UF4WI1q
cwtjmw8czOsZsN7pR9tw5coShW43/d99X2sx6+okJzsgmyXpsrW0SC9coOfuka2USKk9KdfhzNCV
fS5vmiX4Zpq2/Kl7nqlp/GcdV+nDZ+isWEfYciqYf6KH0qx/BIABfhLb9T4w0cAQKzEjhd/x9lWQ
RgOY6T/He3UNC8xyA/ANpBzBP/jHXqy5cRM2wwoOrZBQZPrfTPy6R33tDDF0gU0rd8CxcYnEy/pU
1V6Kznvee4mOCa/3+rY4fwaapHRfi+2cPyG2jhucG96VW/VjDh+vfl4mdRIGNNG6rekCGN3tACu9
L2P2tWNXqIcZFHBb5fDm9i3tYCeliiEIn6LOk4CRSec7uyD+GVne0+QGePZvcG718JfL/3RjQCsF
rMZfrIDl2FSRRilHTAKgezEcmw2DTfEdAgaNFdQAwVYKt0Pgzrj87Zr16E5BbdhVub5t424t4Nqn
8wKDKw5k9I4wKfsukBFRC5vq+TN6OL11F3mCYJj53tti2rH5uiin4mA9LGBuSpkm/8HKru914xE9
h5ZaI8qzY1STJuWFNVy3IwAFVU0/uIaAgOGZiIFzpl7J4IOgF75UZ/n4ObfHpprukM42hEEIPh0p
90A34EXBEB5Hqa4gG0x9yKilmnceZCKqSQ67SziZqgMEz1yhMYlrNrJ990rhAkmSfiGeEd3Lv1Rb
wpYPWLqP6v+MAYvJ+iN3eoWLOnk0b9DD1CuYlCulHZu4BZlLRXaq2c+SnUWO80IQMh25KVle4f1B
UDwHXun7PfrxO1xKEtfL1ShyNysoTXhxy8JkoPqEfrPPvLwSP8rmMtOIqLZEnGqxtUALtyglSRjW
qWeUsCW7OaUVJDxAgrlwMWZGJiGCrt/xE3NJ6Z4uGcbVjblSzbvUDdiC5gBKbz9g+ML/GHAcYNrM
6QPj0zyq00zJ0Ez/g+y1WdNHbWssVLP8K29+nfC6smUyRhaPqghgCZt7Hcl9nogwKx3x1HlnJaLi
9lbaNmH316f4ed8ctChORn3r+oSEdb0AxVzQgQMiKUH2O+Hk2Hfe7tQIh5aCNiNIE7RHtGYWPJ4/
DzzsmajkEyU+KvAG8VZDh90QMCnGRrq1t0er1igBQiVdMEfCRv/35GCXYTxDQHe3iq3FDP/g1ec+
Aa87jXOnp0kSAjEDCZscz9pzmL2ZDFYgKYdCkuTjP3gjYu9PR1XHCFBKMjOTx6MxeSeNTT69PbCu
v9aEOrS9z0bS0P0CVDzIlH1Vh8pv3wvlLILTowEKnI92snosxSoRVQYHQDu7GZxKhm2OJZg+fpGx
uElm4hjPwPLGpw8XwClGr4cyuI2aRAgpEn4JSdFXTp4UpVcJQwBQ+cE2yRuXq9VcqtpbHXV4LZ6+
8+apv67osi31HiK/9T4Du6VuzU69qB5DKZqzIXmyqQI84FWnZsLJQrTXMvibJ/53nH6XbTwZM3Uq
Kmj26Ha5sxGk1MPsu2mYF94L+or/FzhxTTTdDyiUkgP1tItwvK0Hl3UpPWlaQ0yUFUa67CJ4Z+N0
qU/CyLN/5uFgYOnk5Vh9lD0J+0+9D14RuWAKMVQuBacGivlwvSckpMtjqkFhbNU9NJKeIE+tZ7TR
SKSmaQhR3tPRno92f6VWSj1VKwnMxhFwnfr0hDFrbI9xWXDjd931H3KsGuw09Zq4Rhgxgu8Tx5V+
m7v28fvzVptyI6aniNsJ/+zU+UE3vsLVDJFNDGSbKp8Row8+jp5YOZC/Xy2vLgEyflzjpR6euQXX
x81lwB93nyxc3mvoMtadb8I90wNMqjBs2GndDtB2eOtIWQjWE7/wlGaurA1A/1ayUXAey+JzFHR+
o5C44no61dyWsJlQcregaJwbmD9hHD09hgeIghSztBCYvi0rHOgqwrR08S2XwHnEqoVfM7Gzz10L
Txzz+M1VpLVQWxKqjpCFghyObHcEgGCuOfoIV3aN9metYMhuDBFlutjCDU7T7yVxCGKHVdYGGumi
xLE4se1nqpEy9gKukkTgb0IwhHCa2g0yUXUO2he/4BTzIE2zhFM55C97yUB+ZPGPbNMaxmwOMDxo
9HThFxKV/JRuZwibpkVLIRnO+4xF96yd/tHcKgrOXvgmUedtRxvgBliAMoeDuo/+EbZDa9Onnqp1
aJx10sn6eVwHOM/6TueFBP/K9Dq3M994G7p9RLfB6xkZrHy9yTS29w7b+gBBiXbrkWcWwlPhbQHp
k5hv9el26iQSC+GABeSRhgQhDe70GpkVCidPgGVCuO6ZFbPFYzxZG1z6GL4qSDmEWmXGL4oUHbHc
wQGxK4hC6lQiyEE/nrNrVnGztBYiAMeW9sqcvn6nq1UD91XFrJykeaBmybDu5eaAr87hNDeJyZgC
dSKoJvmYgNcFKqOIypbKik1Rhfht9D/rG6yC8XfK6HfkdrYr4fRRP90u69o+8OYufGZHICohXBsR
a+I5lObGv2nZBeyB6Exk2FtiIZGKUUyAVLhN/zx7cKNvU1u3REDdFgO4T3qqAfolcNypztLcP3Cf
aDukDmGsALf59f73E8WCX7+OwOsyzJpUM3Pa7WyLoE0sy2cE+mvseOv8t30Vkp3DA0uK9UOb1kf1
oA5db/3DQ2lZR/uEXPe3tjDypjMrExliPpQFTsquNzKcAUhf/xtrzqzVdversf6AvMiE757WMEZ4
flzvX208ucIBlJbW+sBqzeoJyCzd/uv9jlBHt1R80MqK/cXOjLXajCEhirfevY6kiURr1fJa19Ua
aMZdco+PYCgjxR8Fo3Ck4XgtDUZl4KOXy07zBliHZHaB4ebGt88CqMVI7RfeDOvlw6uqNHrDKXvE
/CXKjDPKmCYpvLjm2ybrBvuVXsYCbHbnxX1X5yX9srmIqUSCui3fJlj9+j83AukL1DauK41KXwhs
XnlVIT77ZGaAkmJV2XmXFWWrHif3jCzZkRA7Nxq0A7XIQKogtcq4wMP/2SuEnic6VRpGbTtrne+s
OtCrQpV22KKsWjXqTgVFqiTGPBbcHXbaWwZt3LNzfJ66sWW1FbAGRYCL58DClZBPVRMVs6UORN1z
GRhTUCLe6bQH0j+fjR5eP9O+yB+NlX6P1bWx9M/bENtpmONrWuDG3AT3l3C+cUHNxTTXJqWhy+ru
WckEe90Bz7U4r+sXEB4RZ2eYz2xSYFLNQdmWFRga9HaNGWaH29MafhVljkh97HawEWN1U0zFWcBn
DcgeH3pKmC3mYVua+6YcGQFsGU62ZiGSv8y1+3SDU1HX3Z2wSxiYllmnixurZ4Sj+NAvqrHhgbOS
B8vs2cb2xFH9Olg3wasJCJ4My3ps5HLryYSwzOK9TD9EcTVbeR/A51mXfJt4E7bZPcf4PVXi8Iuj
RGS8G8aLAVbc+xzn7g2nDm+M0tuEfCnYxmLwYrnrJHru5O0OcdftnUrPIe1UtCC9RgPRZOAo34Iv
NfDppxZL7ZdYhmxs7vmRVwzwb/JraMZ39yj+drIKMRI4+UtfqqEtTnL4XrWGXY3gm5LT7lhZTzuK
9zycxbAlQ5+S8RSBROYv/eH+ePs3m+8aYVdvjm4X3eLRHn3u/CYNY81j2+jIBSP9Te6FB99scpFU
uNZDMN40nvPxwK+A7fEgVIYa/+NzLlw6tq015V2DTJdN+SiB5sXKm2EQ+D8MQb3F2j4Ro5eacj0w
r47yuY94ig3Iidu4a2DboykjKShAR3Pc1fgSasYgTArbQSZ6i/sYBfxRIWMS9KSteIKQOzG/KEk+
r+2kJVONDmdjBG1ByLBIOpvq3X/XyhPUBlWTVjSgqSFghV9CZVNSO1quyVcz+eFPbzJ4MuqV0mHL
/1T1O7zlZW0+fRdI57KFynrbclo08LqmZFKd/7kF1R95CHE+i4pIvND509W0jRS2DBVqw7/gcsoh
DCF9snxotgC8ByEDHwpCG3BH4yB0JSRd2aW7rg7rg1BaAwBrqHjrXv2piRRksDjiXO/CIH1qidY+
nnLIU4Ffq9kfWU3wo0AgwrKXbq4Q3JwgJb1XJCx6bvZvOXp4pNTlesWbAdniRPfhVlBMm0sbQxuS
UTwrvY4cHeHcBvGhN3qZH+1UfrmR/2qksyt+XuioeyIXZ/75B7ZJlIQi0CJJSD3eEivr7yWGUYAz
uv8cSgIZLVGuuJG6Rv9GfxU3ekVaZRGE2bLAZi/n6omzAOlWrRgqXdmkcivXF+4tm0zC7yVIML2O
TyVwBwCIsGhK+mtcLPcOsmYWRZ46+1nlRMMMCDO3FY7nPTqkq6jYrTrfMhKldAgrjRsH72/KN977
CuE2SgSYn+KGPHKKOkW5NxPCfmZ938kHkbw3/Z36tWiEr7FCxHDtOdBtjCp7W2dTQwSPQ2BmxULX
kkMTAUQVnmzhtdK1bAwXEFlXpdrxPCKSjlmfByqSEKu8Gw69kbI/QwY6wtnETjwwiP8kgyeCYNRj
x+5M40RH/7NDoYIhUrEKChuJrI8N1DV+UOnHE3oJqlib7XDR3qIzoVxz694j9EFS4CcBjuRPXzI4
vVAQJucxBETKiZMAF2OKvXPwU3piD9PWvxAJ3MvtdcuWM9vHipA74dZafdq7kCm7N5Q4GfA8ggku
YsqzrZ6bf1FfcDD/hgOsMeT7SnuRpbzKpAGE7JgRIy3+SIHWu/vftCRjVPh+nwQkpfUgPXHqjXi+
h4+c57iKrGGR5vp9jVP+pZ5QAW5F/6oCaIAnCKxaMUp970nzMdulORyg8ViC4NyRR8vwQ0emGJWp
1c7R1/ulk4mqBpBUJYxkyT7QK/PavnB6hZ7wtoebqRKWiRV2EVVZl76h+ij//GrpSrc/vUD+fp4k
99otMoB8NrZgpbKQutdsKxFKM+ggH6jtyolqQU0V9UX89l3HD/ZvdiAjwb9HinT35VQSg+yasmgm
BNBhU0k7Ju+K93FFJR56wgfmzWi2AeAMsGVgJbeoxFJpO37VvI0E8J1FR6kFXYD/9DJuVcQX++zy
rJ1ppaoeuVdjMst/219ngboALPeGwCIJ2rnSdoFl3teqDqycBgxgo3GDuNKB+vgaL8NFFKhgFjqA
3I8eAZdfqEv6JhUnirbLMFkS+F0Ea9woE4toSf1bzcA/s6sh6cxmcz+pbOz1wVqlaXfuP0lOEymA
wcW3n2whFj5mUtAQ8B4AKz4BiRgFC4UuRN3ctqThPhW9hVIKVx1Ye5C1jLwukKHaL1Ol1BIv83zN
MmxGHci4DW87NC+pnry4MXRp9rbp/2rHLKzfhfTXHrUjYHgYZAY+ImVbQiRU6xba5Gz0Mw4zR+Ab
ilylSVJfDJ9tfD7cMRJ/5yDJxQhtH91148cVpHOu8DM7qfmPNX48WjCA6w1T67xYNyjyXPXswrmm
iADT7Lks2e0B7XBvcDp9KX/WtpTgo0hVxFOSuT3xnZdZCl6SyjuWg4D4ImIK7cqu1K1NDsWx91eY
e+jTmY25nrQxa8lJF0p3I6uJhZLwyNmgCQru3EHnHERxdeDNf984hZeN8jSsAu++AL/n8M/sQu4l
FRktc3rsjSOnOeEOdaepJpKJiVpvYda0z9+dIPTy5A2dYoZ7gw9dQQRQOgF09iuYDJGKo2QiI1S/
FEtNA5ta7f3aspWcXDdAoqXxNq83pmOVd3Jqkn02oYf4Ue702YOkuUAByoXVRAFerkNMzCQ7U1Ri
QQfux0wd5TjKwQ3bONqglFzDkuFi6M5NSG+98D42sWOo/otn1UdRnpo6hUi3mwvh4c/4XG/jFYzw
HA8wFHONgl4Fw6+4ATsKqz+F4DmdGcHN0p8WZGV9iJ09/YByLqG1KERlipz7eKIC39KvoziwOrHo
o4vsCRSKn7nEiQnX87eECcI1uyb5Jh+/F2lryW89VkK9+eInJ8CqfxBOJUR1INBKrWFoL1GHzd0o
ECQE2tPW0IU8CV2r70InWjHxX8bQ9yN8j89R9LEyfMrrqSRofpa49jR1exty2qL3GDXxVIzET4UM
cLHW0vyaa+CLgpKfwTDjWKMu1jy+dK92NWA6K/cncQD1G6UvBuMQs3u/q56UXiwyT/ordl36dd4D
ZWdq3HIH82kzgntFMSLPW19EkzCTSVvacdPc/Ja+y9dbkcD5g3U9V+TxmJXHGWWbc3JOjlR+pr2O
iVYbTN6O7/kH1MEW7QKtVj6UcJNaRPfmEI10VBlqdpKkYWN+NZlESU8hIS4Ah1k2w5L6UFJWPhbM
HLO1rT1Gk4TjVqYWYnnr8LlR2YRoB7/6oeQAgI838rZ3Qc3yG9flVQ6meFTOPq5kUnvs1pMVGl6S
7Q4T/wBW0+dj3Gr3f5r72F8VVIbfnAa3LU1nzGOZJEHKj2L5vU/rihud3tPBx0eBUnBR7tInwH25
BpSwqp6FOdW3fut1YkgOAAsvLDPoOjuECg6gWdrHSZfh/FT0GA4U6AwY94snQlzItmGC41cDyYDt
vyS5GRF1I1eQS4t8Hm0U95y54aYaffrULIjt9npPL9dMiBDgjbQAgYn4fmdarNWmXqScmLuLTj6h
N4D7SsrxU0yF0nlDOcS6OyrSHDHX8ws6zdx8DgntaumI/pekCycVGsBlp33Y+tcYV5x9YhVmIP9d
XLgwxD7MGy4OdPNTJ2RmDVsr6rIaqQzsqxrnt4HFtHmxzXatUNq3sM4tryoshv7C2HY0mEhnlAR3
8lzK5/X0k10NaPZPNc892wXOsvu6nGuggxvHrxXUwR2rxW0e3JILKA823MA/hPGx8qavk4nV/9pz
G0kWN9uk8mLSWnYBLG1MBynGM6iDVshu9G76AJX8H94lk8cCMuU2/PMdA9jkKv/YTaUjBjJPofWM
CIU1MbS3ytidYDuCL3Jsdt/bxo6LPA4uPwgwMqOHn/BkNo7BwDsPXILokHXzZlswBAEUfzzvxFlT
ORqILoFbKtRy4+ybfdxDKTJdIjON9YuRoznwc8AZKxjAHIxxaWgP4pUiGnHSrd6WcesuvEPeFXqn
2oFvb/k0Zxq37IXTzi1TB6MMrFgSvASq3T/DmfGvANzEuC9IgRM6u+wlNVqJfLmleSg741y7Zf5L
oRSiy0RJkUK9acHoLom9T4YNoD+KrdvBN6tB/Jt8wf8PpdYi2M+KQyMq2cRuwGNdDrw27YLCrt1P
gqEf8pwMO9xth6jRd3nWXpQObMe4TZzwKiI2UdTq2ZCLaj4DpTXr1SiPxxW0CwDaQJBe9HjAafpG
9qdR07fLbO+71kiV4YXdjfrul8F+BXGLV+m1gz719AG4Q4JZctFG17Sy3dIYd4IRMDDNO5sHjoob
/YS3hyPjKkS8p6x0bMte4jv5UaImb0GWjrhjzcrwxhMUMvHTi6dpWDjAqmBk/pXf9B9zAM+GsLVC
HA2mvNV1u6tQpxG3Sa+t20wpeXnjDjzWWKqD5sveWv7VFbavsyqsa23c0jMu7F/jzXiLs96as781
m+b08Oel0ECuZoL1cJ7kz4+3pupXO4AJblZnnw7QDp08foI/j9bZ0ppotMWnkALUdmTIJS018D3e
DEt+TOWwES58kLIuMjDI9EkjQwJaY2G8pLlY0o+zthojFTfst244bDgFnNlokPDiUE7AaTEXkKpG
n4X1HPdC0gEQytRWh1cW18PxFcmU/v7YJfAzDBbUVgaR0Ryw+JGPK/idZx7nagGhNw/ExSdFES98
PyxPtt8uV6rNm4uiP7jjW++ivONYf43DswIEXK3UEB2Mu/dY6Sg/IazIRW1dnpdQV7S44Bw5omUV
x5Hw4v+34WKGhTZhNXR2p7ObCqfes9ZaO1cb9rn0rKbhgC0piWmpaXhDZoF07nzKxVYFhozbEi19
RII8iBNyBXDVZJNkGfsYJwuAq+uAocwiGvW7rUrlldVrbhtowiZoWwmMBrihk9FqBx/AFVqnBlQQ
BsKjSXbPIfkJaomF5b44r4jPBgSSoRqM9OVEXBjrfujAvSv7HFWfOVTzMoFcuvt3X7RRigfR2Es9
uztYyrgKoLXjeDVswlPAAa7O9WXM+0p2Wyh0dpHcX+RI6MWJHOVj6l8OUqkmnS4g/mOGbgjalSdE
sqJBGx0y7rm3hI+DIx2FrUcKcdd0Aww2IEsg2F7huD7EuI+JMzJMaubE2XiNZv0M5G1L95CwiZuG
80wCXkhnFnFWdewAqq9dujo4v6wBKTZA7LuAE7Hq7AQcE2MVZcoESRrsqe49gPT4P8602GL8jHF8
fuXCfSRdr2GKKt6E6+VFbz0AauNy4hiY0tONHL1iSLMW89WvN8XqOyxyi12kVsJDtwB2YXmwl9fY
FD37BsmkeLPzcgn+k+/GT2X/xwiWn0mAONfP5h2V5l5TsoGoJa2hBiLPtv17gPGbN3BDKiet5fcB
n1NAuNd7fulbfCYtPdLJ2npGBKclr1CV9m42Of3f9lrYjWvDjZ8aW3TzNwLmsix3plONN9PxwZUK
6B6FXYZFwHQXTwkmJHoEVjZu1W8ncsMvETsGAHuYwguZfs4jet+TPiLYg7vv6QxnOx8t08svYDur
DGHvD/PfkzUa6oiUFZWwZ7yz7IV3DecqU9tX401hQ1b8RnsFJekOzKf/TTQEyudDta2ffGImPN5i
bnFjLYoCbY95cZFaq/Mx+GvwcVdWSjSVbRheD1kHCqvBCNwgb6C5dpnOXtt14q4fFumrqoTK4Lk2
DH8iy88+9XuWaPVB20Dygv/bo4NolCRGWuzDkQJ33jaVl+OYWE948chjNZU9DqGckXPdce3tcfKL
Y+x5eTcmqhEe0CD7FwcxIC9fu5oOPyqr8El35/vvQ1WL+YXmxnCX4WUpACDkNOJI0BLOnv45ALok
b8N7z9KC1Wo1Uw1A6l+G59h+eRUDSDlWJdhYPtBizVZT8So2YxCuwkVm2YaM28T3wYCPhEDLHpst
euSLvFl0s07ZLnzFELfzgIFZeDbu+pD6rxwWyp6vQRS3XwBAnl/OSHPQ6ykR8IGyEwQQ5ko8867x
pmhQFyaJEsuIMmIcw9E3WIWwaCMkmN18vVcMOTUsxuZDoI4RlRXAVM3pfCXyRONQGoCEUs0NCQE+
ZHhT5Kjwp45EVeeT0k5nsg/l6ot/pKIGc6sBaOSlVcl5XEvAUCDGabsO5nhUVyZL2L8SGGlnkdbS
TPkoJQPa0QNZ7owcWVqZqQA2vHz5iedwO2jmDYaPZx/tYM9XI6N+qAkAqItrfZGTj9PEGT7uY3GF
2Q8Bh7BAgkHIiNqLndZBOWaxFpVGEJIT/vmyaWyNcXKi4sNKqHYGnJcN711+L8sUpOf2t9U4NAIs
wwT0USDzhhP274ZFez4YgOXVzmUYcTobwgiEg2UnXFm7Ht55MXOLXoimkK8VRFAN2M+STeFbNkFy
upcuHPAw6kNPhzp3boNjV01DSVmNJTnO/rNmksbhB6s4hB4AvsSJfOIH2T4j57SU0dCIdu5cs+b4
/oQ3KL1G8XYzwMNxCsjDqv1Yxu1uMeusf8FQGnyEkOYSzdm0YBF7vaxe3PFUlg3T4Far57OanBFm
3T+aob/+TrFYM8qFPVOQxcok4qfgwFbbWTPQouM4GoQZTd58BX1QzGe7OBE5QALcPodIYGXeAC7z
wVPwRH+371t+xM+77sCdsxpsrDkCw0wqta5KELGCe0nQIzqxkkHk1tNxRN8Urs0txLdhF4AVeK+3
ShMMgo4obgi1nGKtfDoSXmKvHE3uZdkHH3NvENqIrV5MRAMso/2BmhWFtiUqgbMO/wwyxv7DDsto
8u3h/6Kd7hHkCstdQ5b1zThsp2ssVeywUFokOJleZw0QW6pum4RwoyZ4eyun4LjSaToPPA3WJOCi
jqSVU1hnGEdyG5LCBkDQW96aNHjngVgEysA4Kif0RIw2rDnAIQ2k2NL7Ufq9RChGO43uQ3VSNSIw
6El5mmt6NY3Zan+Xyj8le3HZCGB+9ccMauXNW+mTFV1VzSq5I8aAsULNYf9+37cDjLsFtxCOVrAw
LqB4el6ikh4du0MJ6CRA4ylNRBZawRry0JN6fV14mJiNckIhFayrmSPwqWdZUhNT2Lo+LG0MjRmK
0QG885NoyWJq9KN9T0qtnURGH8FyqymtwSDSgoD0EMT8S3eEXT/cPP7QOm1xpH5GdEroL37lqE94
pF4XQZyEcqq/bYxyFPVcMZ54/MsK73zI5l8YRLXsd9JHUnQZtEWa6OPqy8c+6aU/EI1qfcXeZ62m
A0yCKr4U3OL3sXyWm3lWM1NFRPX0Gwk8BuV/BQPc0zd38+741nnQnf4SiTIg8xzlMeDE1B00X0j8
IS8HHXSZ4FKit+s3KU2aKqD5CYdD99WqwGwGcN8vzOogh5AAQqc8i0pe/04AAf6+jzV7BFMZ7NqS
QgBvxn3s0oYuRfXq2pVwR7Vm4OvlQLIPg4hfikOrwaxLrLuhYvwMBX/LM9gbkfw3lmPEp4Tw7SWQ
gpW0AcnBw+2vOBvJADnVleSvqmwP54ojfej1DOcfq8MKTAlmX5SX0T7ucm8Q3q031Oat/eWJhWMF
/azNfRJHQ+u/dRMorkusGbFR0sI1FiuWImiXyYsta6gW+A9EBTVJ+d/0eTbRpcUNmmQ6Utb/qXWd
URaG1NQ1JJWW8Ojd1teTPAuhLYGv6wJpywpIXiFjhyYZHf8OLrH9vWvnxZ+6yvJ7Df5K6nSBPTH9
8PV9oSHltzNxZtR1FkXiLg9T2kAzhgNsMNdJuXmkspqGj5QB/1qxVWcUvCBkxdxk3u0LLgcNNhh2
GrzGKtpKXhvnC5ASpJbeOMclWJ26kdxRXA3Ws+e0g/GOwmQ7BZUw/14wz3m4rKkvxDBLZ+A6/ZV3
brCysJjQ4hb0Q6YVIjirT7S25OUztB0yo5Yijqh4YjT1L34B0jx3xXzUga545pZiyazb5eDH+sq+
xt3aOnqjWtmPO9LBZo1JBeORUS5CRSisUQmHv2SrNXxWVB+9vSvFJFVieOtqnE7z6gQa4thQqo5A
Bx554jPYhACWgw+wlu402FkQ7v/stQhomOcx0qyIrMOcdtbI+07ept8J09s7vd8Dvgt7ilHKNgLB
nBeGpQbCdfBoNwuPMIPhWXx2MvUUc2/6voiVEm+JPVY+5jtL9+Ek8MLB6hjuDJG6sMJr8vIFdZDm
5kbnYnfd90NfAop85EyGnSvQR9tdDdoEs5aY75yxiW232WvcF/ArppNB5RynDqZj1YC1FtK9cYer
3trb7UgSjhf/Nci30isFA9Wg0u3NcGvC4GGxdZcdwGkF+ORB0JQdKcdBsff+Hbh8wZ9KtslAjf8K
ggHSdr4FNNk3BH8uB1aeCbzMp+fOSNKq0NPNOTcK8zDRNxDnD13ZjgOzsrzHyPsFyufsXR2BBY9a
r5Lnphsp/ETfjA2Rj8ZXycdIfbi6xKsP2Brts4gJvPkcVdcYlfHB93hHfyctcISMU0ebfrcpOFVd
Lvvslv+Y9uk6o4iWweoatVlfI+Pn0fMcMxgLhGKM3u4Zy/qXSWzMfneEJYn25I+AfEjqbpU5amVl
3R3/Sg0syYVeApjhLBLIrcOSj9V/3KCbKeIC95kS2Ywg2+bMfoXQ8eb2Nz8rQYy2NxfO7irBiAuh
Upza8WdJYDKr4ZBuDhtd4rjWiG5iVNTG8hUzvKSXlxy8Rx8ObRVnoVff4nfqwGtYP81xWvQOWXtj
DV5aY6X8hknuy1mbDHxAGB4mfJF1VtmlxSmscqOKCrb1O7cij5yOdJaaWmN0MAWFBoptbPnZScHO
yYl7Qb7oG5QvEPZerzCc0CAb+wI6DgQWRUxKPjG6uV9RxEPVXGDxv2J3uPShc5aYzwtScVrQ75+5
1USXVnQPs8LKrFGaMzIsrUZLSl8AQ75IJkocbR8CM7uOmWalZhnIpvsBtrsb17p2bjSh6THBIbMX
Z2gR687naaEtTUPU+APU5NA28VRtRwf5PjsQKvA61Y3IIY+B9s1WrXtVvPOdgsc+gt+tCN/Vxnz6
eDinzeEsxKUuXTxr0bLJzumo//Ls6elVS/oHGt0Qdvwb4HM/+05+KgjSQkHFcIu0VwMoeRSadIRT
lyNLGbdmKjxoo9bKP3CX4p96zGayWnBCMjeutGPSELpT6NZI2tFcfTQjZzJijQpFy/EYt5Qj9jDT
bFw3gJJR5oQ//LVEEJGlFck/dUjsHXSetrkL5Z7fZwpA0XUcguz0DdGyCT2pDzbqrJfajNSDUYxr
H0Ivhob6Yt5wkqPazt5qlFbFt4KvMc7seShKmxZZOXYrj/bodJqaLpgA5USAlB1TcnQ2/y0r4XD3
L8unUrOllLFQi7PPgjEpRsUcgPqR/5buRXmfECPu/mP8ok02kbSW44Hsvsbjm2m4JCwPW5b92Seg
ni2Xm0fi1N6UjqKvuSUGMei4ODTdFpTI9fZKJJQ8qMl7ubVEfcvikoVpUdYfzjXHpyQlAvZd4abq
xXT12gUjeVLKfrV872t1DMiLLCnb0yYd8ZUkrhawB87dGUNLS7UPupivIm3/pcFgIgVNGWb5hF/a
m6cHS82O8AaaOAo55oAYSEGzRQ0eHl6a2gPDFGNReQyaH0z1EMN89P0SIBmssC2m8fAT4yrbQ7Zr
vdFWLtwjThJnqbbEVqIP5E9ifsBcE1YcYAcxDky+tokY28zhIWgNqDaCW3sAEJYLRx4t2rq/MgVo
0qXppK3w2RnW4fmopJBO871YHk6jS4l43+wcrGmM/4uL9xHDAtvw1u5vnne9tHD3Rs4UxjCbZdq9
508P4oDdn7pU4MJR3vjchh3L1fGy9OcmT3/wAARGT2QiPJ8esXC++cbrbrKbJq4LsTEkJUpeFKH4
T5nuVpv8HkSP9ftkYbKVpAlZYfYgI41WC2RZNxCfSXC8MlJbcyICRq3uH9WyFzaHBSaC1TdnS9hf
yjWrHF2GUSvRvFUwFbpEJC3pG0oaEX+RK5Aq30+JJsW/xVlQipAAUtaVNO74YrxuU5+rlpuaXUBo
dtlITp02DWZTuFTaF42NOJQLgMg2Leqvo7YSaqrAuQf3TWT+1J0xG97iuMUy6ctjNjNk75vwywEa
BzIwYl5RLNQYewmFGrv0GX6uN/uGsKMNaQM/ckJpbJrG+1xRzB1BKvuSHm2Ox6OLfoMQjenYk9Ax
hsWjQCo8ozzYzzsjgYkhSvv2w47RQK4CsiSoIxlBJR9kLxQfCyfVNwjKTwZi0TgHP97BvHOIDdB/
nOXamylB1nAII/sCEejTlAF3hYyn1Xq5mZqi2K0iSKkyA3n7VUVWWjHsUgDk12K+IvNgfpi9dpBN
mmh4L9jeVKGJRep89CbBE463NKkzgYGxBo2uvuyyES3QgSsbS9wBnWp6XQeYCb0pPhxTWUKiFcHi
texe2Sx8lbqHzeJv9LTFfCPMbrqRP9NZ2+mErY7Yg68O0h1klCDQn+09sbNvIe3lsbSSd81nddlF
psR4TKUPYK0V7342tP8J/Cr0Y8pKoEoIWOfsokbuZaAP+YcjfKnQkM25Z5gKCdlnQBSz+Egoq1+i
iH3LOJQPvG5zwqyuQvf371K00wLcTDw1d+1VEQWJtV84/FqWxE662j44BU0wi7eZAP71AsIiT+MW
Mob9FS9/eGNQGHkKr2ymmOJcCTE4+g6mTr12R/XFvy/1jZMMPde6ydxlAhF2MRCzhqjUOKSpvmw5
A3R2h++61JZ6+NY7IHzZIMigQjfiqcFeTbHowJ254kd7NFJUjDZLzUOh195C4FGNlyMPfqThvnDN
SmVSUphG6+oSlMJKKb/9LT1Zj3W5tEGl1GwMsQdfyxR6M+5ycCYz+9uzKX6hiErfY2EVBnOgAan6
YB5yhzfOkxMhAhWbd/u4T0BL5RjbWl52Bbhg/N9EItLYUtrRrqw3GPei15opxiH+lMLu1jcXgLIx
QOWNFXslzx51inQVI3Uol6Iw6Wll3Xt2A8cOGYAKDoEFsX7hs35noOfBr0OA6DxHN1XxWK1L53Oo
sZ/b4ScOI9jFMDS67T3rE86ebCanKs+F0hYBTyj5u6jYPhTAE1UxA8/veZY471P71h7jMU7Mp5iE
LOV75K05NPkoGZvSi2+xwAiCMRfI4LhE+sqwvheyujlwFw4+/Lh0DXJHFvMBFEKTmRNXAqhUHvdg
QQoK1FFukMEeBp37WBEcwDRV4r54PM07YS520n/Nu4ExxLrXFe5Q4E25jKP7Y/p5QdGWKtxIW2z4
YQL/mYGb35bhu/fuP3QL5AbDgq5pxrlvvYrxb0MPYOsWi+gMk1coxgnAgN8L+cDBlnBVEvByEPqT
ycrj1BGtx3SsxI8XAYy1ALJoB6ckZ/71QwofQ/bbCpwJFSK2lt18tAc+ZHYPpJBflnFjb53fdGFa
7PioIEpvamwkhX5LbMpcxSdxCNbtue+wp+iIGpnnv+/nGQVsRiZ41DXCKtbTF+Z6KeeFtOe6mnbO
H3MFOLeNRlnr2TiTHsL7M/N8irfX9tbSuEXmrjfn24d03eV9xDWa0Cvqv6zL8AejiBshFksuOYwD
XjPRNEMiYtlp0MCunio9O666v0Fic7aYJQd5cHsR4hcyyEeYG0eao0CJXWJp/4aBC8SnzSd8Weoo
KBgUcm06LH8yttwYssZIwI+FgJAZMz6II/ohIgKf6a6B//XlIIe2vCAQ7fyKJ5AT4FBZshW2kO/A
XdEko0WlDqXiqUBkMD7HOos3a7zMh5+vlFAlhzV64Af2MDlNnMJm2YYc9Ok9kx/PBVcEbNIQC3JD
Bz+h/LbCol8CWjl2yYZai2fffaL8NZwLdzudlqYJJ42pCTeUp5vqMSeQ8T03OxX31Ch1cNXkWxgN
q27SBSm7Ghqrz8zxB9PzXo34ry4Zz3mk4F+VANBnEqYa7rsJGRXlGFsxpp1sriIW0kb2t2mDvZuQ
MEvhKFoUT9SNHNY7/bffwy8igL4cWjfYhqM9vzvl4Z0KV9OHhcBfTAceNtCESGvhR1Gjka/KwWan
bGyxUTSWf9zd0d5WQzphpgaMyIXvLtJFG6OCbFFtoGmcorszGYKnq0YE3gdK1+Qa6cnUOEiS5TXV
Y7XKMMMXHeYohuA1QVsHuMQ7I/GGOeUsYBVHdO+LbuUk32jBirsaE1wKXwX4WY+eyVoD+DIWdn4i
ZEzQGYjZfAGXzMLYoyCBQy+xbGs1LUgCzenxezbENnW+RLpwqOZSIZFT/S2A77iYu+UsbBsym9nI
tTf+O+O70xGAIu7MtfrIp69PLoGOmmWAupMkFkY/2cKY8Ds4ukUT8XJVPdyrifRTZJ/QwfnVxPvi
5YuyGSxmJP43w2yl8yNTtCrtoDfZRQ0Hg4Jinei0dsVDyUfv4MX8n3VUEQiL3kEiOEMXZTacYiYw
5qI2GsJXabBOZjntqn8CbDlXposUhaVj7i3r3geLgwjUz2xWUHJRWmnPcwNLHnOqARHdd4sxxxoF
vAjCukolXnyrLBm/8Av/BpUNncDIyaX8Zsl+ZFVcmhL2dqHrKSZTvhglNHUTdcvXe1JS0C8AaYqw
9esA+33ivZWB4cYR6c47zYhb7hSWWbUACwUSS+ldDLM+3zmdGcmTPGCVC5Dw3UeFF623n76o5PQU
6/VTXi+V+lmafvOOC6vPju0kyHCVXGcvyJyWtrK3IRY6nSTUgfQs7sDN4oO2a5PbKCBpkYdRJsWj
NpcmZOcdOMm0IhUrEtxKSPGWSWiRXfcr36Zme2x7uQurPpQL0OtkXnd+4+SLJ64Y6NedVxrz9D5Z
9n0HfKA2tzW2oqeN6EY82KjeOQ+9Kd5yOxotnDnheYCXh2h/BL0yfrjLkIu71Ra1jSPTJub2l1YI
7PEMnVWCBIYU0ilKQg7w02jHFDhBLLFIhTN1S7MqfzihOo4Tq+FGNVggaSXfAbczsjwy/kE3QE6N
vwzDk6+oWaHZgh3R4kzH7dsq5UjZbhkhDkfg2QAVcPGXpRHpDTxSLgmVLkSALvO5Tcjzf8GoH6rm
efbbY1F9wqOCpkCmgdLyPpLx4AJZ9u6TEdQf1T7plFzog06mjcJdolRlEfA4wJYOPVWn9UrtcMWU
BISBEytdtE5cwJVcDYy0w6X+SyVvvrPO38MLlIevf1+lSAYnoQTUYRTMD6zUEkmSBFoj3WbJ5d0h
3GfhVZUSqW9BOAC/722zVSRE3aUkzm/FQXY5ZaqeFltX41w0CW4Y2RISvVE89nUVacnsSGfN7kek
l89/YPKA39qoybGgKvnjf4UkEa/PkW636wSgR1nA6ApeoGpKC/n6tiRKD8vThQfj1VV5LYg+xx6J
xosJLnxaBq6DwfrkBD/o5r4z17YT1ox9qIXYP5eRmY36w4Xt7BHZFbFE47KaVbfGFjGWoxUvbZNT
/qGOoF8KB6UmsoWxYDEtp4+YqVC1LfIM0zfIF5qShTxP41Qd/asj8OWNauO6sDGRsiyXQtqAByW9
cRdMkza4amCxeDCHT5/9X5HjaJnExUsyaW4iWgqRLNCsoclsq+Y/2LyGZTmADkhYvQJe6Hy01qYw
RofnG7lYMBjEJCACvECxm8lbVz1w35mHEHOo0NwLWGxFabeLklR3nHSgP4nXUtIrJZGkta/lB8c9
AXVCqmyl7OGPO0l+Fow0kijy2yChZOt3Af13wsR78wvuL6anS/k5jq/UzxtIzaqC88dr1P5DmqWt
jpHbBSEcpS/4lIBfNtTH2pgf6SGzkID/0do0q6I29WrqeR5VFhwHYW47j7N+71959/8P9S+4CKG+
gjRlRVz5ethoj1ndkxY9cOistUB9vMAOfrn6ysKwzjTbEnhuMCrfmHH2CtusxTyPjV4MQlIZbKbY
OwfKoLMNnZIdsJIDKs/gxQGc0a9M/sfZgkOqAvAS8piUbCcwLx4NKHZQznawADEzk6VF9DJnHOPY
b4HsipxJZeei35qG1xF7/88TlbDP5Q9m3v8F7s4YywCQFB5EBuLN5L6fmG/68DKyIqOcdJsRlaW0
PKoypljcJxBG7fS+VayItWNYFglCdGROT0VQJUie8gUxdHdQyDDNBb5LJ0cTMq09tOb9/Zoz8QOg
2qWHMWI2PWeYJCaGZTvHjvx1UnT2zMMV/Eoz6+yLnoWo/GUxjh5QcLN+xON3Tx/58mHtH9alpVI4
cd5S2050h5wuN/c6URIoKK5Gv7ewwl+Ow4c8ZJfjsfM/4QDmqSuGn7aAUY+knFy7aicTHYW3Tcw8
WeUOK4ujOXNGntJKyeY1PLnrEVIrJZyX0da8yMNDhKAvvU4v0rPzFZfMA8vRvs0zhIKM5NdBxBdl
tI0ALnnyvDLoy11dAzz0BpED8buZlUeqoYmRpwzgh/MyvV/3ft/DMmRr6IEroN/Guj9+jbN9HZ08
S8JI9kAk
`protect end_protected
