`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kjl2K2RYtlW/tH/p9qU6nWfvXCPC8rH0AyjOrfdCktuiMUu/eJ6vjas/6jPXgnRM/O1N/k84ZIETdpYirG9NhQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OkSm7uWPyCnElDIacFBushCpTvDB0KtVE8fHLrkF19yIn9bS/ZRMkngEhSDK08DUxxSh4QIoD9SewcbC9lSkzUWmO6yg1M6GiUsmlv9BsIDFUH4D2SlfEgcZLkLJC/TqYqFt872j9HrwD+iea743KSiNzIiT/w3ImW8CAUtw1VE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kVVhZEI5Tt9SNC6L2ZrvhFXA83jYXPHomQ+u3TuRFFuzRqWVmi4iLvDqx4lfxFfrrBwHyNC9dgbemQs8DcRgGLyBlMDG/Ni3yA+THiPQ+JuaQMzs4loxnr3B9k0LelGno+0j3Vf8RoWaEHcMzKdltZViGS6wbHytI/ZrefiWMMpAnbhWThGtoLrzkIxky4uLa/z+ycsu0pOntVNINvX6csOWVoMUv4NE5hPzLwMqD9TQUeda8vxMSe6K3mxdLs9Gl4VaAhHny8Pqfw3FnHGIdktzBu/yTjFNGMdL7pwR+JYOogKJTOO1/QPZvb2XY3E/fVH5DgseFPNSQff5tMTQ/Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MHoQqG6VrEMnQe7aVeoV72LVc0222HatINdmzUecaFjT8AdBiMdXTKew5inzQHyLJ/WAvbJNVTkCNsJNqrzLcarJKusL2PAqfrOnac2zBtNSBZdM3ztWdsqMoggG39GTmUcVf+LLOjQbzjZhYaXziRjyZMVghsV4O4rE95GacCg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z+Z1roBl3KLH7QNAZvxyjXw1uKpE32+glE8gqkmLXV/NUGG68eB6SpNejXqpoL0arO2K3/MsLBSqcsbYjwd2OyKrLUItcEXe/xzl/WiMnUuGfkfbvjLjPZwqI2qw8grqiefkjAStJBGAbQVIXAzNyo5/yZizoUa8qraFkJQfSHK5wiaATwfqBvYcbO1q3gRf/jZ34iLGdkjjkHRTjk5b9r/EPt8DmbnstQSzecmPQ26P+/6EVW4NzgeZV6vfm5VehaJApaR+BL87aP0mQHnqDOG/D2b/vdbYkXEPASVvsYWs4KfpE9FvfwDWCEZz+nsUZBPQovy6A67UAlYF78AQqQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 169698)
`protect data_block
73CE4b9MRcobXbeUclfYZb7/xrGfb0aRBtkMMo/5BEOLrx3/KDDMkpSCH79/o5I/XdKtdZHeHSYl
hO/AUxbxEqyyYKAufDECZ4DROBm/N5dUFqE6s48ytFVaszPxM2mW/PHJM37jrqR+cF2wf/r5kEDq
7JDX0Z71MNcu+RHUPhwKgN7ylkrjn1lXdrdjLtYciIPjoIQojVnvyT9E92osiQvjbcsEBSrNdi/x
ldwLQc1Qpkz4DRm/Db3AQVKNsTE4qrPR9t95YSLZwkSZj1I//6Pp8Pir9hyGAipph3b2r7SoUcO/
/VYC//4PGwZsJHTc+rJj7EcmNGhRKVtcZ2fy+LEtgXp8zkTpxenweQt74Wx87GaHE+HrZT4VCccV
LfFiWaM5Iz8CcrG8EkV1peag0oJJbYQeBuV5vVj8ydaANVjCx1iVW9Ykeo8q+T3KDilVB6ke/tro
K4I/qtxg0L+5bFGtYxTQnMdAF7YEKbc4caglf9VngXJuviG7b6kX3LXuYKGOTZSeKCVzOnt7g+p/
HZXISU8xMj+302uzxPE/rEqgVZdaqgP0yN1OwBTt8oj58IvBpQ4kH63MyHfOG5QtKyiAbaBca9T1
6YqJ5mgLRA0FpNluan8nKYv/dj/cFwuWGb7IXrm30tWqcFcnXulxlDJGzQuNfDBKXcRa82XUCT4e
rY3qZE0XiCC0bE/ZwDRdqfwl8iJwA9kG3HYsV+/hKQG3Xu8R3a1YE1amGfZAl4hZbkmQA0eXmexA
Z6XowkvTVeRdBhCaRx7I+q+Wvqm+D74ih4kCYQ3T86CAbg0SfJ4tMiHCiFIiRv/yqeioORfMcyIO
K7h8LB8A8o5Z9py7wPGc8cCa2Ua6t1DFXMRk+pnTINLv/u5DkxE8DbZJ75em46a8/qTd17FOcEjO
V2LaFUXENl6Js8/WwIF8N7gNmupSAO1dyT+xJo4sLTu6GSDn5obhLdAtCpSQTUW2PgalUsTvrOOH
ehzwMWt1ca9DMjH01x96OYppNx3FSZMZPG5NIbm24SfLWGVBm7wW/zm0y+OwyLu6nDLnLDpjwIKv
5DsHQg2Y5bSkg5B26CqZMfSzEcLnieV43zA/Q0BXW+qDkIQii3obNa5k4MIBMvrLTV/GUkfnWJSm
07rshWu+F8hHghVTTcbtNfqzktfkRgi/b/vVtCHBKdvXXoEPwb9KV1gVUEfG/Vvshht+AGhakyN3
H5WglT14vbBwEC423Z9aoeTtta9S6T6wh7gCZMopbFWjctkk9DeXLqkNz8WtVVyk8Acvh959sXeK
rBjf34N+Io7RPt6xg80q+Ium5Ri2Bbv/ck7rGsnIV3DwmpFBGlYgoXmsgYJbnSZ0DGNG4OLYhw7z
ooICuhoSy3qAuzeLAZYOGlene/Gd3caXqs+Q3f9ug1xPsM/ZXHRhYRhNHMbaxM0nT2s9b/13Nve7
Nv+0BCuGGRAYvu3pMtmLrvojVBxihnyYS556g1EWQKUc1/RCUqiFC/3LrFJrA3qmm7yK5D4iLrL0
YuNWT3nOOM6kgw3YHttO1mYwL6OIjyj0s//8krGN/7qNmxaH1TFBuW/WAhw54xW2GE0mkhlGzvt8
eD+a/JbwlqEoZPBX9PXci1by1OCavYUweZe+LHIOhrnaqzynxAnJwCycO8wqzbXKJdtb0Er9fTRL
GQcTPosa7dsYC8xS5ezbqK9E/naVFdar6Tma/kzhLnKDeKsrV+tmBopmxXmvUlio70TaHKRlrAJM
F35QMwcDgKG+cv5XOzpK3Fb4rulHheE9YHMikI/DXWlsPiRZQFiHTdKyTP7eOsqHiD3jGJ5jR1wL
unP6wtNEIwEfs28sjVBQBFkHbU5Ld4B16IwYp2e0FImVDcHinkY62OGrKolff7aGWhscK5ekomhu
Yem4FhnlMmEURczYGfDlRKIL/9d0mvY1AjECHm30LZqykefFv7eil7SDQ7aOnUm79Yj0GS2LjoMC
JiljUQ+0JQejiyiPQo8XLdRj8POeSDnP68hZntjFo4M1RSClwXX3BjRDE7ylGQ8kyO9Srg3T75EP
WAunz4r3H+TpF4FhbVrPTK6Og6nE2+Na0FtPoTfghu0Ot5xkw+cKDbwJBpbYnvDSz/zfckcSs4Lu
KGBP2eembYaOt75+oP4kpMWXzSvv76k68+EHhunZFHcK0lBvWq5BJg1NHN54h6eLbivKtESL9Pqi
zDwgaZy3rDVHRXCk+/obmtr8dkRV6syEops5WS6XzCYAwWSKmCSvxJr+oSriNSNynH4THZqc6ZFR
2UKVGdlL3PJuYWwqMU1Atfo8bjyCLcJPYfxXc9zBZdIjOJLuhxIWYrQcQ+KZz8KyvmkQM5LZH4um
Id3HlaYxAoAP7VDI0Sr/Mt81kbH9xdqJrlITLIIfoiKbQWIas4sYqOnslPpSgXXx7U2JVR6jmNrv
u+L8+HEUO2Mt+YkbKPiyd3jTdabQN/vHdd511gXsqxl64vIkijxq3llNJbyyZ2NhV2Sg4t8lPXgg
vosCGBEdTQvMJov2yVav/uJrZcdkqo743McCC6Eni6o8IHB83uUGlHW9HsHbLPAb2nwjajD6u5Qd
NMfxbLJAzMH7TIqufTW8+38cyoC8LaZ8JkSu7tahvjbfzUrygwA9/s+lJ3VByTKyqEEY6iG+U7TN
K+BOWExswiEjDGpDRK2ObMjl6gbAx9BZUooVA5lxm6QQ6qN+ot6tG4IgKUqmN6lWL6YxY9One27H
YCGaVK/cDr1oTeaPiGs3oyxg4VqcodzBdcSctSnd2XbKjb0cUuMTRLwg5f3m0BwUqwBGzI562ubC
8EMMh1Ld+G1cD0zgB3sM1qskz+l0P/NMFCX1YR7zzTLwRLnKAAs0a+gN8Z1gFktKg0thRhFbGeXY
oBsfSGDuYt77CyYMzYWKAKjBrZ2p8yn1/C6QHKcvibFd/Xj9dy5AZM3zvBG6+Qh2s8FhF+as0jGW
1OSF2PzlVpuyme9xfQBGkOaAeTaPXjLShp58TxHnSEY5MNeeZPZ17HPKxibHfWjj+WMOzH1GGRpF
Dx3LGY9jIlZIxiphB1fi47E0elXwIrtmHzySeyePhaO0ifICI7kjeNsuVbfp8V10AQ+64O4+o5/g
I3u+h4oDqDI+katY9cPAvs01hG6I/76LmZUwYKaNvMKNpnEnJ+6Z4ESCJGOdCscafxUY8WNl5Kfy
JPDF0H/rrsrOahp79SodkTtmd268g6+4zwdvJEw392pefIXc6alj7ZedavALXaFjHSFuetcIn7pr
5sk8NxMp9waIpWKBBvQCG0xRhy0KWgbl6/EQBFQqU8MPO3fh7DBzCbzgzUpbZnqzYtBQi0u/dX/j
cVFvrcG5EGqUk6aXXKwD8V67RXoJO8cGqG+raZptSpeYyXtUc9mzvZn4Z1Lf9fUqiL8oQcMSv5u/
fxDNEPiBOBFbe0O9ojqSVOtvFtEzEUvhSDsEqriveiGF/oE9o72BHZB0BHyKNFi6TjS1A7+3agMa
/GchWWdkStJf0jP5PTyQ5zLgBI13OcHt8ySh52I8pZL5hS/6YxWRjeZMZrwsViOe1SRR5z8Uner3
arEk9QFScQcnLMJEFxRwPQoOEWDxYrq4dE0GzpTnqaM5yk9LxaRnauhMNzslZpLyDzE+fpIVvu6m
HldifmxRjgf0uZgzrln7rChK8hbzH9Zq+4AhOViivH1fQAKDj19ziSb35vXGBdpTgvCAznT7H8Rq
FZOPvAmCL/cApv9j7eqokSRJJ4a+qdVn88Doo3f+EqvLgk3qGWlgKZETWvpYmL4ztcanO+KdV33k
M668rOIthxUZ6dj3IVqAuGUxs5oixPUzzcue6Tcy61biapy55iYolhTgPGDWiQq8+tEIVBm7BK4G
wq7E0gznlQWDeBZgm6ISxqIYRN5Fo1vN+juzfoB7OmI+USStHZhsyhS0X1ePhNrPD/CADlQQ0Ma6
rKHDi7E/LfZSeiUfWd6AZ/nhl+604eJkYde8r7f/NYGwc3dCqwDnIYHOBLYqokc5jKP8kzUYqUSb
xeXkHWUzcmg1g0krDfFSIXMYYS7AynHaDX+hvFGyZ9MMLyCZXBbGh7TWP3AoQrE04b5rz7vyjRTN
pSuSunSD0B6DA5hZPw+t959Qg4SvOnaw71W5hMjrMymRBWV6VBUYfY2mKxjg29K+ZekvqhLxrKLc
j3ANVfReMi6tciRzIBV36C4O9P65OrAYnuZEZeByJAe3pKyHe+a1lQoq6uPLN7kvUTRRkxP/0lZB
E3OprUnmn1SDqla7rPdpqibV4zEcrR/LYbIu0UXI4VGN4R4mnBsUljgxk0olbYHRLVdejRrCXcYi
SDefcpDJ5ux+6/CAoXXWV75cKomXvRyHfTmhCpjIBq5sRoKiagA6jnv+nlx/qJbIBqPI5+OYre8M
7BIEUbPo1ZGgOEjuewVjhl13+kvJYXabABTkCkm3VBR8AyrYlDj8ce0C/EEPKmteMWtdLDsldSQq
SL1Ft5mLj3xVlT/DrNXWV52Zjbv4O1S/gh7P7iIe3NdhAYwmzPjsv4VEtVCqfmXPb8xWPbSjaCuI
ozqOK4Jfaosz6uhJG5wcbrucCPbDRPSbmCv/XYDa/NksJ4KJIs5ButqU/bX9ZU1D5gou/cggLiTf
pL68HGSTIEmM2+RCAcQ40yhaVwMulkHG+zUFLLJ3yDIvk2eqfYWfbwYibfqQpZ9pt+3ibq0w1FLO
pSkzDLur7xtN0+I4LlN/M9ACaXei2Ig3lRrxh9YghTZ56bZYNC2871ZvfPtcg4UgcWLtMkhhlh4s
KbcDEhBqGroW2OBi3ZY9ur4Xm1yFbFfL3YyV+0nzb+mIJAboBQ3nY7PHvIfBFqX779/LH3JECFx+
lcMM+acWaWmWTTtDxuElpDBehN8NI1Ba63vGrlr75m1wp+OxYLEqV3aUNbBZKxXsR17XUen4g2hk
7DyjzyIo1vLMD1D0RRkFANG3ECzzidoMcXFB2X5cEHGdGZEhR7586z5qbwzwBSik1No8vBrWU9fi
lstSpkPcmkZw322/tiMAyRwolVCl8gjDELj1utV/uwVYb8pgBgIXUyrGIaiO6gKhG0dAAnjD5aWt
9WBfcK30AMqECjpQqKUf5RvDAHGMTcGmLMvPUo1RdFpGcZdef20x5FHxvbnzWFjARS4TFmPNwh3A
NAX19JIzRyZp/vIcUaqZ2Et36oYtdytyHMxqsZ3KHPphEs5v7GyCKCU7Z1+RbPlUYIG8bYCn/ALy
9nIiJkhOymeN9TPzp2BgE+sBC4TB951D6VNdWq0SjzbmqoplZrTL+0yeXeN2KPeX9IVTMU/aHGjD
MFjPVtlTo9A+js9wVSuxLa8pDgt5hNM9h3ttPPbVAnVplMOnFT6QVtZGopuCu60qMM1o1QuzXBqh
9svswzzCSxoFfj9WjjrqJmx+td+5JBG3nDqwZZGJxzTaW7k0wwhb/+FNk7vAYIMD279fRgmWz8YE
63ldKWYLejgJ0yav+tAgWBrBpnw6JEe7ToyFG6tZR+QZ7GRE6mz9kuJfMnFh95eOO9h1OFETyBk1
sfhzci5fDfvOOA9C3irloJP4skhLe9qgFn6+SBQSeeVCeDacxq/qWZydl/5M5rpKbroIyNWdjOXq
zOnQGoYEKfi2FsM06QI62FFV25y/aOZcLQfy5hf3OA/+OfoxxErmFZhbIPdZgROpV1yFQO36XQoq
afMhOELoQl9Qjnhac0HWEAsPUPLtuDeesxD4KmDt2hrAskyFn/nTtFWz76H0s3CR57TGA1qdcllK
iEoqwF2Sx5W1GjfpiHRvqmG7Ik+T3+2LLbqlamJf5Li0ZqKoDAAbKOQZdZR2F/ddIhPc5gwyjxVC
6Gt2HSxOOaK5dWgQYQ/6ckHJfA+K7Hu1fY9imQiSTcHnufsIJcfVQF7UMPR+ME+pM8iHIO08w6OU
LHOLFAMCQuLRC4ZkE5x4x5aiTfM+lvdxK+In83gbQf05y1pcaIlsvfIw06xFOpGdZd9j9K4rccGq
sg2nWlIarKKmlP3ogsa8VxH3n0gxY8Y/bka4W9T8Wf/0xJi2Nf/9AFDugmrfW55c0YW/mpZVzgxD
8krL9h9ugJXpsIXp18+pvXQL3UqmoV6jMNzxfpeCXGcJoPLgyg4mEq8cJGkQ686zRYg/MUKJfFW5
wYh2A7fdV5MFa9n8QWKZd7B3RN5C9upvJdHv8KWE/zlvjEnCc0gB4IkEpBkzVbhY8Eoa8rmQsbRF
q7ay9hBKDoLVo+1GMN88HqI3MdzxI6gWZrn0323yFblpnj0oHIg3zaEy/K5sJ7HVjst0EXZDeG1E
WdGwqbtaUrMy1trLJjpAE7iW3+ygOFtF1ZsFMtR9MlpNFwBTLeWTJg9Y2RMmVSHJVVt2w6Y3nYl+
jhaumlzo7IZ00e1rfr5dgrpzJ/46+pLq4kiOr04tnesDqDghEFvz/SMbnpV0yHo1um2oXHCfPf7E
fWBYkqmp+aVx3Unm3+6fnuH/E7uYOLRmMhlkvpXyBfJd1tsyfz4ghAbS0x1FAw0e/Y+OuSN4VKFH
4iYC4KzfHQk2KEzgQ6qcxIqUS63jGsMbJIAxAnGmUhG0lmCFJ1ttowi5MG0HlKSTXhF8LHqIPo1z
iZIZEbNiROXuPRSE2NC4Tuw6/IcD7mISFedUefjXiZ/FzIXIO8dGmTCIozMxB8n/nhLCQFaBSlKM
4RLIw3kpLHTLpwcLEcCYCQQIkWg/typ6IViKDzZk9fFcP7eFJYSMBTlIuhkSFSXscC8Sd3bDad7n
uGuC535aWmPeDkxJQEFJJKDqbnsNvuZONqcSCIESnviu4LMJS/e180HsN0+MBvzbKwewg+fxMWcr
bSu0w9uqEUgZfRdjlf72Hkk+QaZvvyThcVQDCnv3e2W0sEIlWLfPH/bQFqPJkI/iSt1y10ZXF7RA
0gWZksYxxousNjivTSLFGd1+lTe6EN0KEP3wgGWVrxyPYXkyNZ/AEg6DueGHx4/CnXZ1vtY91Csf
b4di8kPz3SI4BwxFn3NokFx9gUWSlgndtVJXzS02eDPWkgj5qj5TE+9tSFVWwX9YlLAMjBj/W0Y9
ZTBO+RDVqkMJjEyo1xpkGXaIqB/RKvABoyyrAJfVd03wliu5VudpPf4+FjztqtIBx8mF6I9J5t1R
TxOgs5nvJbGf7KqJz5tgTOwt/rytXGDOqVit9PJacyO3jNEs+nACS57eAv1cpKUg1XL4VnnAmNIO
9/C/bkILiDkojry04aHOuCrk1pGfC7xzNcCNkcIpqcTxV9wudfrkB4jH9Y5PWevpgUkx+Yeh+epI
MGmTNoQ6sBmyzPlSQeh2dlei8DnL6ftpmNvHQhfhJGn5HeMroST1M5sAxBp7HPtEkIoQ6v1MDATu
mK4xpeRjWwUzlSPsc32IngRsYiNFuIcHxTcHhp6gvtHjBnNf7rFKj+KnORauQwuti+y2E/OZWgkX
nROWid64b6pRjDysa4Mquw87wRSp5qdtNhExYe5YmhUmqjZFFTqhC2MtLTe32WKWq9TtbzCbmyO5
+Fhfi50Pc2Q6IGH9/tLrGmUqj+Gn2mI8VUOQT4We3hJYx2smNqnxVrJmoF3q336RNumKE8frwMXN
kMeaA7uE9WWDWujdRzhUWV70i+Wrqg1RgTt2OfwVIMlBrbozFcLOuKcow5ZCJU2uqH4ynnMicY2B
HFZhPnmMBlLLS6gT9UAKNWrS8/dx1Sk5VKcD60dCru323VL0ZD2MxW8NpMMIkwV4aqredlTebgkI
kz+y6srjoM1USsAD9E9YoL3WhYZy/Jisn0Uhmv7vCrP8cln8uH6EPKoKVsTkIzNDboWcUyz4ioTF
cf3T2Xg2rk4uz3hqZimw4mtYu+B5y4D0LTy+fZdk3BWfvHMqmiq399+v0HWqocQve8Iw1k4XQJU8
A3Dfx2Fqh2WJcSlEIl7esBMgA9vKscIKapAEdrMtjEbiK2ZVW5VQveMjpznQh8aCWK/f2fQOTyvj
PYzxqwxdBpdXQttTGa1uFS73UMoZbSfX5HPWOnukzIqGK8+3yaa0pMaYSmKv/9okpOFZOrVoQvo4
zQgZE8yOpANGWQ8raNoNelVYfKzHAq2m6if9ye1KghAivXbZFMyCb5NZwqUNzLpSGm25/T+E09rX
NJL+YJ+BxZdxFi4ZJF7O0oW7zjXdfGhpCbLa7+1NubdA724gvhHnsN/Rs1gxXfZqPQtx2k+zeRAF
5bE7M48ghQr0fKK0Z/I9WiOwz/tbP/yY5GgntTwo47iuulLm2LWIQt3bBH0MubBvAa0drHtGzV4l
+dJNmvpHOFMNAf4WuUaqeumq1LV9PZIjs2zGM5h2CWQMp8bUvAUseENJRmWDqS7qmmErWlQQCXPX
DHryk0I1+euVSbf1xD1eNqG9uXIG4wxJ8j7FBBW5iT8Z6dOGKE71LjCF2PufepYCo7XmedAPsAsO
g4FTpGXkBECeb1cXPU8a6UAiDHDdrGebuPOp19Av3ZnFogMur72ajtEHBzmm+PIusU3w3ULHK/zR
XQffUoNftRwcGhEpNzbq4WZe8kzHV0vHMiBRX/d8+dfJynvjSr+X2lGcmJkL5MVLm3PkpxjXHnEb
hL53KCASjtoqcFlaMpNdZP64FTLR64OixTufOipXKa6hGWjchTCHaycQNC47bfXWgdEpjPso81MF
jNYcpG6Belly8oeHZ65RgDw6mV+N6fdlBimPKE9/Pu18Mi87uW8vdvEpyJVpuOP8jsUo9A2CM123
N+izvMghX4ANmU5U1+heb3RDksw8hN/Y4DegnccJsR42+og/VNLt7SVwc1i63vkNhPopBNYo5jQU
fw3LhqbGxVW3cadLpb+Y7gqWMZj6Wfe0iQ4Sh5kDLPN7lvavhpGAtEkLnDKjieY3t49dzO0Ufpuj
CpvHiFia+lyqK1Z0w31Q0muTrbOf5QrdhjiY2fmtG80BMYLXsauIIFumpUQ/5QJlk2yf6RuNxq/e
72KUJIyMKREcRnK0gjxm1GKYbKSNnuy+HpfIwKDmv0qXx7kCrILD7KH9opCO0KFtTO570MNY/3uF
wPwagMWveSl12dxLyUoqJpLN4GIuWF5SHBB1GcuJ5zuBZHMadDIF49IOyHP0QqV6OIPPYDcqa4b1
T5CWEGeNIuvmH+sUnL/3UIlSXcVxjHE19dorCqqccUOWxI9pfZ+4M+ZROFw71tIXPX8kMESMl3OK
3TGRG7UO04ntg/lcxg8hB6l35MWe3gd4YQaGB9YIUw/dE9HR1oMFj55GeFRF2KAFreq5di88XbfE
3iV2assmQ7yaQ1weSX6C5EC79PCZun1B5jKpEkd67o6vm/RMgOJ1XOo01r0uYx7hnbdxUCG7JcVD
YQXw6gCP6PIGHlunyiDi3CFzpPGDaRUpW2EbwYPTs9XZhUrduxTPTWJbv9sKYraM2rUSBL3EXZeK
g6MfqUSXFTtkfKwwGjDMmEFu8hvteCAZCe4LaFMqbemdR0+7ifePEiIgXl+g/Qw7YbjJk1tMh4Qu
a+p2mE8u57xY60taGYQP7l5WZn4nwZrnPBBkQuWFgUgw0LqPNpG30qTkLFzU1m3tKR0zvLA9hDY5
XuZvufUUdPAjFI/KhY0F1IC21Ouo2TtOkh+7MCqbvqQtiEQACzeo9dmYWuhLS8sJfUAa+WtmtsXs
SOcEJJCmJQYnpfDBMx8a8/Bv265PhqNl0bnEAPOArjXHTuhG5INtd0RvZfHW3LOmnxeuvvKiH8kd
POeAUTQHSLy7QYqFBGRrBac5k2w2TcO1k+tudYSMH+gTmEiDGiiU6oP0BhgeWd8lzW9oM+D4PrFA
D1MIWZNLrR0gEINDgpLSwKwmw5ReaYQodrFkUhLc01YRBuTFgp8H3sWb9PusoYHkuNkou5Im75PU
DGimKWiM2IWZXLsR7yZntcKu5vR4oCb4z7mA0YuqUPK1dJ2E38/J7K6MP4SWptpkp45etsl9KuFu
UdFPAtGfHxwfYKAgGPpXL9KcSupOECTCm0F6x8urH1bCpKgOWEbC49RknExRNjKHGhh2FYI++/DZ
EuwX57nGXWZ5ztYamyS7VsKOLU2r/iOaxHavGaftN9zZ3FDnuAiVZP70NP50qM2LrSkZQY1LlGzo
5hT5qiL9gwzHDhCBdwF6Ab0w1XrmmXmdJx3oHd2ZKncz6yEAaGezi12vWG+hcTHio6ccXGsgadzh
tOy4tRIjhPLlZ0BysiKn00Hq5cBjCI6QXQgAZdY0EeUDxforKTRQ1M2b/ifpRjwhIXL6p6KzP6oB
1KDImSNsRJMzxX76G0u3eOZi+zdSRyrPI3ODbFysJygtgigJuBFDkwghJRv3VJwM6u386nn1Ko8P
9uaUb3zZ4K4QrNWmHNukkgmWtrM7JMTs5q4m9YDXtLfsLm8G59QaHaLbZsvE3GEIwFGgGYD5mymz
s5Jaje+bfYaDZFDp5mrGo++VGxblPQu2iOP2qZINh9torBkchvwENktEQvpkh7DoB8Dm0N8qArXt
84dehUT5wOMq0GSsQQoPIAt/SNJdbp77wp+RwgSpa/gOVPOHdocArCgZSjJ3UkE+HxV21zUKF2yc
xg0GCov7C6jJsxnTtPLHS5JE4qF+EzML3370B2OV75NclVEXjJDrN5KgkLPhKotcMqkcNhTJgc0r
jHODeqMJtqBqBOsiCBRtjYgiNi3uSRMaewN7UaIK0IYEoIXng2dTSH9vnbmqENyUEh2VeZ4+tEHq
isUUv8ychNn757fe1oDJpVpARA7f9dv6SBHykhGNFQ4oRZh0OQWtovx++dCV4BSQ+5mHLUME3mWE
WUWbM33abuDNDcEkqmzyVMUTB/DAjk0tSX3t9qQpjO8YEMy1/UKpLpIas+EJzWes27MmUa/+KWS7
EMdJQYn7AJo6czaaYSELM83fz3Rwkq6fgQJKBsx4ufIUmGm/Sa7ZCpNtrZOO8mahd3B0PK57Ydyn
D2jASJLdLU2N1JnGPsbmi1mP0uXrO2DmpS/EQBnPKlPuqmdUJAudFxTHfnkKx1UjN621MjpyFbXY
o+MZ3UnX4sGsVBLRK2KTuJ7vUhu/sGmuaQTNlg7cGYqZzuLq01450Qda/bGkK7yUwOuHHj0mrYKH
gqXVUYYrhypIytO0PW+O/VnIr/PLB+nPYPEHuLYzlgpx8+pxfilPf13oExq1zUP+XFMLVM3WSDFI
+v5lnZpjvIAkkioD2n5gTajYcUt7fEhMj7ej3zCY52osMM+vZVG8jKoqTmpZmPOiquraL4FhlyC+
mHKZ95+NWI5DThqalJraAXiGf/rmi4eW8KM1kyGzrDnITod5bscI5fPxBYDX0/jP3kcCJiSR5SKw
OQs3MFmMLl5M6wlkN3TjNyHXHu9Th/n2VnAbnZ+WUYUje4o96zewIOKdekicAERgLOND21Jd5TXf
b/OoPd1Lot6kR+HVZd0SGOuMdf6RntZccNsAAJEKmwwssB4H1JTCzwwPIJhn3usrO1se3RYM4Erd
kalauvaB+AqG83/Bfe3iz2Mfz5DT0e0GTtHt+dcnsciMqZxmAbMVGzFqWMTkdKNp4rp+d2bEs4V2
YGpKZggBEN6PlLj56HQEuW297zJo8hnHjqVmk1xZ7DItdeBSLvZJhyCwMIY8JBkwXEtajVg0vXvu
u2T+uzhF1Fdn3AofoK18nYLNMNzM2MJ+hZcLCdm/ahOZx/QV8fOvoDPlUmXy/+MzkyB24GSR4Bqi
Bbbh4aLuweVwwClZGyTBI3Rm2frcpm2MOO3GtgzzO+Mv3L9LPfhi39inQFKxfeGBqgWXrEjWVpo9
tiVW+nd7Dng5B0b0biTucZqiRdnC5R9/HmkQXbXcQC5w2AeK3UdPixVBBFvPuNs/3QidnN7WqBH1
U5eKu2ARHAIsi//v7HWfjbEyIwioGfmLvTc2sBKGhEMfXWtwqX1yadApOhDyIvY/TYvQOSpND6J3
mw7bA+X8GfuH6pFXOtfWHCMFp+WLbX212DdihWRuqI7yRMTx8jZ7s/uhNVDCcd+52DrN8/AHr69q
+4NgFju04qv447rI1uaOjiL/qs0n08/PXhxkD+oAHCR9Eez1U7cWTg7semvxiYW+trsXF7zbdiUu
TticzyMV/MdX3Sy7F6Xp64TuRS4GxrSv5Uqs34rmvfiuy6DtoUyj8eJ44WJwkXolX5p3kBH3y66m
a3+vu7eBi2keFzmzL541QxokL0SLQ7bEw9hGchtN+w2UtQm4DsP+b3Y7L1D1S5lU8XHrb9ruewO0
EqpkjAgh29XD2kjywmGzfS1zyP+Gwp9tS2EwgZac1rM5hVw5sVlDN60FNZSt1v9OqoP7pXJYmZnO
eG+ZkrYYfG2jLTu2Gwa4LJ5I4Z8UMm7+Rz2IMET7ErS5O6vI3X8ha0BQEdFma9xYEXXc14gINOPH
cUPJSP7TOjyUcoccDayDerNIsV9U/6twUE1gzE2ctpTCnADoQF/IvotZlFH360+EKtoGydNmIbyS
OErkq//HCscoDymsIL3kSxgEVlsfk0dONLIl8iw9wK5+eH7EYVtEM9OUh10Udf6Y7+H0rJk0Gwb2
M47uI7DT3SGI9jm0Kkhnd/Mviw8GZlFNty09BqR3curAjdibKkTFQQgI+i0gox6qavODI8r9zj5z
bgLRqivek8UWSRituukz5jU2wJJkJcoMqYASxfrxCSEwsaNvgar0HMUSxbYM93vVi5t2FhlL9GnH
eOylpgPxchsjNs2tXnRpQCPP5VmW0ubHQe4RFYWZD/6wVZ8MzrLwqWCYMQYSAXzPT8UB+IdnGx6n
AwOrz/g2V4MeCnigtRl01bgGGQSPIN4JEbYAv6WL4jOQ7n2KM2bWqwIbAUAFsVvrast+CAzgVk4Q
a1/2YpnhtCHjJyVwYSwQsGgJHD1hP8qjn4OXMcwrR+vZfRZPHoOY/ZHreSkhWD8Ohfpfl5+Phfxz
3ib6PYTbaZ8VIGHURC5/IYwdVho4Lc9i4hb27qY1NkIWtXAS9l3opNS+kRFK65MNE3vUS/XKT11L
Nn7Np7yTWcdI2TDeEIikXb7V/BGQauiuxJ2g0OHpX/RF01EaSzp+y1/jnD+tK5TUlM3Mr3HktjmU
fA91/nEzPBl29OosLiB0di8HbrA4ksOoBfaLINuRgJR6TZvu7O2toPfrvDVQ/Mn1VyiDpXPnbhMV
E/yLG0+xfjC52EG/aNgFT9ylmYjXj7/j/Jm34FIAxzPzqoCWxhUnfilFyizX96KxdcRTCmWYGgfk
7h2V1CZfOLCQzth7LmYjzC80UlOltyHeifCfw/Bn4w8CkqPqpUz5ihLDmv4vN6McilT73NANWi59
V/V8Zp2UIWQjiku0WGEmWuRyR9FdSn8LSrIGUGx4C4PyGKEi4xw605RspM6ZpQcvuSsgXQnBTIrR
cxL0Utqys5XLCtCNfHeh4EYOXfLik+42S5h6iPuIGDXSdOi1oGqosj50oDtIe9XPpamoLZ4sEMl2
U5SwEP4lpwerANIP1LULoFiVqytYz746DzZUBTtm1fMP8x8KdnwQX4KgXLDMc6/lFK032F5cDDzQ
ncFCTE5OEL370WlC5L2dZK0Yh4T3+fZO94jH9T1L+dZ7N0WaAL+k/H0jcqESNG2QvNNdFrcV9IjJ
Is5zLHAauVMhgpL6zyj4OpWXXvdHLBjxPiH7Fmy/j/+LZ3IIriBN0+2g+249zf7QGpnER3USZTup
bdmAZ4aUVeTrl+mqpT29SCnHjEsTeJ9LrseN5l98Y+VtVRj/HGtsg2qpo3uHcDHrkWH2QV0HSXrV
GbJk5tgSG6j15cLE7CiMVEI1J1/ukKwaeKVca+WQHZx3EhaiOJcoq/QBIVb68hbz+b5xYCAzzMu1
+jiVogCPV0sL17kB+o5gpBG1bIZ8Up+SillorJZvMku2RwCrQgyzcJ/41yVN7VqYi0QkeFd2oAMR
i7pIAwjIBAjFEnfZmqucmFzYYfSb+aw5LPHW26sLmvsoBiwnbkKqOsBkVbtPTGdTOT5yo83kPhg4
w6jgSg188WS3d/ThulHmRxH/jceIJt71HF1Hu4BIUCWlYXY5NDiz7VaW1qdB9aQNJwQNUr8ISeUE
dsXx795bgM1diC1ra06nb4fl54P/Vvzw1APlwdFnsE3ojDraX9ef5XM3Lpbet2YPgHfm+EjSbP/9
0MKPll30NO91Hga4lkgdR1UmH9Todhuac0MLX++pcqTMUbqamrxW3fP2e/3JmK/cw6v+8DMw4nGw
Yi/9JQ9WSPhCCuKixhN9Jl11SVVGtHQ3beMOSO4LbVH7uFH5UuzJ7OUNt3BoeY/8MeoZvHhXyeR/
OTqgd+bOuvw7jpCPGYihKfweWs0o6VYEzB+ifHORm9OxT+K2WHqpOlFek5GPWuxTh8fjR2vi72D/
VDpAV8Oxx6KASVqj8jVdOy6wl1mVZ6si8UDGJu+I38QFTBbqEuFSXBZSg5FlwgYmxbcLaEcdHSKe
Lazu2OnoYMGrnEO65wxHsrV5BUnsXtZvGEGEzdESZhfEFbX7eNJaryGU2ntWQS6qOAF2BgID0GM9
YMdhWyBc3pCYTeLcnsJnDGVumrGjdFxnjmNJxUXwo9FYAaQvvvhJ9IF38TxiJzqnIsOKYjbpek+s
NYhZvJmRJOCWw18YAG4iZuaxYuIzwfltIERlCwBQtCYDaFcMRT8oc3mBBB4JDQeQIjyvSr11ri2v
XbegYdDfxFrwiOBgcNttD2QAOJVmRrdSFKqGX4cIOH2mjsycRMh6EY8Vbu8EXo367dVfQ2iMhGW0
brlp04sa6uSOXifyPqLTORr/MXMqh9BfuqcexMBju29zEB/zxSnjnOA1396JzPgLVN/i2AJ20WLv
tPqfIftcj0lMQnxQfx5+geDNdjF18R6hoinvBZi7XLf890b1E4RhFRcvHTHDpZ/j7d2p0oasgFp2
SZPYdnqlXsr/g5DVbLjVPk4as0Ad1etmMH7k+j/BBTHXoVVfL2wOZ6z32Rm9IJ7FO6b8qZHZWk8y
ooIhLukgmoi11q4Z/OGJ2KqhZaa4qvVBL6a92Y9nhGdSqA2fbNgkKIPLiNc+Q0lS3eEguFy20HsS
MT8iD3n0tknXpZM2W4cHKlAWyPHXbvJBSVfbbx8+8rzuQ5GQZF7RX4nvfaMFg/hkCaINsPvv6QDY
Qs02N95CLE4+BE51an5YG/NROcO1dzUZNx6NKQ7yTA3a5MY4Y89DpLBYyrBPKL/dJqiVH/8qdss5
EvuG8RfvVb3HF3rCV2W8in3yl7qCqC+Dsrn5T0QEcpeGckV6gUj2ji9Hd5w0kMHp10s4LZBAb/1t
MRsTPQvZ1pHAKf9QkMARTCCnG9jr1suelzJDP0RtPkVQcyY4ODejrUaJReAVwFvyfAbOF5a3yRCo
uRqrNFPdK7HVcuqWxSKoQ0ocXwKU3SWMrdHoy3vFNaZZ1nQ5tJOCOq8JhbqhLGUhlCRYv/r8sGcH
RXJqI1VPg2y5EtlseNO58JcTYIZqcFx1NcZLspTIlD9WmKQSIB98JyCrKKjAuf/INbZN2Qp5zCGW
xcnT34TGOhcUWjfrplQEYEhFpCctjFlFWkiLlFyU1+3P+SowU4gUvKdw2cKQsHnDRt2EjM6v2JK8
q7c3SQFFijcSaeaQ/Tv4ltANJWrti6pT6oULWZpRBl9qVyWDz7jNEeB4i6Xo9D0TbdNWCn7ZGDQa
WcIyALijSM5AWoa2eoveaB+HReDM3T6u4q0PagOMbF4J4y4pE3kaQQkO5777BF72qFx5jtC6Q79e
rZeqjJ8Jyna/HvOk9azt0okq2ldnfKlqcRDuvgbGQf2GolHyvCBnowNlsaV+/dOPSPpw4/TVfB4O
K1yqMjtp8C3uUjUS3L+ZLkWxmpDDCp0ymOK+OAD6e8g1FFQnYQ9oNiqzothRSc1L7Ut/mvqS/NXQ
se5xQu/ySZxdd6T0MsBgJR2bUB3B5RhnA8HutqazE1xsf/f06t/G0WwdPgKi/IwUFnHvn5qgGU3b
+qBZhgt5oD+CBA4kLlCDxWEgYmjQDvKH/VnbwnH53BujmGJaF03TCgjbeJheTvQQ8qmILUs4df7T
IM8OPqhldfizxFrkijUDXGkksGKc7SlhWaoSIDmpY3KRd1fU41WAnQiPhhBNJIIzvRH4B9kepKKI
Tnwm4Q3xRDO4MaDxp52Sw0nM5wrkUr7MGDGhMyvND3PLBjiD+VATN0eT6kkpJXWzb2YlgoRpoZqC
qkcnu6bDPK2ZCBPfAHzIA+nd1PQCCoIeKuZks+xEfVDapfaSeFmz9AVm3kK/QV4/m1d8PMuikd7M
brh9KdmfsCJsw3fod9ZNpKf+G7/1TgdNw5NMdMFnnilU89K6W2nAGFZ+o2xkZMg2Wj2/IoYtrpvi
ZobNjxjzHcQSNVYcCqzYpB15vr2U/dVUu/4eez+UBlv+yytY2ocra+QpAk4r4YpteiE0VcXImnrW
J8lKW9PCY+TgRUJXNtR/ZNmi4xg3fQGVM+oKK7B6hHuGce7aylxHX5YhopBwgR0tTxy2dl0766HI
WV93WnEX13dJze6gg1mSMYl5fzpGi8CEmZo+P43xI5kStDT1c8yDqdDls9TjBUIjOzrFWLX8W+eq
p7I8EiR5fc73aqtORS20edg+iYWcoRfhxDH/d5RnhH9kMoiatYpiqjInZdZs/2jLtmm5nA3+UHdr
9sOPD+6BDEYJBAmdjwUHDFWZhJ3rzWLGDbeDiDWOQiRH8JjqzBUKf3SWhRzNnCJpawtgxmXTDe4P
s9/GmQBPD4SZsSkrPyoGwlsUwf4T5M6cBNpjaJ1KpjsNpk8XI+Ihv5bB1Js/Jvv3o1Giq4nMl53c
N0qEy0pYP8Dfd3fDTqI3slHCOqMWO/h+HQrT86a/ifvQMHPEVWwJK5guwaODD3WL4nSerWe/apLE
T16GDXnge6sWYftLgxOtTPfJi3BaLCqdmTJxulK2cx6rsnHJYcdL1bow93Ao4oPYYvGGXCH/2p5m
ZH0vlysjkxqiXOaaTzqBrq+TadvxU8bNDlhftvr2SC1KM0i32ELrGrvgXc6thUXfRGG5aqgZdAFi
z4P6f4KU4BqFzaTHS6hLHgumKXCylAG5VFE1Oh1PdG8BVEHI2xYNCCwyl3UZzsvNERq+5tLOgGoe
FqfJkndE8aJwojHYLHD4YEob1/Sg9NM6PgPAnWHjV4ClFScIJ25ziQIjS3A/DtiqkzG68kAXLsGF
gnqsNnEm9wrD2vDJ69qAkKCsNTvQen8ruS9IXusVKJp1fDaBp7ZqFf/ByMLhHMYW7COFz8+I2INY
2cDMLYPJluvjbxMis5WWVqCD/oiMUjdry6dJBSKwTh21cd6nu3ULKtW7s5tVWhE6TUnh9zbbk5sz
fUschLPPJd/X8FQYaO39sWadtDUFV73NtfkGgAVQTbbUTIfAcph4emqHFKe7H5AM8W73SohGDzts
1JLmJFYJF7wsqvAbsrfjEhMKg/v9UvdpmLBBSjgHq8Fq/kb0OzSxzyW9YWR0z5htJvucbSYVgEQc
dLUh94f2Tm/BuJa4VIOkQbDRX6gw6tsbwFR1kgtxnrQek95xilSLiFfZoOKwwIvcy2rc7b7k/b4z
i323+beqZHQW8ZT2LUlHhSDZ3EzFb/PtWxjodFT2Gfp43RzSOYYonNCUZHQPrWjtsgOFxiY7XiDb
w2MRAZYYNJnNP55CnqFVTKMsr2TJn9NoF3vJ0OYXrSfnpJum7GEiDsy6IVKWn8phA9L5I4QrRslT
C8eyogb5iWyLtQLP2pTR+QnXSyafvyGqqKZfD9O5vXwpXQNxD73kQY1EidffKhb6GnBe84A4jEfE
SoERZaMATxykul0dAHsZkfJSOIeZ5kLHAp0cc+XpLB963jqe0Gm8kcdgvTFPy27rhXy89DoRLlq1
sgtiPop8Nu0BTeA77JKJscJDOBcjhwttOTIgCUJCSMllMCT/J1hAnlJT34Z03r8b+9BKFg5mx5Na
jUrxDi1o7LXZiZPkCwvxTWW9eahurY/APiuA2/4UnAcALxZGSG74qsStxX4xuCGLcNfYOrPsxvqu
GMi3yRQmJT13qdhRlgK5w1KiwveBuO1UDQCXXuYCiqIHib1JUlMOIj4r9Kq1s0dV6mCku7L1fXrq
EYn+ILonCTTl+64xOMGfPhmCzLH1Y+hPBYsyHX8AwSwb9IBxlXUpxHkLAaXkuIW2D3WbNTOlzkYH
2Rm9Fmre1+D6tPUNNVF25virsQpXQLCfNNGuZnTySHt3QsLZiYwEXgjrYTz6cnqAkCgSwet/mY9E
mUwdCyFzU0+WZJqIlMXLuitg8f0WSQbx/d4x9oKe4JRbQxX7Dw1lsJWKZkbt/hhwDe+SS0/Iz5YA
l5yYWWjeSWXj0agdz06j6BapnF9EnqMWmfm/oM7H/mDznFA6gG9uYIEQIfus/Hifi7UScSKAihYy
x06sQCNFSxaZoLb52E7e3eHo7xu8DxZuQ4oZKUkbHKK/woSKmcVKAQD7MKTKP2iD+NznAfByT9WS
gKnAlUBLakMbzx8ZEL0vuFdWzS2fMg6sNTul+RH9eRM/vcSXYt8WxrUwo2Vpm3kHpTSrqBLs/pXR
nq4daBBmv5GFh27J8chMffRPNXTeCDxH23KJDoNOHdUrYlhBWyC6//3vLb1uqBcR2xpwCHGS7qPM
/KFd8A0Ma/iwut9d5jXN+Aaei0968n2285MNO1ztkEukwolnwRuhScgkCPEcO1tkUnt1bQjBA/Ue
phwVawoPkK7n0KN6B5pz/lOBnsksLojMMBTFqFkJEdHg7g/tO/3R909rojAPtIxGwVH8V3yY7c8X
SMfB0a+HprJtp+NG2Q84mpX/W8LObZ6nk2ZPrIOKDSj1pWXljWV/O8z008fsdOjSqTFKvBcpxHgx
vGxb8O4e1cFpIROC66PXKfovNCVfB+BMBwEYLzM7KFrK2oSv9PQZq7c7JfxBauH0Bon/l1u/dnUt
pRK3YHBoYzcAOMRO+NHG1fPBMAUfeUekiwvg5IZ7nsCynSLKF3eqy+HzRX2uSGAiHroO/eqB3D1z
CqqeJ5Tz3hKNtuZwaKjC2bcMEqHJQ+nDB4Ql1Onxf7+AgRh6P0YaDQbJbQic/QSFiRm3L+Qprm8q
APJUkH0kPLDzAy3DUkGC+pra7+6r9UuTYuwy2SsnGTZihkre0wECjOLp3SyIAT/B/5pnlPCEekSq
hlf2reWY1deeivWS4BD5pm1FkjN7GVWotlwAzVeTaNS1MDh4ck8CAhAUAtsEwAekiPShoJCl95Cm
GqppPSgd4/vkzgDxXQFwdlWU4arCibxLyxtQpzv9/kBW/M1FS8xNXcyI6rc6kZaZt4Don7JB9aOJ
HAOagsYQCJGxHALymrda/EQls952Ku7jahQe/Ftv6gCj5aI06nwmJe89t0xlQjQNwA+pyvG+maZh
LNJ2usU62151fDszMFHKNi+zWySCExujyhRzkVdgXTOG1opkx0ln9i9oqJANZP5XCzgIxwSgxLUm
blDDSbSWgLR1J5NSXPMGWMxm4gzP1PTTawvnrMuN5te0zCGOZE0YwPuF2zCdbSN+GC5kf2zNFZjE
2JkHDtbeQsA+6b+qqGpXOpW+QXvrnGUv5wT1uouJmNZgJfGiX1d2oiTJMzThvGJdOInnk1+WLlZP
2erDbSjQlOnA5mxhM4whNZ4W2OqPAi2UtQb6Pjk0ueBVx2Hcs4iKLVmBuu0c+Z10iNDnIi3nCOdE
ZGFtNR7WYQYE8gLroaSUcxNMpqigAifXLXiQeeux+dv4XUFsgxrfSeMDWdMULlNXEf+/0j9dBEe+
bLwgsU6D2VE/S0BUY4H6/LyETJ08iAGrdRVEUV8V5cADSLaqloeqJs0duT7Ela1tNotWssYHnyE8
9HRTfAYeTjZYhmc7QNeSXBB2Om+gFGyRbAfY1yVXi/Fj9z8tTDPLBN//cvuFH3j1lGEooSqHOw6e
z2WMMWTa0UVCAstuSMlmV2USIIp4eNqJ4/Af+fHKugdNrTCofqdCdsPRSDWFPenPt6bRepLZdHar
I1MAWge3vjjCVpQ6Qfh6S096q6jx2H1LpGJ5phKQncONCxWVXE7rghakcLRKxQni7cKBMIlwwWO0
oWvABfcico0AZ0Q0LwDFLY5l9eoT1Giyc+qvq7TJs+xSWYQg/MuIaY79UGx6MpbdeE+Ez60Hixwm
OSKqwz8gIK/gSuVlJ6CLZy0JdqoLSzk/PIwjN4wZyztx9GOaUsg4LjUGG4SRLxO/2eGvZ2sjOQfX
CyRGUq2fOGHVWUGsaG0AFNzcga1CPqxVyowWNp8uUFxib2BAEosN6CR8gxgV/3kt8m7mHXy/O1Pz
LGOSHz6QZxNIGmlyfgPQbNgKe5LbzAZVRuGdiQ6UTNFv/jUbWGMZFhWGpDfwoAMlVHNfzZdFNeMI
x4GZtl9EZ1z7e3FRS75FkQAxgR0Xg/HWeP7ZpbX2epEpQDtvUKYLCQ+qpjBBHzPmeZ5V5jlTDV4y
VxjscAwILfZ92uN4OC6bqGBzvBUh0dVUrFdrr30qSJ5GsVn2T0Rqbfvbq8jkaFwtLVj4SvbrZq2H
/X4LC4SG+vosHACRosyBFQzDrU5rf0usaehxQ2TitafdWVF1pm0c07BzCULrQM0J0rwBf6d4zaUI
IoCJysULUxpBCXxLy4YoYX0alLTRF7LdV2GuTr+WUfMQaGxZlPssL50sKpvZaPsEYKFtCrz1cw5s
/Bf9dhpYyELAcgCFxiPM5XH0bmcycaMy+W75xs5TLb8Z1WNbf55iKtJneIJMouaSZKSu2i+yiOOz
xwoD+kQGQR7Jk1vyaNdyAc01AYsrH2AeBj5mtolxesHGfw/M/tOWEpl+1ZqiGpBS4Xz/lD3YDhl1
XUDNN5psDTCuMRAcGyoPDsSNHrxDC0PLaLVnOpnZPkdvOJ2+zlLtOm5vxSO0QsGoq0WxGmXnT3Td
BuRt/gk2kcHVEBI96cCkkzuWSpMEllVEGqBAMm0mQbgkWQh9sQxKNnXxOfovAOJ+TJJtb/V/K3m1
ZjuzNY4xMztql6QDSz3lte4sdAKgtFAal4iCECNE7HB9ZmI6YTK2I/UrqiJPBLUGCXbR5CewsVEP
h4W+G1fjOz0HhWSc3f5Yi/OJIlaGQzuz7/AsLNPDX7sOJESbGhqdTYAqNH08HfMQCmEExK0MZyaF
IG/13twH3rzv376Nw7cGFSFmre5Xt4Zb19W+hJAK+H1HlQ1TEgvojpvciWDVp2w2rkNeOhYh/caW
jIRwAzCsjrgGS+xQWGEYHSr0IhGDbkwg9BX8QxdWHXeQp7QnUVU8+C9p22blIarWtC0Xu+QFQ1Uc
JOCagnO6Ber5Jdu+WELzFuJPrBXGGTPMpfis1N16nSfGYxcZopNLsbQynVTfC1ZvCJF/I3PPFdnI
frRZKTsnKyK9vRV5zzEaM1tJYaxHNUnx6R00dYjT3u2kAEQUmd9u5KwaCN8kovQ+9jy6Hkrp3UaJ
adboET4riqe9bq6GDThydHzvd12BcLKfnH6CXG1+UFLZDXL8+edB0sf8takf/gOOHF1XxsXj9BrA
JrwklXtxVqnTe1szvvfm0Qnnau1M2FlqsXvEin+ExuefBxEIbuxVuhYjKilDKRZbLHO6Qos/K+9b
MG6ws+pk0o2NeXO01Y9qRsbUTIjluMYwTQHUVA4ioU8K/jTcHXcLrJsxCxgtMbPCp5l+cpIAmplh
sX1rZ2PNMHxcM2eOknjGYKHVmoAq/c1IqScSjZJdUh2XJA+iLN5lGccP0IArMTnkS2ekjbrfYvwU
e840dHiThS8HY/QXNbaOe9i+AHC0V4z6UrUu5vVZqy0cjAbcovMlorrsZ3R55TmTGiOJLCl1E/ML
AN1Ek3og9zK+HId6b0GV5FyOBoRj+vsbTC1j6uwscscFMs5QzF0txuhgRZUD1MaFZXFMCRw5+VrM
ooGlud5tEa3eNUaC3rocF5r3ydN/R/iWWeq0JSBeImaGNFyoTNVBKYceFqAk4grs4cBo2fLCjIzB
pdS3z3MY10Sk2lq1qFHHAE9EeVariuka34wGv6RnTl6TJPjRQeydHMf3M54BzgnhV652TTBe13gB
WmD+nxvSuMXzKj/6b8Wyu2dswq1KZkZA65bi+IsxPaRHVlj/CHMPRsgRFPpj5l7Ts8mWvchDo6Mx
9StdraWKE08rNT27Rxi6ixAnMIIhmwtwDi1/2TA25yh133YY6GZ8SWUDQnaGPVm3tLjdIatkrZhe
rY9PceSieBCYCcDLi3UyE0Thl8MHwF4GfUDDRYcw8X1XGHT9X9rwb65MdGp+2YdfBSgFxYPoqyKK
6WZ/gtPxvWeN3x1GEj7WnJ1Rz5r2W8lfEhbPhsvvTIefNKPqnCNsnHWQMlRMhBa+TA96biO9XFA+
37eq51PS59nhvrHD3WwYClY3DUpK/eccFmzHcZT7M3V93uFCFupvNHPtoE58FnsSS2dcHtV2DFWh
Tq3NcUz0VS4uSdWpTd2FZ3ljpw3zlaN+Ycy0uCUpaS3W7Vs+XB/D1k9AEPYGh0nLwhYsd43mfokW
WQ5tBgJWMgpFITjIasLmRotaY1QqDOX3DITUthdh2nEYA7WVK/OYCGMk6Gyv1Zz6agCd5VfUkXnn
Pxhe2NXhOpzxbSv9BctxrV8vDyXhh7S/UPF8eicI5gs8WhyA8f6EMmDz0g7Eoxs6n+Ubok9zyc5V
BRLC9tnYBhPZFp3IaehWA1OGY0K7h1VZael+gEks8DaB8p3Ul/CKHhM/nS7rYT1lrbAkTtbzH/4U
OkUczUgifbt/GbMouq0nXGinMAxO6bwdLZT47BeYO8XQU5DzVxDTehZky+ON27VPdTx7rCaT2wvl
zQdB/5inO+eW8arvlI4HWOHAZ8cfjhttQWkSXFzVC3exg9gBe9WxmavRlp8jJJjbYqLn65djJ/Wn
IPuPRiVcPEYC/NfG+8VdvBR4dTQJVCuNtsYxkYpiN+5IHaWXNfE+xcC5jkt+Z0i95GSG9sdU9xDW
w1dUFVDFFcFeWkASl+19H06Ow812D6vcbvXtHIyP9au82eAJL0Umz5DfzIQ8zudvndDGOuWCfxLZ
MSPejf36FNVTWVUNo2T2E7yp6IBsKT5GcX+2FhZRzLCMNI+zhrbyYA/sS6OhgCkHB4nQFAlSk9U4
gBMq5JdWIOUdyAmOBEAhJRuAabiU7qAfKomHtAzHfXewUVaJMFJKazdY0L7AE/z/R15rlT9eCZng
appCYM8WOU5QSDL8GaZA8QYDtUgWGK5/3TC9wkYVlEH2BlDKWNNAo67N7V1RBsaQDnsdkx7Z/ZnY
NReRMIK4Bi7HpZQkUSq3ko5DOZVj9FJYjM8i0OreiNXt+lz4xVGnLMdYtckH7UNIEVch2H5ghmdy
aBB5geAdN7wQU0Hg8f8T648FXNKFddOzY8FTKmg2VLxeMRJ3lHdlPYdHHWFzok8WVCnV/9DJslP7
am7emZ4UlpK6NAT9aQU9T83SQsL6CxKxeh4I/nFMQirNtZuxByMo8KFj7cLc0ieugNUDl0tqM2N/
FxFu1BuW1AWLOY0d9tRlWa8QaEj7TVWcYEi1O9lCJ39zQT7JBuJe/uZRYKMLmh8xOKFHZRTXZJiv
AxVhG5Ib3v/iNMybY8HY6dfKQSK0OmRPwGTJ+5Drcv/ue9nu7G3ncdgKHdq2hKPsLvA8xCW6VBiH
6uodrlda6vqJ6/Jo7VEp3jR/4H5hO4Fz4qJnzW3awZUuJvfpO/xmBQIutnTH5f/lYGaAt/yTRIAL
NcfA+/D4kNVbebljbAdlPFUX7TG46SbC0zaGGvEMPfYkUVC8Q9liHY82Tb3ItWflIpD7VQthZpOV
d8e0GWI5/3Px2npurPQdbMEYQFr3XUzLNZo7SWmJsToKQwrnQy+9SMl089gOFAMtY4Lr3GIb1qDV
jHixSa5k1PNQDm9fRmfU2rozFHHJ94Jbyu84h8IW8F92+ZeP4qhQEOOqX44/aYOLj0kv99jXxmtK
1o//r6uFomr2PtV+T1KKtXkUEGpUTmIcraUBH1eCiKsgvPddO6u3RTVl7sIppE3PSu+udlCyPsPe
jCV6gbYvk8yTMH9Y04yg995aLXaej6DpMseBOLB+Lb5NWkUDXpvCR3MzFEsLwgyuSY0RSrJ20cz3
ed3a7Um+O/jNr81NrhEoyu+5k+8osbYfiAmlx2cIZhE6cToynOBvWoxNWSDC/fOvyDuSgNQ2Lqwt
FUC7YFYMcf7Ci7IGln2z2HoysYDn96/zq3u5WY+AesOQObSUgWQ0Y8/NxUdmd+52ljcNkeUD3Hmh
McG2j6XV5Yq+2ngM7N/EyX2FRP73rP/pUoB7qofAr9iEh+qEI8TJR0R9JfIvkogiXpHGzp/HlZYX
jmXGfbvvMTySC220qJtYP+aN0T3iRK6K0cUyy3hufZlkCE8tHxQmOmMcPR/N9SGWGEt0JERkkXMX
xdQoeufUZNdiCzbgslzlJVCYqsK2fqtOWXc/LVHS/4Y6AbfHtMMEqVwmNSwKbF5ruVa4M63l2Ht9
pSHL8p6/pKfAI6cwFcnlGufS9zs3q9PYLE9f9kspopwj9N9zwOWM7UteDsWDDPkhSLA4j+ngY+8j
2OvcJ0XA0apzHZIljzBKI/UbZMd4YiENyXiqWyIGkW2B8j8pLWOFv62/fYRD+Rl1Mt45R+mqx7Yo
e3PkocJhmCOAMHAEW0aJ2lkKSzMnaHhqrdhOofeqIzZjw5jfZ62EtpGi18nfMDQfCvyzjHcVXfb1
8fCBT69tCX3saXOHNLc1i5xr46Eniv4u3f5ccrGcx7gOxy6HCsJQ78HBzgHfHybx1V4GH/IlSEWj
2gwvaWLIpYFVzy76RBS99Myc0soCS0YnTLCjPBDN/Jlgjb+JPEfX9HJSihMp1u+WQmTBNiawRwTg
T0TFvpLRlKRIIxoSAGpezWS5AOEuivo5CYZmj71LxKrsp6CWFErDUW+f9OOaNtZSWseuDc1Ry9+l
52ojkTSBaSQ4CRVRRUopvmg7icIfzxzXDUs9pGczwxvAcXg8meNJUdcomqcviyYQ4khR24wy5bYt
FHWMuArVuo3ElCPA+v9iaILT8PMTL4sgoMQR3BNiUSzJUDmurdUAihG4T+SQxdJcGBEJA9wZaXvi
lr8HtabSPD4G2OflK4un7oQMSB3r4nIbdxwuhKaR4JWmpPrHb0jsV6UT0kg4MwCsEIh1K05cMUsR
hHF8DOOrezsicj4XMWqi/pY6JaLMsWSFYGKs5KBjKczwQIGqD7fHiXumw+YFgURU5Lzec0T4i6ka
KLAkXHoNw36gG7p4gEt9mm8XqsN79tvOybO4BiB5EY/3kKqDU3eLk9Eq6SPnK9ebg74YPp4iGCGg
YM3DuzhHx31i0A8MHmOe1TRGOyKiQF5y6fHQBkdvuTtTd1SXyci7b1q/L0pcdSNwV1ktnMUL0lji
y5+WbsEt6svWu/9VwlSXfkgO6MDVzq8LETqC7LYYh9nVqOdrRkZVfQ3OysanfRNcJLz9w+TSyZOn
6C8RxzHZqfyYCXMx+/RU4YIMkwcVGaN8KhLLeuHSsKhiuHZYpNuFOXz+/SQtgR82h7Q8o0u7FWqT
W411DcT/MGIUriaDXvIs/jx1EJEpmdqdlV9RqX2K8XYCvwaF/s30PJFQPvHe2K6GhbGedKTdIllF
bUzyqf2QaPz+wpxCaUN+XH65q3+8+f0bkp1bwhkrFzwh3ZllEvEowxEid8v+OiMUpPZL+HohQXje
bmf/ZeOM6n+TcQizBfk0zYObUkL+MABHPDVivy8VY6CoInESPL4VVUoUD2SKAogHnsl4EpWHzMe7
VpWCSiUQf9S1331UeG464sAKFF8HuqMUdiX1wQXfHEUz7BalPMuTHFysPPvpxxNNVintOtyXy1uO
8OSscmDWALV2q52bx1HJiZ/wT+iRqA11zV5gN5+VaSS+JQvuroWeHBvC6fXXdy9ocMzwFU9sTqbk
BLNsBWsoiFoe0tkZseha0hCQKTzfMhXxyn6OGeJrSYiQkvRUq01V8R5A49exS7bQLD3cZZUQkrPH
TVuwrK/hqk6NJ5WKUdJ6ennxA7E6fAwHCfE/SPiGwtlaWS3AC/Gjlmu+V0YImiSPSMHjkCZB5lfW
M9zCqPwPc9jeP1jvj/w96l46QWPodxM6wsZ/8xmSCgfnxaeqoWBWpfnF9i2cOnsvaM04JpWYIa7A
Fcdcsu1mZ7Zp8rkTjMIDyjdBPDRKYpWZOrhxC681jeYzhGbb9LXRA38+2VcpBQ2woUN0qIasppDa
VCJBGUZXHwYfF/VqeYG8tBH9MaEOhBgMG8RGJdk2oGwYs550E/5AumgOM8jkkrfAyBolw54QrVN1
EaSdF2u0WX8neeYTXwqsH+bGYbxHxny3ki6CKAaqu+iwO/QRDq/V0GEYsN39bGlzEQ538dyB+7wc
3rDK4TM3AkOc0ngZnllpcp9DGLBXt9QBosi4DPAZG9pk8YL67VgpQjvLtzFxJTMX9dYA+B2nwtwk
SoHYrDRxv1B4EkEI5Ysl1SjHdMKKNiCGQkL6obbF6imMKhsyMaT2jNjW6mwg7m72uR9PEhJCjOmW
3INflRMgevqlDK5ognaQIO2hcCw/Heg1HlpySZN4OP97PvQdHiDigE8dtMubiJiv8f2QLHBDNVKA
vcLXCv/9xAq01V6BLZe3xIuR3nMeWOQUuxcMko+NdE8dDxT5H7oRStB88UNUdeKHnFIUlmBoZ7GF
DdhCXYDAIvpi3zJUvZRz01UDacKKHNSxGMnXUqZ25FtAhZbvu109wUDrtd6L1b+GNP2p6Ei7n8Tl
re0Y9X/Ga3fP3LLiqnEFZXXiDsLHm0zuWGM5fjMgFYNuSV6j2ri0uV4QouVH2EmU4+SgMtV7QnHM
hhlhlNOSLMgp8VleGK/B747G0bg2L9inMBYv0kuzBQxi63CQDoSzOb568bUO0pInZaX4bkbcfXCd
EkWzZfqlWFrHTs2b91D2aT48J6gf/oc7HMcg7wgNb2cdLVDl1J+igesG6H2BvQOMpb3QlWJIKiAX
zgEn/D/4t0si5Zu9AAfGI7VJ6DXOWfDSNi66KQBLykY2r8Bo00rr27CgOzwdeOuzEXc1xPPXW7hp
0G2HB4QVyz5EOgFIYPcg/qM8z5LCm2f8LhhU2C7X7ck47TbTqtOh3VYuNqGB0ClZBI9z8xe2wZYA
XOC/ZNZ7loGwyxfbLs5XkUAEsRk2DEPO0y+U2UQRGsmx+7ygkfm66/CzTkB+i6FRIMKg4qCf/qSz
E4RrZMy0EJlIbdWs1AsSCh9dJBZHmlGfLQR+AeOtqK/5R7k8NdYbQ3FJSS9FdhQIGgxYXhJKGpgl
90C9mujgqguG1q7bWNu4aSVCDlCqmlSwJtubrUeUDt6LSrA3cKZiOm2Q58/IjgaCpDuWhslMe6Hk
BmGDk/eeAAzKQynM5jJB56vS4AZtiINn6amfGyqbDvISXdLuh8+6Y2QSYrhmowlLLlYuxXG9e5ss
CGoYcdyUWMKtf82XY1G0vRLLcJM/Vx+k8UFXvIXR1AwUsCh1zLHqMgbifdEG4dcNQw6RxKd3mXOV
o9a9za4kYEIHe2Y78KmGxpJlTqVPqr3lzAbQWPC1OhWilFGfRFrAWh8saA0qOMQglk+o2NMP4pa/
GG5efACuUusqAlR3czcu4e3vWt0OsgfmwIctDt4adOUHBervoEUeEffq2MziHaOPE2zJ4OfEMPCx
gkORaWOoSdCJfCjsp1Z29Av7EANV7AYcHLKK34rAx8SB0dix4ow2MpvBhGqxmpGGxcLPt1AmT3ky
Y4SCnVGBS2duYGMJvaFV22o2NIYg5e96sxagzj8IRQCk9cPxcaqATXmXT6CQ+Z83JmfK/7Danp3Z
jckdhw6DvyvgPrWPRvczsOvBRdYI0wf9w4wnfmr0GI3M26EaAP4hfT0cGN+KU3FJtSynS1YbhNVn
WFPzX1aeVfc6iNKn8m5Ya1RzLB99a63xbhfc70VHNo/6z22yMbl60M2RfEa4AIxapwOGaGFtooij
eLSi1IMz9VxB9UTJdOHBp+Hu0TB2CqC3DVR7ZuXx1XRWBXyI8uU3AN7n9J4b69YFVuOLkDaLWAlP
mcIsm5QWfa9au3aW7t6mxFp4INTDU/6/NTsz0+cOY8/Jq67Qyc8ysnm6kzsyJIgjLinI3381jYOw
RcQQfkA21uf7/IlM6Zrn1+l7QlqvKt5kP45cN3HPmcp5Ce/w05we+fsV3Fm1kVgrWGc4XbbmeZlD
wTF7LSuL8guxv64QZoNQnpsTkTpsO5zoxKnZUogpC4+De2tXueUJi1qxcZp7wI9j7rCSbcf0HmJ1
7Pdab6lYr+wm34h4yuOIhWlHSZHu6X1HMTEoKdUEqc/XKdytXdWFPNi3LH4g1gq45M8iF+N1U1LO
judFRAlgEAfnvqMomGrYHXUkOCI/FQrKtXJcH76m07B1s8SG4EfKfkrxg3T71DZqjW+ZU/eD/0ng
tMkdM6uhwMknfixs3YZwCyrgg3uHJt71vpy05w6Vnkmx+u3QsqMTMpE6+royxQbT7OSU8N8blmUp
IJrLc+0OCXmSNg/zJ34W10HuCr/2yVUl6+BxWByfzEwerGDiGc+/K4Iu0NTFLN2Jwz+kwrywG75o
peyC7zzU6pG5RgtC+Z2Caf3gb972AY5Jr99GbG04B+qtedDXmVzGU/YZdk6P1gHbqU3NN1AlzGgi
laGXSwn+BV1bQ5MAS0nYMTgwz7JsPeZI8OoK2ioEkeoyJPa4nqSgBZ7N7UF2UV15vS/XBOVkmiEC
nQJCtEvlJ/mCHetJPxhRSnWO8HSAVGBEsUzQDsY2FjU5nc2Hpktrs2YXVp0uwBjnHkTgB+5QbAaG
eb7wTG10jxZ/u+KNG6ix/HcnMcza97ODUbnK4f8lq/WWxE8LLDRFAE77gOaVYpeK6rts/FGainYk
xXFNWMbTN4X7UPkjcjBCvcsKsQnfthbrQ6786ON8fzqSJYxv8Z32wo8GoBo7fHhlw5uvpq17ZZPe
jGmmPm8AQtktDkaZyztqB/Ha/+KbLfiQ8cgT0rA8n+6oT50oBUGiV0L8bi/fUyYhNFb3VGqE7yxN
Jk7bIj7c91npyrjJSLXC0enPBGj8KWe5qQn0JA8ZeFoO+RPkeqIl2LMDleYdhUhzbsavHaHEccbJ
edmpqkGwspPcBBXj9SIwsLNLJ5li5iYHJaNtc6Q1/ZDIXQyPEudxI2U5J/w27dzh0hiSn7nD2zw3
Myle9UloJ1Hk6RhPvGHU5hbPR45nFk/aTS50kwhk8+I68omCIyO7wOsK68+82klQAk3KFS47GVHt
+Vt7T18Xl8G5/LqJW53Nc5MfcwJcO/nVEkLwbkTZfK9XJ56t66uhF82Dt11u8GuzWgqUyuxcop7K
Xpqe8wnFxe8t2g4TYlHltQoaislFO22F78dKP2/Qm7MQAUL7L4EYkLpvxGP34jW1mQY0glhnp0EK
QS00XzsndYtCbTqMYdDY0iCb+ccLpa0x6ToSTKl1c0azSsA1TS4GATGOQswiNoHCrEyGbK3f/VP8
+cayFUjp8Ezck4c+YkVTWIzF3DkETVrc6QRYWGM96fqmcGuKBWP/lCrn3WCr7qPnc7qNVFKoBHk4
GfbKo0UtgccoT4xMhT3ks50Gg3VZAUfwjEmbql3vjQ2if0w2piUMds3CthFM2wKWkksL27w8Bjcn
K2qc+aOlgHIa046cXECnLwpMInYZaiFz/EMDBg6hrqpgzJtpEOFcmcK3/p03tGVQl5Rw32969oNx
ur3rRCRB+GgAiCoqWEWvAny+KpsCsW91RMAhwg8lipnkg530VkxRT8laumggamOa0mGbwMn9384n
KZDD2fMyYEvYYFrawCOfTlOdLqIEe2kX7avmVKE1FhbRuAOLCMlla/gBct6eImoePY7MSdca6Vyu
keWWf5LKe9YCzIofRXYeFCT0UJPZofvDS/+nnOZJlHKDi/79T9HLKKZYjAbCKMbjP/UJTpqEbIUy
P5JXvsvGygF0xsiCYwiyL5mQmFnJT65lLDplNiVuRtUp8xg4kW9dHoizFRpM03/sXhXmW/aPOb3P
vGO8aklqNbnz53Si5FuBDHJu3n3YavQoXnft0bibss7xVhqZQwkmGSQoqjnaTKrVj8jT2cSQpEY8
4wgS5ZaOkzlf4Q6AXnXed9PyAOefZnYtNrRLJMeZD3YVrzqdFs/PzcGZ6ZIlug2trArFK4K+u+Bv
+7F2riW3VuWbG0c9M/4Add09mF/KgyF1mO9dRH/uO7pBEKnfvEf4XjBlgPzGNz2NjXvxIbYdM+7a
22JGgBLcdBA0hITSYMl5oiz+pZgz4HA7B+yF+9WL/Jc3OsPfGR9a9AFWHH40njfxhD0RVGUG+7Oo
tD0R8j0BcyeqUwvZcRVoV1pVH28euY8gmzKaCM3mPMCFPFUM8p4+CsRClzhAH/BEQGmdJADxJ+Dq
A5PDqX+pyjQKvby2N9BHel4oZwaQAe2AllGX5eL/HcSpihYwNt+MutJhj8Kk4vFlgad8ntHpQZ/k
HGUV5fSIOR1jMrPW7/jqgULqr9xCbQix7yQgMj3LURZDIDJ7O1o9vVkEtY2ndrfu+fTVhz3tyJdg
omu/j//Pj6Jvv1OuuYBMM/RD0OypJmnL6ZnmqF8U7IESmftZ1mxXr9OVyRJww51XaBjcu59HwkRz
ctuXoYnrwM1kzkTRKxAIqnSeJD8ndd0/0Cx15vkAK/k4ASper0s5ITkiNF9CQnj7QhUvzpS4dmZ5
kZ4sY3//8cEZmk8asF0x1FtszpGlKN9EScg33EUmGyUwz2qaTJwIi+4GnDWv7R6BY10uUvHrmSZl
c8mPZb+IIFF5/usdbsC3Qbu7nVtKsQcPw0vGC2FEe/+Dh4OUNmEiSprrZJFCzl+OkXFcmtDkX6oD
MT/1NDARQZY3YjWikk4A3fAXQvjM7Y3jEbOztIp20hG9SDBUUVM072C8R9Vg/w1u/iYEM7zxR0RP
pDeIKmXEd/F3xo3kwtvZmtPzRlTfz/35yYA3PDTWeFoJXWG1kky3jfu8mIZLt3I74B28ZNiJmjqv
MUgcWvD4WIt5gxzRgjg/jceO9YWUk5AaQoMiH6PuPHLEhTZ0glSpQHMJv9ax2JbrakvKE1vws8Hq
1cD0LRiseWvATo11esrdLvJtqkUu3KbeSVVmEjibuYIWUk+jCBxDijtpMZeefcaGyDRaHXepXTxq
ipclV82OtkqPpyIR5k84E/Al5bHqlA9VIh6DGH9Js2XZEkA490DGwB40JYWvlWlNzKPTDpcwNelo
Zfqq/WsmqEf9c9Q+FNU+AHjA/s/6brBbrjKKQ4O9CRMaxKIBCbjn3mSMNzJ5K+ny6PQ9V0G/cDxz
A/mg+p6gidlDk0urpq7kPsGO+gXq/SYC0SD/Ybm0g/tD88OjjwGMaSifsBMay1tNb5QcOgnWM1CH
b3iiIaxIhU7ZLYI+gmXGyyOVfQBNabe294qEqRTNRBXJisXX/5hKNqEjrJsjJ+zMuy9bJiO1AbWg
LweIjuD3Ko1XgEFvSLdkQPG54L0wdXFLxsiggkPLYGunIXnVKYr76H95MQ6s+sPEEvXkySBHaEzf
Cc0ZR2gnUxhpPh7FqKZebOell+Gkz4lBeJDuqom8k9gXFXLUupoxeqLnI5khqX+T4mpa+W+bseXB
9qkB+Cd1vR/iSmx8K+lI05ZufMknuowW3H4uG2eKR2n5TL7qZDMSN+ipYCkScelDlNwZF011ea0o
NicWuZa/fB9eI2z9/QK2bTAOFQfnJ4b3k/wmyf512UW2G/NMEREZ1RBmZWus9sQq4HdUAPf1DBO/
noJcALJBMTxxp96GeQNy9tkBynEnTrX/s3o8pTRTHW8kr5ci6GkxPSujX0/J37u1rBUuhQOssk38
K5hZDh2cr2UTrINDho7wsaAMcu/w0gzET5Jh89+cjrvw2dT+jNPgykGvkW+G368i8woA3+I/B1f3
k0WZH52CsfWwbq1kPQnBQdkkLYPR/IFLBfT8h3PaasBuBk3FhXmxLEk8R7gMxjKPqc9hGnYFKKnP
udktr8Jx0Eap/e+qwG0jphCn33u0NRs0duQDdqCqAD74PZ9SxfcmzW81p3TuIAFoXFMDLM9tEtz3
vob+zHZ0eMa10zQsKFX+UJGCCnylPIwkU7M3E0BRCoR4ZEzGMtRDytJL1bCasILN0lbFkAcilDxi
DtPv1pjzaADB/FEizJfKjydvULAE04ILp7bjcgPC7mJNMP4ikh3flVgTtDN32G74YKesr1Eye/9w
QxcbLy5qWMSlQt3AnNPlDHbHa/+imSAyx4W9+Q1qYPkskh6vzJ/66dnw1SqpNxZzt7l+zRl510+R
ixtwCl+/GQ+MM4AXWY0hpwUEJQYYsMBzMnRJRMyNhx4JVWQJHSdkpMLTKXd0kBYm4zUpRFe0O0YT
LQQEWZRDcrp4d4nDNQmYP4lvvD2hVwtRCb2oCM30Z2bOQm3EdGyUYYdVaMtUZhsee6XDQVQRNcYj
gaQOIyZ7T6C9fEK8KFXZatL4V4dUFR7kxOfVViesdggGpNB2OlySiy0PIBI/Dghg4AMuFg77Dl3k
/bnikcTyx7X4xH0GUIqkH8G4r3+DxgWDiOsdZODGlk1tDTDuHTyOo07yKQUSlrTaLyy+a/3hjHRW
uh7voIBxMyxZfwr1hzLSsuvg0mY90WVb/A+fnYkhqPEJ2EiWSXfVYAMBroxZogU5oTqR7gYeGbiJ
q9rf5k85MErmq7QRj709oPW8J4ZOsURLAFuwm2tpX0hUYTjgdSzVBXOUHXWTqml57PvMc3zp7lR+
mK7EfER857nMFA9WIQ8r2gPRHJZKKVtIr2KDU26ZDFzfNzvcxqOSMIR6dOQaznEJGQYnQPzj6qnR
/TFHKG0regoX8naP29HaPbQbu5d8gAMygZyV8WPGCMTwk/Z+twIeUAbZ16XMPeivFObKN9OAqwAk
Y7ah4lC10vqJMEPHpsNvPCJY+d7WANNIvuDdw+Vju9FxkXx/4veEWuaD6w2gYDenDUcMP4BZGD95
GLyz3TnSuXb9AWR1+3sJ4sGxZSbaYbQ8mZUfhZS4sJ80oYpNtsqrQoidV78PaMvHi3NguCyjnjxj
NKm7CP0Dbbqzgp/QexqutB59FdWqkHy7ybkfv0b65ByyPxMm4GxNDIrLtVlIWLBBvFq7xFrVsPiX
ufEgy/I+s2raHInm+WuEEFJEWwDWwT7DbOQvs154pekeZDnD/iZZwbcCdKMePdLCVMLL80h1LwvM
D/xXR49XsaFYKDCy+AWLNN6vhkM37MSyVCoiEctBCZTod8Q1vEqyV4/dgOi+fASoaevMc8uojgTf
35MT9d0HYxV0kvHpnFsAsndstYO5AGHCqRMbp047wNEA2H4mqmSme8dMWlM26shwmJAlCu3iji78
oFNEZEFXBVyIplUq7yXIckHg40Jbhc2ZSJjwf1FbR38lWyaP0gkrZ+bYEDCyT8ReHO0tkBszZku9
wqNX3y1k8W67TB+F/iZBTM0ak1vht6y5vbXLUNLvIYNVmBcB3CO7h7hMCPGPrYZ35rAQkn/asQCV
MiYeofVklhtBYsAeIa8iq9fNqwBoSUHYRu3go8cQlutpGShtjLrtOXm51+bDpNZegATO044ggNrD
XPnBBYWmUvMLQLNONxLgcyTPky+oxbgZ8gHz+xFr8UdlKyWPSt3WjcfrhfB12Lgx727Za2ctUQV7
tAOxkIPEg0Rbx2bAmLwCEusUtcuwORsV41rU3nJv+x6m1n0qxpHuqisZI3M7pUut6K3M1wEGhsE/
JvQVrW8UtAjGJfsgSDTmI2w+I5m1goWFVh+7vDH3jbCzEd71glxMxl1Ibw8rtVocNb9+bl6JqfOj
cx/TwoAlf5fol7mcc5m8N2upGffn0fYcyMTpwBnMjl+O7JB8EZBwcWRgBRlHvwLDxpZVU4Kw1AeP
R1pYDeJ/NMkMMMf7TDbfTOkunsR85j0k/dKzM/5i7ud7XJoC5ZMxfp2yZCs8RF7++6YBUElN2xjA
CLGLGRKiIL3nLxhjIuQ1afYbdD4sNwVcjm3VfpL6SLrlVaUVwyi3EaBUiA2cluDIe0DuvF0iCeag
UyM20qwdUoSxPfU4vK9UA9qF/JM/wn7YR2nzW3f9YLDvxpgG+FAlCP97HqVuactqzm7DsbZymFDl
B9C1IkLfSn1CUO3Ve8WS/ZGQZZ6T8UZJhfmXdcGeDeXFpQ4CEW4/bKWDmdasc5pmSK/nV/pTAzGc
Kji3sdcT/biOLZ/L4G+HbBpVWusWSlZ7JwVsIIxdvleUgqP+uI4fUKS3Gdaqz9Jds6HoRElk9tUR
dSv5Bx7/GpOCaZfU6qjHuuqAWulNv99yx0dr1fxFBz8zhSY1c/pL4rYvS5mh2xeuZOBKcOKrwZEl
tZK8PO0JClX7/UxplG7+bZfNYcVUj9pHzQ0T+3glTX2G3+dsPcxdKEGEJENBYq7pQGe7/iBsjqS3
qukRI5PSkzquJMJJEj0dN5wayLY+F5udwXxMU8/LIMguQx9HGtKwqhj0vRH6KCccNyl+t0n6SNfe
Cq0F1Vm3uPuZe+0MDGUrla1YbODa+koMgsb35qpWKtnG++nBQIdE5U5QLSvtySIMKefkTLGPtxGU
x8Ym3+TaI/PcdPBn2yahBGXUPDZ4erh2FJoaW9me+UPkLxLidDBRTpMBL1Ox71u2VVoc75NRXa5i
QO27PELRrcLjZKmEDhAfI12OJ80FEO8TVxBu9CMtIrxyxasKd5uNhW09UYKZqMLSJYzebN3mGQMi
Z0eTMgLpgPHxzEv78gbep3Li7+IdFVNRUndeQv2qBQoyiS/iEagL2O/CWdslKtw6fD31sRWXKEuJ
JQtoilN9kKSYQvfc66+hI2OG3QrB0b3NRR4rRI0S55BWkWp5xzvRt6Z6x39pIt1Y4Hdsfeftn9jI
xSF/VglAt6spX6TFhSh0EgW1of/6MGsLeU/+VSQLuIKB+KVgI/bkftEcnqNUNhsvpylOYAFU7KYy
akAbCeU4/kiksTVquCh3VH7/2qbZj8KWXvqJDph2hfAu1NLQzKcdCQb2i1dQRA4ZcY9VwSt3fbTB
DhrnI1RvH2RQffH+dy7od489xrV8NI6Oz30vNBAKJV65vt2T2rHBDvHlVDEIErQ6UoEvzRkBM2jv
rufG2TARm6x+BUHQdTyYnsGzJDASAEdo8MiPL9meBFQWRBv25a77+RZLAzu0Ep6VBOl5MdP8GtHo
P7WB/U5qNAsNnTSFyfrXFQBUbJ8IsIyEoqz3LbnOvFHVyWtwypLSEMVFmB7wc8mxM761c/lS4quc
ZyDHHMNBayYzhHxWur3VZJsQVBHsg7Z0j0nHlqZZ1Pyra66EIyhYH8LNmCuRu5zRNn1l844l64ea
zv+qPQ8SFmF5ncGsjimNAt+JRp2bHa8J+6CYp3PKAtjjhse64jUNikxGFXWfWZrwF3uSpHO9MgD4
nQafJozlDy6F1cFe0ihrxXPULUC7SQZiRlUv7OidOL45iHhFzCIwNQKoU/UQkzmKow8E7m/On7iv
AlHLTFy0/IwBhMm9i6p27lMeq2i4pIWs+85HJXo0Oov7WZs0l7fp9xzACimNLPJs32FEWdwKv5iu
l6lnabx7DlaFHBhpQt/9WTAViPCC6WUS6jKNcHH6cxR/DORpYE1FpFc4lVc4UNasoXLMaFW47qOy
iJlcAuYH98cjJQcCYT8g6TIUId3XO+ZsL7HsTx2QmZbcBONVWsyCryp9v+bqv9NCvEuJ3ra4R0M+
1JHpAT4Ws4exvlznmqj6Y0Ir2gfoZNU0JcgECUaYI55WN7Vbaw8VKZcu1Wz1M1l2wV9f3cvh7027
KiDSd3qHXF07cwbkKJhdrtxOr8p6RMxGdBVhGt4xlZIrWi/anpHxzuXWB/RYGs64jMpJlBNo30Rq
jFkSRH4sCehgH4wnWYEVhg4Jsd372lvSY7xt8u7szm/69AMmalPzJMzsKfos0HRe5C1aK4f4zrZp
J5Fb64zrf41zxdxf49gwgBnj3nG9mtnfKD/zPmx8AUBhXxiQdYF2VfEWkMRhNwHUy6u3RG1rfJzZ
lfgMZF19OrOC6koL7wDOyXHsLZlbayvvGL/YDJoIOWM1bHEkml09b7fSH58+RKCb9ApTQMq7Yr3f
NVwJWJMZtZFqTtW++Z9Vawxiz0QiZV3XVDL/dUnfnxbtLeAzaVUnS/LnBDHOe9V2ixELRMVpFauy
bmy2O6v4YeeNCc0HogAHt6m6cA2N1yyPbsu8cPIhCXTjesTwanlx9zgnfilKVg3W9Y4ufuZcR7uL
pJdg/ftFLXZqf4P/Rr7ythmm3C/tJdzB24DKPasz5GFjUEyPDJN8X1BJpTUSF5hBfZDfpp9/yL1l
1jEg1PaddAW9Nat08oVs/E10Bi7o0Vwu5gyPLFgEhVYeEz4ynjGMWlLk7fG+knau8UtfTJgaC50P
E4DyR1D+bgMFI6Ciz+SRram3pgOnXbPPQ27XPZSiHK00oXtAa5mcVoe++nSIfbwOOf8lqfwfXbbH
rmVgI2TzLvL4FtXmO3u8hKsmd17Oaiibjp9tBbtHBavie6OSyNli82cm6BSXRfwsxsf/cl5ly+m7
M4oiIj+nEnOSGcswW5Reic5RmcG130jsSGyWdjIKj6fHjAHOXiOPlRV93GEqsl6sPqCccxy+AdBn
xgKqgZygNtBCVvi7U/ETagMjq6dRTNS5E/q3YpArWI+InpUNvTi6sF8SDAb24GnSg0Wsbdod8VrC
Ut6v08UMy6Uaoh+67LU9SpOwK8dd3cDIF7FN7ZqKwikdynu0fXo57mhHoassVibP4P2ElijL/4Gc
ZDdtGwGljyLG5QWB+QU3beiVaSD7XO+5SPMcWR+LlZWk+PH1UMVowubYxS0JUkXRpi+iSSIq0oow
GeAXcL8DOSlmFK+t9RgP9iUEuOePQ4MjyEg5LA29IlyQwGVP8hIuJXIEWGvMCWgFo7jILwuwCyS3
QsaI71ilmed9VNtrlLfnCjX71IAEoXOMMK4zuefA1V290pBay/NMuCD+wBxDp8vzayEHX7x9F0gv
3S1tttUhzw+4WuaH6BiAAf1gcgGyz0TZRbBRJZEfUarNo6vl/OAYJG5Bh93hs263dkc8nVybqE+B
s2uD6WEsxpfd09t19kXohdC/trOW8dmI7BBpVMPzUkg1KeIdthp6xvSQ2ILd45JqHWwd7M68wrgG
vUAbarl8lo58/DBVsj3sfkbtJQTPEUy0yLw1xoWRKZdqnNuj3TO57NBkmWADbGFfYB0uHSg5g02D
B7nFHdLmiAwMg8rFj4duH8Vfrc8lgQeMnNqeXN2DOYN3FCbng2ygsbnP+KMuXaXRKFaH2WCv1vq+
JCQ2JqZKQfit35j2niWPj7fI/JAF9kjIo4orbEOjDOP3QYQ1vrQOC+imRS0mTqXOh6Xe2SYw4PNf
ek3dFXjKuXsN65hwV+ki22E4OsFAk4zqdRkAMMHZ8oG8riG5k8NgIhPK3U7xFiC28RssOJOLkYZ1
L7xfLDAolMIcukrcLkhYYnkpIffMiq63/2qIDvN9BB5z3XQKGi3IyRPXYL9TPx8xg4OC6ltLEsLc
3PdgtEfb/TfKhKHNP+P8qqzaqJG1DSFl3Kbr4Aa8KfUMoDyxs5oOMqrSnxjHJyEzBnn6eMMiCZAB
pMHUmeoiw8FI6la/BOxdABPsWmGzQpPIvgNNm61A7e1W5tApLHzvkmKuwqPd9UQ8Mp1sGTA/uz63
hEy9j36f0gKFiSsoXuZ8EOSgePVSEmELdwZdRYYRKLgaRsacy3CGO7cj/2xKJjzxo/aMue0s+VKi
glOxTfBHwrozI3g+GKIdWuNgntbK1IpuGwMhAcipuXarJCmdbb6yVPOVtY1RmOlLPJ68E+4VPi51
sNTE/XxU2TWGGpm/rQ4n0WTdXt9PBT9RoClCAnucjFby0VirMcgcHDzZhlCPPSXL4vAkLboUvjaN
N0zJgmAR5SsxOLdjHM/4dJW1++zhV5NMMIK2A89IHEJqUzFii9k22B6PUO5B1oeMcHyD3L6lBcxh
J6I1j8Z+tBfszkPWBZoHIbdz7pXAgNvyCwvEHYKGlt02xY2uYwmJ0Cttytpd6cEjSu+J5I8rkV+b
d57bSWWE/K3j/8kKuvnJNMLrj83eoUv6Toius5AouwuzfA2XiCe3T4tQ6ZJz2J3MKOzqYOQ0UMVQ
G4c3QSiyMKr/YWQ2Gw91XgHaDK4XlPMaKeMC22XESunfwxHQrjGtLIbU2VymlRUxi7AVbEdj4kfk
Nu3jGn5EHlK0fC2IqkyDngEslMExQjKSTVppSxNISybzwd8rRKrNcyLXAITwxuWNgdv40D6vv6PE
coMJgZgepZo0FlZURD/sD+g2I/T1SP831y+KhmDJXDijNgAdrngJXG3C2IQKAntPv/RVG9ob7yn7
JvxAqv7zY6Y0ywbLoF3B7zirYXRlBrmhDpfF7w5fvdGshaeErNzPVdBCrTVEcXuDezR2rSnqaAgm
eDNadNOXReNYYncQK1u3wY/olK9mpgdy6umHtgsDkEm5KOTr0CmDf/uw+QKIKEA/BbCah7Yw7tWh
VpJ3q/i8iuHjDNZmbBMnob4ui6N+aswG6JapCk5vLeuqv4xAGTzYQKmWEuCLcSduXuunQD42NBi5
bfncrB6Hf00alJvphHUGI9vjSl1N37Xy+N1eCNtWh2bgMcIrjdpC/ohAI6fIb6qs7wSPMYoosPiS
ZTmMUrsoMHneLNK//wr3ertvWRHl1shQl+N96HGWyvoapwIZzmGfe9rtWFyV0QQJ4wK5R2EAVix9
A0jDZs/HXX78Qso+3l/4WqR9NiIXjD5pUqtQ434fRq/SzFoSwARKelgH1WPzSvBuSNaNomcnjz5w
Bx4o256Yj1ZG5csnrlx/Qu8stTVe6yt9J7Y4ZaONeqir9qkLAIMchT1FpWD3EDP1z0Rv/3ZMFKnB
RCZtojCRgoOIPbNTRZi0dUrG3fMJiYQ82ZVmcC/Jid+C0g5PZ24TBPJ8lVYsQvio3GEt5+NeV3G2
uw1/Bnh/4MNJ4d1Og2L+V3EaoiHiN4IS2H9Ac0iVDfJvUGaWyPJyVXiBovmNCfNMZ1euK1yEceFe
p/OIrjMrIonGuglGg0US5Pqnd6SzT4vfwd0SH4WIskoDUgvyCLJ2TCkrxXPT8WxB4mgrb/3EQizk
tfEHUvH77j2+DY8RDtTBfOcFrYmXT9YRaL9xwtHWxQ8fBHt8R72LVLAeITc8nmtPy/wU86sVXM6n
9sFRyPlw5KoGH78QOUIzSTct+ONL+P547rRBn8XOKCX8G9aQsm23isQfgdWsn805ZwTgz/PbQVKU
tfEPCpbRh2ei5H+hMzJXxPzz307HEJJScmt6vwVXHosZVNfcYO7SudPG9FVcT5cVQWXfITp0UeXr
qjOZL17aPywGem6L6PeXFGE/O43sQ1mfUxcm7xNLWuZJbfgA/CNzCuRsZoeoEjMkzuByOnrTaOW2
8RbchkHhgrTBqL/8+Ukd4u6QFJ1TtYGNX1DNDJpV8VXfBH0EVQNHdCdkZX2RvggLHnsnzTd3RWX6
q7IRlO1vKzG4f2Hm92Qyhd0nuddBNlzE7cP1stTJkmBWXUJ3seDPwQCbl7aGF8KBXx7vrtWruXb4
VDL6Iv1RhmuD/dZHGIdHpQql9tmpxTDqO3U70eVnUAuwmBRVBih+crXIW6R5W0k6AHS27k1sNOf7
h8UYpD7rK2byr1cnQiB2NSahQeRUNdr3IX+DiMVM38EE8yW+5mS1SQwbwQQ1T9SUJrxeDXD8tFaU
Sq1aJq6M8NRXfSXOFphX5eSPYVJffUSU7MCE+7aO47LWg4r+jBvWishM6xuK0n/6SwJLMMoxULhZ
EA2JC6ibrpNppAmb837yXy46mXBvokepXiZiJgp35vITubz+1LLQ1aH1zO4GtHWzuM3baJrtD/sf
ZRwHoZwNRRjgQsJanESDyeA09tqRm8rJzM/awO7FzG2bnBg9wZZRu4iqdXNXhBCY9D4u58IGny9+
YAphYCxtEu3BqvyaqqyenWrhfvynsZ7xjekHPDC66vwY708bY8K//f/1vQeTCjtfUfSmMb4qYj42
u9dijhVqNcBCvGF3ceNhGjjSBC92FmbKkuOkzBo+E2RwyNubY4093XwyzM6/s5T4oMmja1Goxa6u
zg2VCSHyp/dgRsyyG8eHM0pE3IZIRPttXG2NwDA3OwMdaJc2FvNIKBQ3GHEtGG7FS+GSKVRK9bC0
EQ/bw9rcISRaVjWpZpnKgGoi6QOyICOf7H6zlRz9p8GHaCHPdQdJuwicWExYqep5p2LM/S/3S2bF
WrPeWmTmUjS0CB/FiYGujHmEHCmbnb/2ynNbYGV/kYKc11QLA84QWgSWmbkF0LMXYkLXOFl6IPmV
d5VtuR9fk04MTjPtPMREU6M8m4yIuBUZyp0PCplEQEAkVPa4v0Ri/5gNJ2KRdnq2vLket+i5Aptq
LlktRJbW2K/4GaEpymv/LpIslpi/uEExNwtA5/UfO8G7cgdjesyv73ZZEnJzi4YW3XzGVyfbRGNW
e9l1GUlLLTL9+kZejbESeKhnPdw6maqCp6S9olETrQLQt7BrqfPhK06LB3eWo5YWiljVHm8iOgQ+
A+tKbQKpz9XzIXAEPkJJ5SaV40qqNR/zvcksruzpUfTIvuvIgP5fHfG5H5K3G6vw7jEZNf1E/hLD
ZUWIJI31YV5sLeRJQWKkbvNku2tWo208HskDCBkGa96QCT+MHKIHd7BNrUx4NznigHz16+0/2E8V
hfzFGfrpKuhTGjkqft7fe+EbHa+RweZmOk71FUyE5zkXzJAboJbWEhWsaXU8uLt3FHszeFib4XPa
l9ZBEIg19tYFsb9aNNdp6ZMsB17SvfUPGZ2CtQ7iWHQcg9Kn+iWBk2gGwaYHpLC5LX2MqMMhsRee
R6vvCmvpKfAA5uagjUDNvXH33Nqjoyi+v+HbQI1xR7LEKePjG2u90IWCZ7dkkct1syzkY4FLF7e8
j8NJnKdgPFZ/PqDd/KjACLfALSbRSKgoGWeMmO/OIl7x9XaY1iNVhWJHL2Ld9OpoJ5LfZqSE/fS4
+NX1h8d7OCOpHGGwfPTAITkrQ5mACUJeyIYyJyGVEl/Ya5gwWjAmIpi31DqmrntferimqXsLIpQq
KdnVq5UXU308pzfYWZnNtToqqQCw1zZiMiQjzJ95bEJKSZtJZqf4p4+F9uTiZx+6K1vhlGeVSFr3
fZzIuaD4DZ6Srm1LmcuO0MiwtArdlFS1GhzbTjHYPj6CFrib7BXaBCXFLernB/HBnYLBarHaaFCA
ebt/rujXqC/XcUAgxtBOlO2sdsIS6q3yvB9BxNlGq6+Bb78Cwj7rOVgN1XcPQ9+45r5IMGP6szru
7zmbM7Bt4/f7oXIJxGQduuMLS14EsjNNCRiwMkNwE816AXITvfVMhT4pDQNol110EsiBonXp8NrF
khX3R/ITRPdrLOrEvvWp+cKw17XPq0eFmwy+SBw8HGooTTS2KVoG0EARmTOTPoBnQDZ337Iyya0h
Bsz8NPT0G1e3win5DabJRuZLKmxHgBJf6jmQ2UPNBPzfzri08T+KNk56B+B+ya3GJ/e+kWg5CWa3
0NsicW3yq/fwvdUL+V0niYu28KV+QehJiNDuz0Y5cnz/KSffbb+oY2M6ioD95RZ5ACN+ZszXItwx
e9Ns1DmyJ6e2GoGJICB3WsJShZNtcCoq3Kja+NoJG/Te/mZlIvVNnWK3MhE/V20MZE2w3cNe49fr
hofw3BiEiGLl7ZlJHaDBVM9SrMtMA/fXBmkUlPl73P9xRd7kqMou6sap8MIehzNViRDg9ivm8Lj7
iV89/wm9w5/xyMTS2Wdnz+p3wlBQsRbtbfxcxugTaLipBIbUpZ1wi27aK19QNdX/E35QE/2fJH0X
nTKr4bpaCP7M3TwWVjhjAr6nbMGk7F2LbFTgBjcL8u/S/y9gbVSa1E3c+F0xlk1vQg0l/BKQinPe
ED5NYKexkBI5smgw4zFO8084X18biCZfuZ76k6bwjIg/fu2NKsO1bxIJNxEXgmTHB0ldYD14UhbG
Un7/rieujjIFJ5TTUKkk+VxoVvsvHo7fdhxm7DCOWk86yhJdlTKGU9KFjnuPo+JFMdYObDVuIcUh
Z9Huu1ojmEJtYDu6DzyC3XeKZQWm0bgPsG22dOzjV/qge6l6LkHak621HcAXwwursjIIdfakEkhH
RPeGzbAY5C268m0EsF/mUoHM3YtnXr0uaEwj2Ig7iKGdt8Y9hOn0877hRQMU9OkzA79Uz1ZUgE2m
L8BNEVMgI78VYyrLmeiYc/b1TT452UqIhIoO65jNQp0jmvvNviOi0IEstLy0c6lUZeCO5ZF72KXt
/iRSSCoUKlRQA9L4PEcz4OYux3KjqKSlWCgwTMAKUWDkoWdfWEo+F1NELsUfBs3qrAqcBVHwWB3F
sF3hXy5vaESUUbCxx+/8uizTXH7/sDzX37IHDMQPXscE6cV/U52zrFbRE4/juJty7+/T+ubMOQyX
qIgPW1s7d17Qy+aYgWIEepi69MMHqqmr9hOFJDpqaGc3ct5sbDxxh+TNcZeJgg3kvh49W6sv7UZG
nfodqJUH/60YIBPXtcsIOICAVRcZOunhv63pIlyH/q6ITqFazLP0NK637DPfRTqIff9cDTlaQkFK
5uojpcXAZwca79QzkCEhAbCW2+ui7Z+mw/79hKZ/OIcRFc2xqdVqfFQW8xtMRNCKj5ht5tibKVXg
/7N2APaibB9aRmSP6Oh6oOIfm5wxC0nEVHdJFh4S72hXut0PNSqFRDC2RY3GKNYiDXNbyTBVOx4v
VBZ/KheED04tgBu0yrvKoZ6gqt4S7f4RS8GJqCXPLiSxHtylQq3eKUYgLP31mYlhino+ZjSvvB9Q
lyvSyHISiyres0cMewyhzhbaGtLVRlLeDwKdD2xbw0Wy6aLwPb/+kCAKkMmkzSJPrsZj+1OhFQLw
xgpeN6/dYPjsVu3PJqNxF5bwgdvIOyFDR2LoMl+7UjUX4uHsgZuxXCybtktNouKiKk8MymUTvAEE
yvyX+SjncP0eK29FRmJozuauzeKzoW6WGEGAzgMiimni9mxsJtEUJl8yf0sFy7nqYbKsomgPQ9y+
zLdHG5VqWVHFzcAWIsY9b6vA6hl7b2YPWv2IF7nDU6hp+KpvZ48y3XIaDQokKG3VBEu++zAPB7dt
bxHXuDEtxtUixJziSTswBbEwgj+qlmXqF/9Wp9y/yVWCO6tDVvbUB3llyAP3Wfp89mgFCTo2366U
vtVgOosx4J0u3PrtQh7g5azXb0jcShHrPAZBkZF6CBE45zE6t2gYfrjRKCqL1lkjWxHhedLQIadZ
AdKKHBDEj8VN86kQkNImw0pfH9vdWoH4Jx6KhSypwzlyNvAgriq/4b/VSyYH3q8dmYI3DcxfRF02
o3yfVe9camdg/XdbhTHMDD6Q0pAX5IQOzBxlb3IpeXRCaIIdTOwaAPSR1FhEIIfDt+K2+h/f+pSO
prFUSzIPcMzSEYzn9Y84V0PQOpDJiA86dLbXxT/474JZgwzEU1xPhJ7ZArpk9qUYV44AznC3reNv
9pSlBZsZwpUumTTb5slGqrBxMFWg0n5b2zMnBFte/FBMfRKXmUcCsseH2mCiyc9XWDaB/LfSQkLM
7Mnic8dODazyECBXZfGtQ984IKCiY4dO5qJ52Swqw45DyihLmEx61aYUdE7gK4ayNfWQj6gF5D2J
4mSBg2jMRDuUa5FQ8FOgXcUegTLKIKFFVtF9poj5vG7o/CvCIaM8F9I2jV/xmLoQqUDusgmuTumX
5m/bXJJ0BghJRm2/AgY5PhKtq4nEQORG5BJroE2monhQY3gDXbIWUrDGdYqy7H7h2eOhoJS8PfjZ
7sGmnivD0Bb3J/v3XER0Dgyl+WDjNfL7z6cGRzIDP16y55a5TUlA2enr4ZHJV3rs8QwBT9oqkmnW
megWR/Gv5fo0ape0yizDWVwHRj46nVt8viWIidSP8DkizB0p2IHpKy3JjtFM2hUCwL4dP0oGU9Xn
bcIsJYR9EA0LFuoo+XuT593TPfkA7Lvpr3Vt/hUgXRK02qwDJD2LBY6qMt5F3fQUouFXGlzLS++3
S9s77D7kSx0terzHHD7XC80XK0bV1W/S7ha9uNZYbVUc3r2ESK+iuOskKK/mA+jCyYi4Imyl2ViY
ON/tKjc65zjIDy61BE4xZEA9hALPgpyMLUBmV12vxJRGsOpDy6wZFxhdEo4e2ZKrZ4iADZu+ZMNk
poeV/IJLwcQUW42zdfvXprbyofrYhb8FC1RxNaWkCcOeP6dw1bs3CBViWyqRWw2TnGYBOfyifKBr
Fr6wCtNK9+7Wl/J9DDQGg36nX+uA/Zs6B5oieltdL93jidn9xvEXNOjlfO6rSsmvlXKWXpz2rX2h
nPTCMcq3ExahMjRV2wwc+EubWlC9R2BNN/8Mobx2VGojt8aw2k1FNGMsOIfZuLRdUb3oi8uNx2WH
I3GYgqd0OLDpxipptNMGyHKDrtGnRTvMwVvCyKhjzeKyQf1OiBOGLTTD8/WgQk6U0Vlqz1JoFjhi
FnGmri7F/Lbup83wGPXSQMhdgm4xNHlLbufxbmfEJQoKT8ydZrpbkGQjpUV6vWjdrZ3U9jKYBTzT
Iwa5KwOmFxK/OG2odtSNa1C2ik6wPHtI6HUlM4ijfQDhsuQKWGLhQLJnk0+bQA6QzJBlk1rkeLjh
0UFxqCrlvWyB1AEs0vsvwW0KRSfcpO2lm160mQ8sML0QXq/1ZNrKRTLN+uHiO2ofZmya/1kkYrhy
lycg9IJ48TqZuVwhHZX23TNxkawTeimZv+rH53FG44DXGU+/gwQZO3EM+6ZlpxXp7qJY8Mk/oKPA
qb+GTqjbMDMMwaIbmZKfFNVz6P/Ir7/OBYhSELQ0SAp0lnmj7ek1PLPHAUG4+CdpQdN9DFe7LUBU
aY6bYBG5IiAsTS9xulCuzX1p7EI5ajQKAA7mpADaBQMGbzHSQ/M5537T+48OWP5ukWElBfkjforX
HGQpQc5CEnzpw3spDd6SDtobAvjeNn8mCo4HhdfDDLDzSC3wWGM3Im+bVsUMOXElAVSW2Ll0+eA3
8qwaIXQW4RalmdVX6s3ik93w2jIXS3F29bwzmJMFkptnTxFcZ0xYkBL99LWEqQ6ADB03GNugml8H
rIqVSgXFP6gAmcZhkcDvaCVtcPP2hn/tlRqmVFjZ+zENsqd2Hqtoyr8ZMKYvmfeZNGI7zpmOZz8g
45WfUAt0QAop+EukBJu4jaWMvm4432KADxUfPQBvfNbQjaTh9Gkyw1pSnqES1uUUxiuF12Jk3Ny4
/dFBmj3CveSNomz0yBLNfBip6eifqMdJIC3VgU29u0L3xx0NleHwILZ5vJDXh+diRZCgxolJhO3e
sJG5g7R+IZjOBx2ZzErhVJu3uIcgXM4coUDCzmD/QIxLhGDyz6/e8A3cWhkHrxftbntxDc5wUBgv
obOrzCuWoocjiMAeeHWcKr6bNNT5fY7tZL+VECidpxUD9EK6NhAnGMwd5sFwjvY0fqviu37oZjfM
l2qaqXRza8kJDdoNzSImHy8EJm1RSoH/w8B2joSeOVcXANW2VWhaXynsloT2xSq5DHCHt30nh1Nc
QZyq1gzDqXCBaLOROqxAo3rlbszbsQoglSr6R32+RKlnAUFAeHJRZNOZ9z2GP7owV/5chXZ3pu5i
FQchjzRx/JJniaeIb7tDay3ZcUvLUiD9gNzM1SkSMF98/lIOhyctG3MGm4x7XzuHfwq2fNf/v0r6
6DBkiQx+JapzzFpN6F4RQUtuKxoQsuPd2AxdwW9TY/jceD+4G83XpIJgHdnpFACBQrhFAIcLi1nm
aZAT5ssLT9H2hALvkvKP03lU2MjDc+YI2+Wx3NjneCl7gsnn5Fhais4Ejh/udB/Swbq/8w8AgIa8
OJTziwtpxU3vi92+iBc1z6gFqa7nt7cYWrLrcL4mmjOPZnuA4SMcgCT/DDXwxXXh4ovlXyQVAZrB
Du0qfFBqEKM/fKyp4aYM53TqJNfs45xaMAhKmDX5nrMbr/ONUwk17UCHxFaNmzYK/cqakKeL6o3U
/fzjPREUSWZR7oV5g43WUSFeOxbP2aeLOIZg/MKMjacQQBoOmen0k63cEVn9323aNzQtqxrwRrav
AuhBBtR6uqGUSNyhd6eaGRhaJMc7DhEPysExV0Pq3CK6nugZyPbenm6UUJPuZLBCgus/kovhSyYm
DR4Ar73pdu/hVr5zng866NQiuWv2Q2IUOUErv0oHtZ/VNNwU/SECqNgDDilzCuQ2Z1nz7AaRm6nH
1jz1T39OW1/P/lhfKEzQV6H1Mn3GxIRMZXaudwgSgBumcyT25wOJG8r25j9c7WloypIUSxCm0GcX
2Bhk3SGHwsxzgX/P8tDfVU4KRSjg1KJE1vBL+MHaCTdvdgaA0/kJeMmAeBxlJ2wnzruiF5L7C2cV
EkOAqCIV/Qs2LiyfDyqfJFuXgtBEgHQPzVKI5kbrXhIVVaUJnlgesZuMqy0bN2X+hmV9VNLtFLsY
kMkX+aVas8EfS5keicEEdOYYukctdZnusXJpYFnhKwLDjrlFQsgpLpkXGNHFe7t2C/OTkvQAuE+G
exhos07UWMNzhHlOZqlYYK79zQix8NxvGYj3jTsEzvu9NqZehKQ+alvKtR1yc6x1RuQKO/CNgNfq
R/XyImp6lqRmw2Q/KE8aQMOgv/z1HkPWNIS5MmxzLfvNDWJNg+2oNnP/JLbictTtxEYfZgqBrCCo
pI0gO0VAG9JQF7bCbhCQxKr1gECttndHa+85DmZGBuFvsL+Nka71F5i7QDCEZ1CDsSxSnOOGCP7q
fWCzDyGsXoV9P+aPZAThH8YlHTzMfo68548FBb4npFzV1TEpA9TKrMM7SeApTqUCbFmF+Gfv4eEK
1BABeSk8fyIuuml0bdm7G55B0SZhH88x7AVXrnVfgAOThjcy7Ux4UPOZLsOlLKnQ/KqMZgcKMu5/
k1n774PCjg/RKr3/WtQV2cCcLPTwclp5Y5ueTA/SDLFLBXP5FeCSjRYF8kNtIfdnYP+KDWu02UOt
pbBlML0EWqgAG5oEYwHbnNcEFcqzBxPdBkcZIj7Os2yF0sNqP//382OrPLePbYBdxrtzAUUN5FAr
lR7MC7Pc7wL0a41rpiT+9C31HPAQbNgQ2SPB4hndOoxZXj+bGsbFol0UAOgF2NtuKUb6Fz/MPnjh
xB1Tn/JCbK3VRRzd/HMf1y/PmwrvC4V64vRPluAvEf99vzTXhuzCuEKuBVhjQmzZyy7EXDSLNJCT
0SljsX2phF0tAFDnPRRy6YK/7eO5CAxxTx23pD2KHiv5ZYYoIJkPVEj5JNzLzT9Le0HmjjSlPUL0
E04dB0/rF/KN6hpIw75gxxrAMPj9Y/DcbTcwgYJZZB4Iw0Z9a+sYCPDPCh0chd7NrvhB65wZksMZ
njoiHI5fk6AOWw7GJWdkwyPtStVB5RvX9jszY/O6BP6vZ8brP+0nUDdKrklJqsqr3kSKUyb1xQ85
B146W/8Hds6TajwesNVJ1V1NjNM8L+xSBOsyKO7kvpfuvN/InVYLcpey6JUzh3uuDfY1Wl7Cqpi/
kheEV4s5Abblprq6f6hRSJucANQocplS4gTjL8/gt8xc1fJ2LHxoIp0Va+5HakSYYNiKKD2cP6ZN
JeOnZAvDsKoziaqEluW6MYslniXEaVfeqfAPQSjAJoAf8pij453hr3nkP+wlAMhkyfZLWVPRJ1Zb
e3ik/x0/+a60TaKH1gyv5dxCZRabW0tk+aJd9mkyP5UZr9GrgZAU7DaHwwu5c66U6ru1D/Zu0s4w
NIZRzMtuS2wfypV7CPxwzWaW09aNCiUhbkGRGBkQrWmZ4QcL7cw6Q/91mEJJDZCQaYVbwx+vO0m5
WWrIJsKbJ83SsiJDoBXw/6gPzCP9SdJRgQcK73d4gxV8L9UlbZVFYj39NVSPKKaggPPwXM6pbh0z
wRNvTQ5utRAaECM0TsRyGAdsx3087SC5Ytx5w9C42aDzUtj/MCVzlpY7YPNY/h+FgAuQLK97owe/
etNlDzAHcCBVq3ltY8lrM1EkFmZLiCSBHgVuyvkHneal8XXxQ1Ml4WWebNyc8lqpDtpEFRYk/S45
LfKko6zVzSIuKIQbj19cLIamGn4RV5c4q2Gj9vFwlxKi6k8/IF8xgnyOa/ZGe59QlwC6/rre7aih
NxxoQocEbAtI9hWIsQp8QzZTwIPaAwdixTFrkmS5eXI6XqyO8o89nd8G0+EoxIpLHXSwpwGAZMCs
BbZcpbj+inJPbYHsg/hJj4K1BcstXd23t4XU4pG8T2ZEIIMi/x6ll9WJwE0yd0h1OHBSzvsjEbna
XuXaFGBkkj7yW4Jozb2NBhSlVrDRHtlojXZ9TxEAoaEWQxSjLvW4iR4wWoOh+qQkWO1D2ro6QHeC
2Bn3CHyKPvui4s7YtWv06FW7+qdt+cOKqpIy+G1a50eQ+aX6JX7bCbgM/MWJeWsSeyvTYU7ffUJq
jcWPC/ivITsllogD0xJgKQ9OgHTtvGZXJYovopAfNCiiatuV3JRKU6D7wWkTI8UWNgqBVePe9Mof
Da7Yqet8URfT9VKMozqYr9EcCHLHkAJHLcmMc63tn7XNEV3IC+ksnEardXUzhNvTwBpUxgWnZMhu
6gzocjWsajTv9sGxr11tf/kraCjyvWHUB/zfEzS9dPTSEFSwi7AU2KHaXE5pXZ/g/VT8N9g/Ooen
AaYpziAoMLcE4/j7EpFeRDZXE5izYkiGy7SFzYmyA2EQS4/gUWdA/vYbJRXa0cPu28DSGW9OBa7s
9uvUqf5E9dLmTbveZfqD4CIr1ut/KDWun/5DDGGTbgiU2rFoPgLBqwksIG2XQh2sF5P/Bcr+1f4U
/FKXrMornRMY6mEvfr4RIJtiAKTnMHR7pU4uRktf1i6Ibt+md4G6fCZma0p3StNC71iqgWayNsze
xH9MNUtplGeyaeIkW9ImTUm0fNwK7LB4DmH+MDWWGc0gDikkse91avb3mW3195e4qd+heuECqAsL
OUNSR5PvxAL/aNkrNJsWYCy1S8aog7JzjLkMYuWC+5ui4SJnYXmjUJJ2n2nm2nQnHbx6WliziYdq
GQnHUdI4VeiC5GbC/jh/xuyvHE9Pcpgn4BjTPiYCTO/AfgUG3eG3XxpCLk5eExT5mcekIKx0x/NX
JpPfB7L4dWTqTqC1G30Pdal3kZFMKfjucpipiD0IZJ5ytxQIviDXuizHb2m8j1bpEM9gsrIWTJRQ
UsWbQU3N8KyJnOlYNNTfNQCKUvf17PvoZTUpRrQmg8U3jdg0qKctQ3P79O6DsAxpooGBJNXBIEJX
tWO9E2h1bEIsHxxOtWJwLw/pjXCkJDDLZZcxpKSTlb6ysPGO1RGvAiB2pkgnhJGtr2nj3FvskaFL
WmYFXhFS6IlZgOlXWXXMLoxRgPz7uPPO6sfrUgcwfSuIkmQpsOBv0iNB0vgfPPMmv5FZDcz77hBV
rroB8YtUiHTAUN722mwgZMMXmu/DHFCxDYHnhQoMycj/t6jmdD3rAqEzcMzqeYdoAqJkPLD7MraL
garAbCkLgib19lHAXhBUNa0nCLxbUH2QLTfBiXKtQYd0mV+wyR+GH3pHBNlVCOjWDGuVWjzsrQ5n
zHG0JvYRJe6BCXG5O86FfJHKTO13cyspwU1ka8i4jCIS20JCF0F2ruwoNOkAWZdEAo19kBK/1q2B
2rl7CqWBENkenfmjUUpJ/LoGI1H9vesfa8pc62thbGFj2aem6cUO4NkQVuKgedXArv9njeKlezIc
bPpU3LVa5QajL3oM1w9DJYyRYllzrmwpHd6VpFqonaVoI3tJB/cypyBasExsAaQKWzqLPGTvg3gQ
muWyy/8rWQsRTj5BD1s5T85QjVu27jJpSiJiqHOEj+NqeOv1N8JSwv0Jgr+LwceL1fxgqOrokbs0
0b8oGw528/svK5EYrNIHUQmttOti4/7Ct1e0fDqMnldPh+9XCA4Lm5DFPfrVyagkKtDrIFOTpuOp
lGeIR2rd+pSr9lSayXw5yGxe81d0vBkj/e/w/6YBNdcXc6Xi9+rJvtXXOLarrOP4P6BfsfKphWHa
OjvJnioxyMoX21BCWzB/pLmpbf5xeaSGGxvBiSIp0m+nBTK3Jy1Gv74RAzIqLEixaLVl47Hngr/2
WFHj4hmu5sBB4R1uhhyQAodoKZBwPiYsYz3yLR1YZw6m++ZWG/Q2ufvdpOVytKA8eliMZpLVvjDr
9+YEZJs/i/v99zCiX6YcrzrpwuKyUoj2U9bnBKdahJuCx3WYTPUJQ16F5eSQuzejSgjFIiD3DVZE
MSUkbj+MKQIRKwztPJvUT/XLk95m99e67JOtKdtdA6dYE2CAV9EEvJWOXZhf8gGlk/f4bmia0jYe
s/UMkb6+cYFGDsozJriOHJOvW/3AKyPySAFh4h7GhSbZyDXdun8kd1PxuZLXnSw4pL0EdPhZV2KA
efzTBsNP0wU7Gh7eaxEU04mnrEhvFAZDHzSALmqmuYIwwET2bSCe1i2qN4m/bHF47QSEPa1cC5j1
SSWjgSuW/dYRyyaFTiyl5KUjlYq7B76aGOfzS82PCKkYvs8NI6DDDI7laPdk8vPE2bHsEC8dbz8H
DArdHuTs6gLjupwjCpczxEjTO1pie7CoG6hVA3BWlFRJo6eZWhmHP/BNO0+a8DR/GcFEjxuMF+aT
s9Uag1Df4iKjHmVOYsDXKrAqXMmVXIyHJNE2FCUlZP68Jcu3LLQdqVIhKR/ijAA4lazMt9tNyYDo
MyMef5HnWWbRPjB9teQVfOMkHU00Xe8RSXuVnCme1mwNk3bzEq3E28PyXTWU/rvSMX1HyPts5Dqx
jjpu5s7zUUT9A+c0t802k+0x4TqFzT7yuzinko+9U49doYpdPbyIbz+YgunONsC6f614+ZiwHvgY
/rGU6q/ILSaxaqEyg/uwjRYbWoqYtOPCLWEuxYFIa+idt5s0IiUfNYGf5ODicbWFyBKghFbu4fKV
a/XYcL2tpSy4JxyM3WPZ44E0OjXNF5YEXGOB+lBboW5Q8jmrkBGmw1DTmGfhjdw315x6scEgr7j+
1incTObECtdaM6qHe1VXJRV3k36odk5o/ARrcZ/GtPTbREm0W7eNa9dTV9bDXJKkfP7meZpgbtzQ
E2fMp+1y3Yw1ndO5HTmtHz+SRghg0FXG7PRzNEzN2wNsqW6FjuPFSFhyi20GVlGdHh1oB8a8btrN
a1+J54HTyRCz4iEe4d5p2qujMylrd5fOtAnNKAE1wAplCcBtDgT6AdXVFjmEuIysQdlG1pUR8Gmw
Y2M5/l2kAwGQsY1D2dqwEh8LkuVFxVh5RQvBIs/1mDEvS99/QsbfTT1JgSxF6l8yO2sCdC/RkZau
gxsyz+dqlNr+scIUy3v65KBuPUBXHOBP/XPbIzBaOCkHFxBJDoEAP4ZRuuV4W90R8bJlWCyv8Uw8
heZ/hfes+01tQowKpXBf7zvu6Nz0D614glyuxCWI2jXUKbSOO42aUI7ybN5uIIfchG4IfKfIkVpy
LKsOjBaMfMzkBZHLJ8ijPu7Nd2vq4vSmcCKqd9A2EkbtLbaoWLjrAtBbOe5ZhXjYgVhiTcNgH9pB
kpSXWKPCUVup7FZnEQDr15hkfN6QeOjaOhV8I8vFV8IQKQdfcKX77FbTM6/5unTb81k/WOfJgtj9
dbr1iA39zPNjm2zJRfDW+dQOuzRRX903+YR5X2d86cSm8apmZnVWMKDcvAsLNMAPd91zoyFVZ7zY
MNKYrHzb467H/Y3BifPz03cWPCkT5MgbFzgRk7BAPj1LRh5Nr2N72JIUm9TWjr01P6SGLlXUwEuq
aUQK2QUWQKV5GEkWcM1RXafrUbf9lqaJZPKyMpLHs6SWyQw14rhsCkGN3myzx901zLj27lekMbrv
q7A3/p9M9aPvga6JAoPKyX8ZFolmh6jIo7gZUETkCxsmstfr0fNm9wXgM9SWylkpXOtdTrA173fG
iDXPIGi48PpQoY8klpXoF9DIhP4oBS9Yhl2Mo5N//D6H3uz80xf/CwiPI+Aol/WwfkxP6t5T+Mw+
1lXqA5QrTKIEs75tx5bz5bm4vyT2xa2ybxfwlluZnqwvTLN6RR6irDAK6l8rMZLqVluvYx00NyDN
TPM8tzyYEV7svXHFJK0evpSKZAcquaHers4/oODEssFxVrsw6MhLZb8Bt+xXL8JDQmwh2k84zRFl
t4G7RnUFwJyBInIFthJuey8FoYzOfET7aMdTjBSzUjZ2g7wnuIdZ/PB5XOEMWH914AmtKlhDJpVG
BFLgeUkuo2sdlSF0j2I7Cqa8q/QZ7uLiOAt6L2eXeXx1yg6I0mnrpr6g0q5PU2IjDV4RzLT7vSHt
GJANGT3/cokSNIESAA+0IMDa2RgdUzo3sTde6WGltBioUEXt1rLSu+C24PnhAAJqs8zLD4YzUX9I
GqEqlAZPesTErzrkUuCFmRtftUaT2KegIrPB58wndd7hbl/2vM5esZAVI9+i88gIw/rBl/JDCKH4
OLowYT5nwVqNyM4QUTVtqITV54oNuJtTEDQ8apPa+vYYFoupLPpGSXLgItYmk3BYjlozBfrkRxWn
NeGsU9u8jRLvknBovB3WNTqPiTcg5NlA0cxcTwgCBId8ZjqO4cq0tDxh3lkrdz+kBcpB4qeWn8MU
A/4C0hsxlLD1qb+ppqRmrWdozi9x6/nXr+G39gJQZxhxf+1bJdtAgs2Esvw1JqccocdBXm2cSrrD
czAUgjd99e2F6B/TV2ZW0RFZUz4uQQrGmLOT0lCRzGgcMG9SEkCqD1n1jRXfbd49k6gNDvK/bA9l
AvgeSdMyo1BJQQavZMEXy5ac6p+CNVSYuB7AiWWnh610FxLP01wqVfy0L1vBnT7Y9BnXwQaEbYL6
dqXtUCKJPE99oTE6FXLdCyP0TJPY565rA59jHSJhBNK7yuQ1MTvzCduloocVN9CNXsFtQ2Yxf7jw
Mv6f+FiDD/Wx/Su8w+RQXxxM5TiElk4+G4K3YQCQiepIBXVOlguI7bsg2/XdUwSUw+6ohcoF3DUo
Jk+UBL1XaEbHBbcw4m8TSwskiD2C9Uz5PJvjYmCteC8jd92Mgvu1Ea1KJdu59dUup1EczY8dan5s
TD/hCnMA1jzesKFJKT76a19xugdFeY9mvanyElU0GNDE3sK6uIU17/cEIkTH3sjzSkq0aJJeh5KO
z61nFd6X9EHgvCqX3aYwfOmEzz6kRDxhD6J/3Q4R6IVcQzxT+wHJ/JQbyid1WNP3vmC16bmOqWdt
ZQx1iWDDGAKoyx2AK0+z7lhnZb9VL2Slu4E5paDmEc/jsJwLuzLwLeIZiMOoJtI5zJj204HWIC25
QwfPs4UfM/hC9ay4yc/FziOePlmWCrtT+F+iqvYjqefJti5B64/MPpTdRfQzeSoco2zxhCz4EPKC
hx/ngK2mXKl0wX7jUQ4mHHNzusX5MsF0bgwjN/hcNF5q3BG2MuVhtHkq6QQVpnyv3EYz9KxjsD+Q
570VbDYsxN2AmGUdlslUyxNu11PabMD0rhyprxSfRnZmrMpoRfl9wribJR/60Jy94nh2l3smARR6
C/65gLDMzvAxvK2scIIO45Lzv5r0pLj7Yisfhfu0Y/UacmNRzHhWqUE+zRM9NO0xO9s9Wcef/tTt
Yq4ITGceUEjVHUblgON4ZPye1caTvZYjU5HzxmuI18LdfAsa7QLLgK3q4tXDIfbEsFRqtftG2ioS
hyBkUotCZHzaL+WeWZx/ChEM60fRsfxYsqwDxpDKmKsiUaCPhoKRDaYtIfRwuMKOwcYtF1oWeF0u
1jZ7JwEzlQGjSm8vQYHqSnqNl2qTybp43xWqE8kOLvjHv+FV7tx7X/OnPH/EkFYrO/5Oo2rASzyU
HItZEzu8urHSmiI60iJNAX8qRkcutgZnUra+K2k63CUWZm7ZdRH6YPFL9dt3sTC+/VEbO5NCvpSk
G+697f9eJw4Qmg0yNBpkv7QdtGBW5Ql6edIlkovJyBHd4tXRMUVKgt4tBf+SmHxd9qp3AMb1EB/j
tlveDPaCD9Xck4ajz0Nkyv8lbgzXAo7uyjza7tRH3aivCudo09Fehi30/mg4GNbwnMta9WWImMui
YQT65/4RX/SQ0bJtikwJdZFGa+Ua7+BEpUqnbtjfGv/xKV4RWztvm7lAcICFSjABqrp8gNPEto8u
nQLuF8g+C8L3RjUmFOZXYI3RCJByt6w4oh8kpf5KTrwjx8WTJ9pd7Z5VBlHfg5XWQIqZ0LChkvX6
MxvYqiUErkqX+x6q9HVbGuFsaVxFT4fIeGhlV88Lg4d57O33pWCCpp/CjAhb0broyafSz9kgWNAr
tN/b0mUHjJF09C7eQXDDQkLwcw0XC/VuO9Z1DSeOf4hDL13R8LkST2PYZkPUIaFKlgE3rtZlkWWW
Q6eUNIgX+joxnFC+Pb+mORfwH5wnRUuAJCy2QFd1T1gV/GTBjJnQwvxD6qDPnZ7FgkNOPhDVhcG4
iQ2Uv9zREE72J2KOYEp9Ze0l+yxTKoPkghs6v0IMSK6GaCYXjeL3Q9iqQa744nacmW2vpTL9DLhE
4F9DpEEz0n6J1IhHFZ670/chHKUP1kdZjx3Cci48PLscayPovNwtvdZ5cacYNucMnJQnYrPMwK6l
Ko+kmi+HUEX92N3ZVhrhQHG3cQ5ItPq8RYDDVs9PMAyWhSD8rxfAnHR0jqzUX9a7E1pL+eU0MdCE
oL3ZzUZe85PpnbBzr/brsc6wL3fde57n8HvkeJ0C5EcjRITdxWiCZRbjNKgXA8SVijUpr2/xfkbR
HYqfBiBJZXWVhAwFR4+cfy2+AncPZjv9pfliwC7fUaDLELjMHxH3CziAudMAs5VmAeR8wSpH7b2V
SH3FCfa+Fpm3mpkCeuLsTKGQ7fd2ukoYcHGzJfTUmKtlzZuC/AcrIdLU2lD8KfOJsvxg97+J8XP/
gNORhFX41LqBT6tBDy1JXoap+wz4N96BAyL2uxYz4hrzxZAEvbnvRx1W0hHpUce8wzJKk2QC3r6V
C2qzuK5Ng+vlh7wvki+OS+o7PcZ5SmMrePoWSpqyIUKICIf1CJ6mRNgyQUZ7rQ2U0OXLbKLjLJIi
fN6uSuVoPAjqCBB8ok+8p4+sbJ9TMJP9KufK1vBFLFNzyvO29lTc6R7DcSUNQZ3XecuI7PovGewR
kD7W/6Dj/VbIfuCme+fM65H+Ts1Z3v3UPFBtRP8yzjSKz25sVbA+ktuJSJhRZ+IGSuq9/Ce1h91u
5VyJE6Y4T8+7r+H2IVSkejGylLGNJe1z+rLNGL4IAh6snOgD04NB5nAMj7UREiHdWIhI+sPakNbk
NdP+hsl24qYeIXeeUW3147qweOBRgFFtUeErApj9FHen80EPKW4PR4PMPHfhpsDd16jFYXMccNU+
ZFu7GbFijGVXDHZIfGxvkUd2MZOyyyXZsy7Mo003FUeLmEHL5UZ3L25nG+1vW25iU3ZqBueSnknS
5ZixcTElDMG2m+KdjPvvsR9eWRR0ArHd4mlvySIGHQoryGPtVUqF/vvCZzxxG3E3ixauFh4Oc3Ne
PqfMHX/5fUOkL9sLCu02ZUoRMm96LgJv1lg1mdxwhviJ83sOht8dylyIUa4dPuAHTsgkWCOpj6RI
JIOlhMYPmI+2vfJoKLnX8shXuD3gA1uIQk44Kw8AQgNpBf4R76a1Fad3F4ciWPBxatbm4ShfNTPi
s+fya6IdP05scoBnTS8wjUr8tOmWvmkL5/Gq7X2zKiSwj5MJdbsx+JHqRps6THTrRILQGm1pTATW
wgbOg06GcMuoHrMPU8LszQytMzPUAPAFxzPiaKxZIoJUas5SBovUxhur4EwOEEJSuPg1amVNsWr2
W0lngASw8t/lDvOQQSFGLyQ9YW/TxkkmN07Nh0uDfzdF7VP4s+ENsByiimQIMnasmrHg2tlZJUSP
/UZQNRBdnxxJsNQdpFLd8rPvLBTX9ANyfqfWFu1IqdGVBCH9PLl+kwZzNA4IxYJ8KjpPXVGSawzN
E6t4hEymSaXIYynIXTXJ5aO5XH76A5SI8zg/bHgE+M037pOnm2UwavL67GA73vjbVJ4be5pJpqRL
foKMrKFQU1RbUmQ6GtDWT1KStfC1Q+w79VrRWvEKModMu7mQO7HGbLcD2n4u5Th2We0cuBz8KisF
YpCrDhA5O+zbX1FWwYlCoQjG2ijcpmqQUhZZkaslAQ+/7ishTU2ma0Kbd60LbwRIEcuSBBBcBYi3
BEgy9pmk7Tx5RMe0wZ11TuO+in+n2yu9ml1PEUASeOV8qpW3JQwdFGqE7ypQlu72zPI0Xp8F2cum
5JoJCjdtqNNEoLGd/ljm43YTnXcN56zj/t4dHaWH+0gTq20YfFUqiuLbNiDHwyGONDuXH6IBnuNT
GRw4njRMwoghJG9y4KfA5POSFTPZkSQJDxU66yO1ZaGhajSc47MuC41f0JantCdJrmH40MeH5Ms5
z1wveNuV+WYwSXiXQqpH5QbIyIi/wqP4msG/YW9dAaZfZWr2lOtXE/0uz8rM1tJ2GsoxcAeoLPPs
TDgWt+SCh9OKLmiOz7s/o1NXBVa2gPbDGwBaxWEzlL/IlIH5G5lgjhx0mdPrOAVFAujtQb5t439r
yPdTY4+Y7UR185bfIN8H/wIvlIDGTPAg0mn2DsTxh0OTJ191vygF3Bq91Aqqq/Kng8kkJ+6+6SRl
wVAgDO7ZGqapomw+iljb2iucACebqgx5v1Jrvg+e6sulsdqQY8cmuvlckI4B//tBUg9ShWnV2uSZ
9KUdh5zSrWOGwY9O27YSe0pP/fWDYaG65AM80P7dY4qHAMM+Je5Flq1JT1t2fwBKcC4bl2s5uKwP
JoVX96KobhzY7RhZtF2C1EHWCwE3s8h8RdeNWN7n1OOUninVX2ec/TkLQmQyUAIEHwDW4PQgaouu
6BcLwOxvm8EeFPg1esOeP1nVWY4jfeahUp7yM732ZtqjcBNcd+/rWHcn45IDck5/iXjr4ILc+NYM
jBNIDEKmnrWg+BExvIyK6h+gPFOT7Zm5ftAAmePhqmjC0R0AxUqHu17mMk+IxCol0ZdSNNzxFcU3
3JIhDGAAf+lW4SO6XfAtHwy6uSl3jWRM7GhtShPbG0CKa+1vJ1JEijorxWD49GfHuDrl32TLITJl
OVaXjIZqjYTvPC0s9+MtlzJ/TdftxfDpvaghiNuBjjE8elDakVbOtH/fwK0STCVLFhK9GXrxLJ3t
rvQvRRH2/f2rwuc779VGWN0J+7S3JNOiuD+Iz33B17EO8UKIi1nUYg5iiVMBRmSdoOjY/aDkIHvi
/pBOqn3r422oaHLgUiJtnjsIdLYUm8NTw49kl9BypMaxVkBSxhm6iKykvz6xRhXgMvPY73YagF58
jlTmesmoo9yCTUNqJbulnjnTYMIkE+tA+3Ioseaadn5hXs8UEIVUPQRRpb+cr06LPHm9himlr1uJ
376j52kjvG3VhEtU05KPPtm+snlrHSygCnCDV3VR7KJfu3w9K4yX3+tVWC3H2mqppdUVtsKdUmom
DyoFJj9OYhlXLi9/0CD3/z4dTttdyheXHIhl4CLnyPhgCJjzSNDuHKPkkYC4DQsUQqVACEl36Eq6
mKJsEldRKjpriYRcS5xR79uK7//XaL0J5X2JMU7kP+1emOB5W6NRhuOBXmqVmfATvUzf3d9/eCyV
GNYpIWnq4Dh702AAPP4ZaszTpliN6PxdALwZ6YyFfNgv/fUY1u5eS+d47RNo295RDvBcapKMngFr
6t+ClwVyima+fwdtvlc6OvQOYV+gPWL2jmx/wM6s8VES9Mpmmm+l4ZOlOczDWs3NgmmPJBtBWdXL
0ipU8cpGhD9tqpu26UnmYNsQXWCRteLNmRTq/mSWfIvE7Vt0iAOhR1BwulBmk7gSKUj6eupuz1tV
XZs871/3n9Cp73OKqGcF+3GNyN8ygP52RecH2+Zcqe64b5ZUiV+q6L6Hnk9xhif1AWhawvFhcVxY
pL8MGvM1Rr0h0vJ6CQkcUoA/RVmE0zHaR2L+Yvpul0oDww8DA+APqFo+FQLiiojerL4KTVQDhR9O
aq80Fshgn6l1DyoscGJB4aJMkYYuq34604DvzyjHlgLKNdHTCWvS+U7/CfOqJcaRUojJTk5W6wUb
qWuWWubz58LGLu8X7iEpcpDn7S4fgFDA6kiMSUTTu4RF8lFhA22tE4T4/fw6RlVrA1w7AuHGRkBR
JCcuag4Ww5nzEmdJJgq/sg/pCAQgLsGzajaxAO2RG7lpDK+3yl1Z1P+x5jvPTj53xu1935GaZSKj
jdQv60VARYbNGC6Np8OLMlgeTuVdFviUe+nMglMHrcCuacP1/JZOjukjz4q6lnDgd2OjNk/IBtKM
W+rmlMylRrg66GTToRXtW609Zgt5mXrTlF9Bnu1aQHWLLFQlWj49GWFjT18brDVZ9zULcew4HbIF
3miKrZ6yTJaJWKjRnWUOIy2eH8yGtHhro1U4LZh1XK9PG6VP9BjezkboiUTLa2opLSgxrz1EQamx
DhGedRaVAQVF55dLOWAmqdXpIoo6FVrvXCI7OLyvZ2QO7iLx/xsMdbmkseQJSMwpWw3C9Qo0kNz1
T37WZHnUnrfWlVHtZv8JsrCOgee49rwWQvWceS3ITnuePFWZyzpnFVlYHwq8k0K2EYpL3DeoMEzX
KQmS4IKuLmz7Ifn54Sm+ZWnxXURaBLEnd7hLl6YCkOWL4AfZvrN70twXyq5QceBCg/5nl+Iji/G4
FmEMr/XCcZudTdmeK2/RqUTPkpnB4BdvYk27ZouKqzOGM6RpmLeSB1rITi8J/vKFctdn87A4dygk
MaS5Ok0RahCgricWjbz/pGWO2hg0GzlrH+5c9VOOOwjFZ+3yGWlfp17ufG+TNv2fS0Zoezs7EQ1q
e/XC2i/xc+81F6w2BzUfey5iBeA/pa93jXiA1I497svs4f9ElMZPsMn8Ra+0Vyz60WxELuTKc672
UA6CsJ93ZeOxSXDGo/JRx6qzQkTXRd+9km4u3YD15oXNMzi8xdfi7wRnVQa4eqbDCZwqcbbU1eYT
2KKo0RMec9rK88A4WEOtfbHTFNfPHdLM/O7iSZmK4kOpR7HxeGZbuWnHudkXQerkLxDvsdJQ57kr
IUHRlQ7ARG02toLBW+qrcQ5gP/crjA7uasDv77cWudPJ1m2QnX5GQ4S1sOzpCo0FSHTaNTpM3ZNP
duUuI0SWEUOQyuilo+D89GXA4Gym66NxmUBg7PISvuSy/gYK6o5E9e1+6/odieMfKyqyRxhhqhvW
tMO6wHyiiLlbkFQS2/tsZkVBMTUKL2Vdgo0njEDn0ptD12KAotaw5eNbToIt/a4eL3a0mKPMjCWn
dHkQrFevPf+QfAWe4/MzTiDcx0JIWLf0NlcLPUsPjhH+X/r7B5J6RQ/KCkWIR2DHGBZoEahyVX7s
Zr2DdOhfqezY7V5A9n/KG/ws3P59uPXDHqi++Vep5vDQcLrzw4xI6QdjxuqBAF1HXeZE8ghmoWE4
z2U8h3wO0Wj5WvpsoP7dGX5SfDEx2WQ2QUpx6AIkU/XqBFY5vT08XyfAknu7H+FjpBtdVvcVdf0z
DILDWtb+P/1tZBYlCjUH0rithiHUQZ1IWtbxlav0E0T83oMTOVLPvnS4dAZY6B/2EkCbOorhskJ6
37V9rphGWTRbtbFQgSo1XilZkPEJgvRx7qtyHyUXOgUNKcuZhn17n7jZkxWq56ZFEa2f5GMj2cvI
kSGJMpyr2qAVKZSOb7OihhTwW1JEc4BijEhxwFlKy/KtcAn2fXwiX+OhSvwafGtu9i3zbQhRL1XY
BKtI+SoEsgEpQ0JE5yQJc3Iai0/PImT++WAM3Zwy56MeE+MfENEBokmfOywtO5mL13/ZBHhmoL7G
43XnjnpkCzWwp9DPStl+kkFDb6aazqYS/ZVR2b4P7iB7IugiKgc9yJj18pOIZi+V9X55kRqhsIkA
fR81bMAzURDQOBq7uFQqi8szUMckigRP4+tUKOeWYGmaHElLtk44Yq6onwBIAcZiDRhMB67bhE/m
FqlVDnve1add8TrO1uedI1Jz5h4DT1Bwew+eM9yc68nXrJyBvyZXGB1b2/9xXnGOzP028jSKlIAc
+xN6WbCU124Zd488vWNiY3LMzb4XgQV5fMljSn4CUKtbmOf9/hikw3JMyV3AYd2fijtMuEEDDjDQ
VeBiMrlgdpHuOUKUR7k7OTfRxQeY+Lhg3Hn5Ak2DbQEwsaf5nHer1fB3yzE03fd4fu7ZKAxmZW/m
EKrTTwpTC6F4EOi/NjSPT/20ehXh6yt2DipjYDaZhoUafkkRMlRL3iGSCHMFyR9H4Sfe0InHNxNk
fvR6WKAx/e4K3lyv+Fy3YfkGb5T1pGu+ltd+lZKt24wKu6IPVbP6OS4XSvE/Th8NvsLuBbbR1MG7
dLJOlK+S9UulCKtqUY6Z1anwyzC0RFy7S1mZ6CXuFXXKPdAxEtYFVuaD8wY2ABb6pBs3HOWl+3/O
YPT5Co9hMzILWOU2D/JdldPuKlUTtV2gHrUmSWUw9I64McsWGoqxG8u3QFnTDO3xoNRg7w/jETS9
YSnNL1/bD/WZXrvQvh7qAPeDf2FE/GjOMUOb+SavhTNiPf+zlPeaLc/j2ZUuVryyFpCQbz79Gj5Z
CFND1uHowyOwdOphNAURuuSBJoJkLnnUErDYHCRJDWrMiVawczL+VXswv5KceEZOMCWCMs+pIbUi
IAmImQXJ/nbjtF6+V2zYBu3ipNynQ9qFPNo+GjgeWe93MvvAmMTPBKKI3XDKgt5IZtU3fjW6RaFt
Sf4vS2b+Kd/GKEd+GnzPbZyDtAuC9xi0YtUZOUk/xYMdBTAdMh8g3vRjqfGP3+OJfcidLlTtTnOa
Z6hxgB/F9TbdJdx9vfYv8N/KlmDQWrHIIGjM20upJ3zMewVBRKmDRn66axgaI3MAfURilPAQW+7i
+DaRiSgD+/aBlwjgtVa0izv+RhbVNY394lvQyMLsUdCzdDHWpSowiiGRSTQqcciJEszLtwHNiMbu
0KtbWeWeoG5Yl2tU1+nMafzkaZbtMurRz1zun+LLy1Smu9O2cj+Y96sa7kMbrLJuBOVaUniyA1K8
WEhkpSqzT7awh5CP26i7KZEx3Mno0zeMpSNvIfGCDDYudQ6cUWNZffBkj9j/13bY//JKudfLsEpC
WiEhxPcubsZZiHs1AmUnFOlQRwfDvpPyKDLNo+QTz5sDO1jPb0a5HFvVH1n9z3iQ2S1ZYBAndced
fCCxjyGIUAt+S/VLgEiqiXNC/8fMugXMd43Z0Ek54NiuQq+60l0rBri134js4wenP+rkih7KrSQE
cKQiwlZu+RlNnyE2ZoWeKqMA9P1tEWQKCL2whSUJvEmr2AHT6GOOT1ShCRp6WfKjOmw6IqdUTWAj
jpDwzxBjFEfE0qcKzMTIjQSbk6J47OWSLnyrSz4KZhi/Zk4ii3nOTGj6qCXH85jSI3Cxsn7Cm+Az
2v5VuXmzxBAvUR8yPRv/w7CbJgIJ+/vukOQn6c0v8GT4CWSXRNGq0Levpo+6r/buDlWrdhF7IksM
9IVGns/WN0QTVeyB670SeIp8wXiDlnTxM9vZ7s9W/Bpn4flhPYLul0W7v08zqMnqXa9Q44qW+YrS
BmNRka5zcNhCvj03bHB9jQOdfrrY9MaTqJ9pDf6jNCv18PALuERg4UFyjHzour9GyntDYmrQMsm9
urhzWjBPprwVRG8/zddbdXx6rHAQXbt9ifoY1IcbTnj9MSZ8QxAnhxq3iLAK/b4DS68TWC3fAhn+
xP6ts5ryMCbQ5JEk6z3aNAOtbhkPFdgfGnBW9f0Ac7bdraQ7PcWPN7LrAWG2TkfO24bDswngkMkX
uoNldPqvtB6CFI5vHT7PMD4PVCBp9Sr0BEVi8ZUOw+67+cfvcN9+n/74AbSimMfmQ+WOEdeB8pyt
BODhlA3ZED6LHLllbbI/JARg7fyohmxNOVwzy9uoU2P9s6urvGAPREmyPBhn1zUjCOwK4hx8GEmf
qU13RCnC5MNwTNzYEzehIj9sIP3loOLIqQ8YQKO4nXK9YiIdF7l0k+uOEFGq4HmNFHc6grGtL2Me
SLFP2e5JdfYvwSFICs7bh4MiLpxAnWaGlbupDiv109rDAv7avP2rjPfW3y8XCf0kM+XoOOoQV206
A+VPuKvytfMvLyNHOs5veNllDIs3zc7G8hslU1EphLZVcX15luNqT84pWH/zUcThnlQPNe3THh/V
q+2JarLvnyCuTzKH3YAEMwrUEUOlQNiVFneab/v9O5vH8YopO6kB6F/GlgKpXwwckzDL1EeJjwxP
4QrgMUu9DQoYTSZtny0FpGtOgePImuo/+KW1jrGiJlVKqtcME1QUCF+VYrQT6R2v+ZDy9RyEuQbD
fNeJivzChPXw1TdyAskeffDyPl/Dab3VMtHDvQW3VJEtJqGvaFfqJZ+ZkzkQbbcQBAuOVLrNgoCR
Ms+Sk5FJGp8AWAM/zEQ3c5OVoCs9VGWMvlzS6YelrOuEpyck8oANI4E3Gxo6ADPPRYc3Dhkbh4FB
+Z0lhRv8I5L3D+lx1qzmfM16mfTrf22T8B4Mid0mR7Lszkpwzx0YZ8dn/tHjSc2KdqYQJQhH50CZ
e2LjRgMGS/K/QCkU74UV7mU4GNFzTvnehahmMGDNkBdW95ggwQH3U9sQvrJYzdvBQ8Ll4NoqIv9G
+aEYXkF9cLFWAxM55izboWrdj560GZB3/TeWjAOrxlJdjG0dH0l88gpqY8k894QFb5xf+yrawcmQ
aiYZ58jjpc8QhEu1MEK1v6Rooh8ZdFxymdKPHszyyCgRhpCHlOqhgggb9h/4p6tyUMytSKfCLjrG
SsVoVxzIvmAyNbnycMfGhe6xhMD3iiaXxEk6EFiLIYNfSu72x9tqg8xROFeI/yd3VNgPloyWMDdG
LqW4Uw4ozui2QHg+SvTM64AeI6MUXdlYSe9ob378N+Z6SdlI9DJe5NodKtTedwtAqnBAqu8EGQfv
PVDUEE2nzP573AliXWo1AslBrdbrGpUMEzeONTbOEChibgtpCrNogNsR1GOxK8Q+08F8uinC6T/y
BuX3cXgvR89BSI01LQD87gGCQ2HkpSKjRDXWu05+ITmgqfjVwaSSZqI4P/5DbkFurexzW+Q4t+md
71/YF3KFvCOjEq2aDjoQGE2ALWOe3vg9aLb3qZBMIW+mA4UnuXa9jI4l4kuJzAN4rnmQsXkVOATG
a5krrmpHJP56kP3I8Jbz5LwrKpkVNL9kpop5JKTuJ4SLxbitpDIEsWYe22FarktV4XyJCFhDPAO5
E3D1C3XPvcwyDMBLY3AP2xYLNpCmTjO6DX4jZ9q5tak8RMfyVfcevodTmXyCtXHq3ZwsYXWFn070
epJRbKkCFbBPYoRDGhrVEf0ifqotD7BZQ3ciJUMeFpmvKJUpO/4N41QC4KBid6GsMTkqx6M+p+6y
AZpKBHgaqGxoWZaT7qhxyc6T9yjgxG5ejclR/G0Cnq3R73Ya1BWnL3FTrjHq5GUZOqpXRJu8fXqj
MXZFsgDgQALTuT0ie05OalD8fQswrjrHzxfqVoFxXEkox6PfW/zdfePHjs1+ym6AQJZJDFHG8xXc
3V4m7nDvoZUi5OOxE83vGdt0eGmDx9QGjSxYGKUSLFBIYIwDdLmhiwqJilvCrPgmLohgSK+M5zTj
PFwGMVrJunvCOkh9Mtrff6LKsM25Cq3Lw8x6t5LiP3EDJfR05aU/isg/DGDUFMtSQtf5jai2FYl8
+x/UTTnOmWcl+7H2g/7ckTIaYked0fcXVBBHr3JtxcltKDJZNO+Vo+Ne4OczeQkCv1KmBeGWEb5R
E0mFwEcy/hubKA1q6kkIvWNqNbixDrBFjHV5x7ixdLLy2q93gpJ3in2SoXTZVDpXJDUelN57KXnV
p1Ahq9WQrqblkO9H1pQqsJQn4fqFG0OSU2/AXT4biBzu+zUociwlo90r77hpkfSXSBD88Y6bYrly
DcLUqtjswSDSmy35XKgMYgheNzBkQVyBXdtAfA/pdhuu80evrMai12mMW3uYURyQlSTw/6Ftq72u
0Md+a9Wa5Ed+fwVZBGADyqPw7hLXKKnsOxBSqo418+alXPR0oE2ttbVw5ySkYIPEwyJ17eVa9cif
CzYtLTxUsMSPXI+EyIZA8PPJyAWt104RSWolAZZx4adrc9CUZ42NBMOHMJBHBauyZU4B4r7RQAV7
ya/mqdrXhWOyq2J72ug19gTkSK+s4KLgTPASuWvC1meB3SrCYTtDqVaGVI+HuQ9KBbLmEwjZ/UX6
/Xp3pMRX2UaUE4mRvNRsHVcOZfL5sjFAajsrDItiX+19k7o7rRgAD76gJ583S8gixQpprfaiJ0Wz
08mcsFoLdJPlNMTEfS+CbkBy4c0bStWooi8v/eJE8VMvtlqDTzRlCb6nb0i33L3gNLg7lAcJFbUG
WqCmgeTaHyx567/j9Hzxa7yRCe3sOEgOH14bcYzzpGrHBF6pNou8rbJ3oQ8tE+G5ShtPxHqhQIvD
cJpqUwXL5itz7vYe++64JUDq0jip7lol3wo4fzCpsFa4QSd7n0cTbsdyJcITWCf087OuYl1NYWsT
xAQFgEnQk4bMuiLeMNffh4QakOOonVe4tnh162BlVB/0GHtZJPsM7PtulL+cMDne8+qA+6yEGvp1
i7FeZLpYmBSqJGE0l7uYGefwJmYxFM8q1FkmiCp6zaGRwb+nkkSIwFcxzZfxGU/qm2F0XfFXzV4V
VKgJAzZejOPc5UUvHb9RTIXL9UOHgbERLmDL8/F8MD7bgTrPlHKzrUlqGZtHaGDzyLN5VBlCLcrU
p32aDAPOlBBwuT6NYWNqaDIGgeauQLa6SHGPMPAqIgqaBg63Q2jrbxPRJV5tW8w0OK1DtPbUxcMO
SX3XrIWlc8JpPUlGPTDdH8tf6J562WH1xh8FkJaDhp1zcEGrqxDRX1BdWaDu0PqH44h0Bl2zaIqi
R8cPrWAjff9Yv9mmGIACNa3WwvP7EYdjTWuNmPuW58duZvnQoKM+pJmDU8rpK4OwiabTH1t/VLOC
+00CCbc/x7fdPNpjpwCe+/k5ekvKrvwvJTR1ZuPxMK7G3ZusvmHXIWHNG4Otjrt0iZXLljee4zfZ
SCczOOJQW0KDp4d0At/iF2Sys/t5MKgi5+JymcxxAOcc7CJ/QZAr7ehHEn4ToNVuCdx5crjm00x0
NaFmxQvX5y5Y/mjK7U32K4WyfLJ6Hgbty+G3gz39fqyL8UYyx85eEi7WNmbfRGNuSs25tPJ8W1yY
tqvLckPYdoFxDVI3b+weNSG4KqNj3duA45lnHu4l5cjlQzrnEAos6LQSy3OQsgfczj63L7JZucX5
3yTvDwLg6sk2fVz2XIqAxHoMIVcOw2BwwuKJL3p7BiKWC1XMNcw4y01wgUmYjX7MjAZm6GgsSVU+
+UO+T463+qblv8Cc6xp4HC8G4jy3brGX2PHISSun/Uf68VsXcKFrNTN+f0WK+Tzdt2+wN6d9zmcH
vgoJ5hFjSTg610MrbPd4KNuKpPkccmolYaH8ch2uAtyk6HIOldje6suVTNHuupoj1FRTNRjlhtZw
JNNwWFbrlJuc1aEg0aZHasd6fv7WYxEVJVKDo/BvwQSvrwl1z4UnGB91dIN80Z4gvTEFuFCBp6BX
gugOxk25l0TtPFKmMRwWk0Bu15AodxsWeEtCA6jjtGVS2dqwh4A/gUXXgVmT891tqGwl9CWEFzzY
ZC0JHPbdWo4s4tiSLFus6tnpu43KyGfwtogQ4jdffK5WjVl/4QMyaHY46NzqRAIE4sTKc/Kcc65s
sQ4BtCdpxoDGwZWHJ/nccF8yxNGeyqwQol309XVrJ8T9nsl0aAwk7MsBgN0n0V5z80iqTBv0CA6x
AjCFDsu0rwYZ3efYMMcpEm0wQ0eT1tusd7bJPnNN3rbJEDnmbmRcQfqaAWQcj+kUFkalsp+/a4dm
T+Z4pyop917g+1dUKW8GV6PGHKTXgfX7jX8g5lLpAL0Vo4W+qjk8jjDOi2WgSk1yUKuNJsihxV66
u5U3j76tsdT+7s4k5mbNocW+IKQ5NmXS+wv2q6KX8QRnEbYVyIoZssJrh5o+z4VmxorvTnJyoTPz
o60TjY8hLGMkzHRMVs0e2PWT2bxe1/VmI5S2gZG7bPGcKvJv6UBkyHmjBC7T2TrMs9L343meOyDi
ihgKzw39f8YBKYDZxeELs9HKCbvaQx+IPaJvInbZudrCvTqirPCu/gt8dEZi/91VjdM77EWmA0PB
bgXG/pddJWdmztAXcxf9LbqvRK3zIpTD4/XzFUnthkxg+pxlPazktOIqvMzvoyoimzN5I1QBt57J
hElXb/VJjniojNIEpHxnXt80bm09XepvxluR0wnof2p5JjD2Oj1owXqOEaSGsbSl3luyRA9qPGZP
4h0o8+t14BPxj+na0lj1AoDmGxCFKAZkSNnAMDhogMw7rIT0IHnGFTR7b28OYGjVIgsuC35VAKjg
1xHxQTe0PZIsClHfGFw6/3Jb7lVjeK8uje9rB1FLFsOPteY8TNL414qsufWSczIsfLst4PMJkUUj
/vDaleBQKjsDMyBtxmc7BIJI+e9x9eY/jv9Sezk3gcngMa/rbllH0KwsMbdxj6dVV6iw71SyQptp
Rxqbnw/0lntfrq8F4n32h6ATrUP+WyYemrrfujBNPuPHotfS6l8E2N7OX0ubnSJ4b5yd5J5ROYQf
RVYBKwrleGze1yOV6kYv9H3ya7azNNrSQqws68g0sP1pZZlY5s9WJnthDP+wvQNSO3/SMBigIqv1
MXy7LqH/ggM+7AfESmQX/5lUgNwNlzTVhRurzQAa7Stzvc43Lq1Y2aGX6Mh/icTUdhxpD5Gdtv6E
+fUYu32ui8cvwV+0tHYOx4WcQyOJciOHWizwWG1mEpLeWZKYOm6TF3Msy8Mw/dDFffxegue29DWy
1vTZhta48rSN9UcCwEucFAdOwvK7U+ZV5ekhmHbnHoseeMBchnEf3u41OMyCdzMgppkIqlZPSwo+
Wi+rgIU2wRYphAz5FCYWPH5lZDihcdcFI0HfxE0LyukkxlyE7FaokkbG4cKQxuDHiEWQTR1BwMNN
PvF7pOnYCCWyiO11s9emQEGsD7ODGWXI0t0cALWb4wxORYqpvmXIHV2iKEY0P625j1fGUssk0hwa
ML5A9ROcBXcWi4SznYq1dKv5ypXqY3AWUUKlfjCpiVRUR5YRgR5FNDnNKoSGRvIZf8SPf4IRHTF0
r/FFJPLEZASc1wCsGvbbNwUH5yEWm4UFsDvZ8BihBVsOeC5kuUuK+S+KFJDz+rRIPhnjmMF3g73g
j35NUM+CZF1NFUE561xltA/xGc+0d2j2A18yKiZS4hnaWSu6e7pkdsAPVqCaqlKCf++mqo5MBaoH
Ld0or9l6XZhhyrrD2CWKKUpHnvMfZAq36t3sxWMNKdjgwtqCGpmoSwtFqs4NrF8dK/PLfeqxqybP
bWoaiM3XskitrQTWWZPB2YsAul9XBiwkodxC2Og13T481lu6f41VcUHmPUzJsACXK1YwYNPz1mYm
jugOCIbzWp9oqN2fPeYPLilEif4ChmrcVUmkOhbu/UIhB7j6cl4hzStpXEBECdy89t17B8yC8eoo
hgMOHA7eZTFsIN2PKNd0LDEonF9lkEnoqZnqLXmTw+Ijuki4m+tTBneHEMrY3GKfae8Tml9ZKIWW
RZEnNnHdhktiIScrByJbr6yV/Dsoue8j9cpqdBDjb+PkZ/FVs2yDoGjHGWZDc4A4BWRoQpELe79e
5pWzuEci9jaGERxdCWsT2h4BwYRrpch1Csl/8o5oeC8yVo9FY3ZLH+HVEPgPM0xhlWv5YhTjAtb+
c9dsQygVyNUe+HsE6jLUfoD/GAasijKqnE3Aq9eVvVtuWVL/31NjCBuNGJmfFGIWyrDtXLbNEr6a
RM9YlfEVUJxoD+Iq4lLyFydcdFkWInKxF81omFL3GtzzyhXsWjBedoN6nsvmXbk0vUQ4LGtxpGnA
DtWT/JABLWx5PICNCV9oXcb+f7jSdctMAFiRKV+eXG84ewwsSIy4WioB3x2jyo2sqsAcNOhe5yuf
xUsmuv6btnwldUbQ99uyzf/Qmu7xyQUfWBozDmNxQR2Gr/SHmphR6nQvRsbigVoEYsElUx6F537I
a6p254Q04XrOpb7hD+IzAj+LwMm7v86x3byynTVpUPI4ZcOzJYvannC4qysLXKb4NuRsRgIYP4Nf
uNMPzzsQy9rebS6FdY/Qs+pIbzkG08iSSp29U6KHLiQmWTrwIVjXo97uHnLdsaNgNiVyJW8YfcKv
U76TDLik0e0v9+TsNl+6j7rA7+fDZxhzhZeyg8poc/J+hBN7qv9vpSFI9o/OCrOFar6XCIN46n6g
iwRMyFMRK3ziM4QCvmlS6A+apk2qb9B3DtcAy+pKnMHd7veXFA2CvXH9c0quvaIDT+UQbOpOXaJn
c9RxQyuV+G4VPxkmAVXhE7QCqi/RumAVfJTKpRBKNgUXjtFgP706JYubqH72MbFI895UuTeUw5FV
ZoqTvrXREtoOUkWU4RCDBUz88YKSCkJ9PZsOHYIMqNXrlFeYxqk2892nKo7IcMrhgnEghUPi+0y5
Gucv9Yfxucm5/meRZMg3X/1msBJUCFGSMcSt347glqJJVKvLBt8B19/FbRgAry8lHUxG64whPWbn
gVtd+MdN5m/nYFG48Zbj0ojZmffZGMV/6wqzIujM1i2IfI3l7etJ2lVi4JnDatyLhl6HwwDpemOO
SX52njILHCdqxs8YhbuBbYTD5wztJkpo7PwmwhThfcH3+TvC4gi1hLMUkbJQXD4mx/N0LuNszIg5
Dy3fF6AKyfarDZzurw4rm+ZUNEQNI9mM7DDU1sauK1M+8ip/zcqTWD1cLR2tNwRhK3QBode5afH9
6i77VGdqMnwTsKWNgi527r8TWWcXkAIheoTLk5eID1SozXso2JNpoG/DPiTGM8U+PaYeBRm7T1Gq
snlnqZJeIEFNU8UGKiswA1yZ9nPcB3GbejFvlQzKxIZwQQcGKWLqNjpf/uYTNLmkRCUNOMjub0PA
4aaGtlHIbMn0VTl8zM9G/q76IlFXuh2yR/aKHLwrJpleRl9sqMQCV0xc4IvPMNO/MlTgfz366cFL
bwkUBqtxFNrVt7gduH5ilGm4exoG+E3G7vXYuEXzkHfYfVTrbsiD+Bav674eWSfXiw6LWOlE5BOs
kVFgLIYZOVtvfcMUCgCcOXfOKy/VQKK37WeZpWdlXbmkTD+zrx7uuT93X23ISUFTQMAO9/8apL2A
ZNWL5RLYYg9PnrzkEQke8U5IRmIJEbqJpmWicHukO7TeTwjac2vzsQq5xipLZP3Wei0jo/RWC2Ay
QEJM/rcRXW/qT+PF78WMtbUlkW18BIGR9Wql3JeQB2DAv34XHDu/T2vu7FJ6y6+EskQvnIXtL1ha
VLJEjJgY0Jd/2wnsEN1SzQytWtoVwivhXQ30tp69F/6ynsrSG1Mw37cYZMBkOnLVSfJlAUnLCH3e
ebsquZFjY4ck7/a5kW9G0nSBy9jSOE/Va8m1If4A3wftjRIZFVnNbVZtW2EIgptSMUoEO+yNW2vo
OqpYmUB+7+cE0Fr6QRE+qtnFcIdCPQQGAog7QpHr35PrXdbcMm5rMo7Mao3PLfyN2DYFz9EexWU6
/UHQdyGlBUrx+dbHNXAUpHLdFLj8SKTdonzA5PTESHTDT8X6XOhMuPS7KhEGuFo6pURBmSBqao18
7PrjvK2zMNVr6uyHj2Zd8oq8rAvPxJhW4Bq2c7n9row8zooS7jQEKJQ8Wq2ad4wUupxXtggdVcRa
7R1L+iBWKb2ohhLIli1I+anjySn746faeHwuDDyVfj3y+DryvYOjX1Ev4jcXfkMqAFmEG5gyeq2F
QnSIXrlzFD0US3MLSdVxkrxvdvhwQ/NlXSlEGNXG3VCbC/KuXWYa3IT5DXIKJdN7wgBVtpe5Ibaj
KoJ+twolLZHNQ3wl0it7LPF6xtgudRBzsXLovUWXnJV/QSUqkKu5rxX3MEvIr4VgEL3YH2JNqanQ
GuRCCPPCHuCPDT9FRzP3kaSNTZpC3TaoM0EU0mOfciXimJph898VWIBVDbXAmu4iWvZjhRQ/o5vP
/lHboqnvCq9a0c/YMbetLvSTXbPVYmR22lNFnbBreXidt9JfBWZsPLyFmPj3MF6bwrroucSkrUZw
+UMzPIgYUAZ5idqjExZJebUHhOODIdmTppqyfydqGnsvMSmreKVAi1bdrRu2tG6h7CFui0wukaey
Q/cGJvT4SdNGaAbOXT7rzH7gGzd+F8U3fxcc2xrgP9WDPUBEtpj2Og7iNtF8be6Rxsd00ygNL9oO
ycuuMY9u7k8Fqymi50VpeJb6IkESm74OwvsmL88Le3Z4Kx+l6WzUJGWBg/NMsNO2dVjWmwxrwniZ
cgKXNOn0g8jT3PpIs9yTjh2ZM5vc97Y8wZgY7WyqlXzeakR81SgF63koAk3sz5Amwcl0SLlTpWSD
vjX7yql90MqNXHZzCNTWS7xSuhNf7Zrj/fmi/UN/W4vPD3ukGAXlBYoPM/AvBHrAHW0RraxDeJnx
hLAHfvWwjc2gvZ2gFZEn2egn9KUGZlywNabdqyNhc3frAA1yDN9tfVIlq9KiUQdFtoBf5GmmZIR3
FkTtolt+oxo/GUepRs7BN68nfFfx/t73ALTBlWC8Kf2mVKOZPHWkEaFkK6LFiEbVcDuqAQmXviNb
4sGq/aG6ErOG2xZ4rQz+UTSTnlWnsAth9/QFQgklMzAFPOJ0ZwTLUBMmJSMqHmjXh2WD6k7khbRa
UyWV69xOjgoccTaeE+GeOHLKlA524INUXTt5FPyzVq8Evm0ZyDH6uz8Cb5cavUbCaN29Hc5tYJvN
9+dZ88n+Q6d3nIy5oE8ZiufiXOrWPguUT3GQuksIaptLRu1fZ2GqSJBMNd011QgmAvJ9rgDnnJIr
XXYZmSGGrDgjPL4o/SZcM+nLgQXKyeaHUALZncXbNGMbjpHE6slYKkYrSShwwE1sW25WD2G48SrM
Fs40DjieQkVB8+SIMvDh62PNlY23563xTt9zqMnRtx08WkbFVusoPwIF59oQzmN5XrfL/hoBMXVp
jU9Xn0YUY1RNNShWNsKxYnR7veKKvwBd9mcNh5dL2Uv5O7kik04SGNYi7XdE87pfMrgEwqw/tACk
wENWRUNUR6sxhJdOkYtUaahxQN1EJmxsAoLtmWrh81N/n8ARLVe+nG443rnn4GSLiZmK45yjkfuf
E+U3Qeqy7tIMrhAHD9vb0nOXpFzOuY/PXf7h+9T32n+Uu2OaPmyEHcc5OLNYWYCdR87GxkMosjDO
rdvf7CB7s4oNpcdKj3IP1FO3C/71//nTb4UhvUHxvWCVInM0rViwwZLPvSyNeSMGKJFoX6QR/Z3P
x8ej5PemznsGpbKmAbQ5Z55cf1mU915Ak9WhCi+pb8ZmROvaSGXj/fABuovZJTr1yDuUKJqNIGUa
GUt3gtvFANT9GCs4gC0vF5ArDCrmGK8cDOw1RBv3xcriDsnegBB2NfklXlsQrDtD9jnszUGoMQ2f
Fziav28AfZS2kgZaA1GARYXuDX+7Yj75sZx79TjUJ18LoUrtBTI+AONPrtGX+z6dDxuQ+zYiTK8/
/1bcFO+TmQC8mqx7RzZHIEMFpccn9/PBo8FA24vHpQIcSwRGdVbnM66n8TGSdDxmKUBk3DDxqcaE
+PC2OIpHPKiQ4hn6apRVWy+yyGkqpYl5BZuFT0auGVfwQFic0gkDhUG9Fqz4l6d4cISISpobBWTU
5iRdOYngpsFjkNPWD2UocWq6D3sHqBZUm4E5YU28FSc+qPWYS4OCJGcwM9UlmpYTaoTGO28gxwwT
0OAx/yRf1SXNOOy5Q6PI9NNYO9bT15/WBsM+UYrmX3gzTJuQgBJhvPQ95OJI6saG4NAXns9/Gwa8
DSpO4kv4eRI/08e6bVgJ0Hu+vAN2F+QuEc3G6ExDmfTKdljHmA91Qrwu/tAmJSn0+5wa9X94Joze
Gsi54TYF1GmFjHQspR8Dd/YKElmPyZPbyozXhk4ztCp4yilMuszqcSRjm7Mb9e3KSh5NAYOjRLyw
Ox07STIx53Gwlhw6LP1/bf9TjguwI4iQ/fxQF61cPGfvYav9ObxdACd2tv6o7/oT1i53RDS9/iji
1TsW4MiDkjPcl5Z7qksVNKU0i4oDLypEj2EaBi9uuy8P7atv9b/OTaarNUFfGhHaKzgBBJJggklW
wqdVwIsS1YtUDFAPVDIIYFUWADwVp94QdW9T4N5YJrr2Q+A0PxvBTWJZju1kls4HXIxYw0wg2OoQ
iXN20HF3XRDJH07Ibs4+PDpp5UJwh/nOQ2WRhh/pK/6HDxfhjraP9mtn2m4C/q81s/hX7X9WO8PF
OIPPMtNd3vTDotxzkkHl3/s+QlRlybaWFiKXZeOvMZsriBzOLaFn6Gu8f50X3+XjlMlinxDsCPxf
EOT/jhFzN2qM5u4wCgUKeOijEEDeJUVZtErnroAnfXhdN3JgRrznBTRigd3PbxLOPtleFpJ4fbIu
oPslso83H1YFOaSoQm8kAXBePnBjb4qVPokELWDbJgiWa5ZNVfCT4M7vuPJDwdy3pkPNw6sAnCwb
H2Jntn5qn0g3lDpUqkAJ/Gf8HLV2f9K0Rj6uaE0EE4gEH3VxmTNfqAzguCGf+FE80aiijwwp0tsS
ie0iBtUdfbCrc14f1cW0OdAQrEV6hHh21/UMuloNJxEqxLdGp9OMX/uYHCpBgI0wqZ42aFkqnmLi
kzyp5TiiKaQUh3zRZCCbD2vEkvGSogtkzgOOC9ae2D8OlNXcPYqH1cbdKsECxIvDxAJCeEctsK6V
SRz4E4oIzTxpgttSQ2+lfTlqthVCWC73n1wySdn+24MIZGbJvVatGfpyN3TgUWG2MtSKhcy3SAk5
HSwe0NMTUgb8bvNRfBs2YNPJeIN9P1fagTu4OjLuCxYH4+t6Qe251r1Bk+PCTg/Gr0Z/9MqbbRrC
k3KDMsYU3x69/AOJnGYiYaZkoATAvw7aaaxFEoof9PC5bu350hTJqUp365hH9DT/8D1JFr1kQZNy
+UdKk/vkeJRUhznS9FMSfyMywct0E0AUSMBDstsKcCpufqvRuzOXjp6kvg3EaFbtiq1QZGBqvNRr
U6AiXtgg7ggPWxXi7PjeaZEulaWSjtp6M++dyY/esvZYvzCL9r5nsaaqCVxdPpqtZSm5VOFUtXlW
+Nu9LyNcwlAJhXpC8wQ5bDCygvVryNHjzWWAsbse5Mcyof0OJp19d7wKXDsv3KyL4O0/beDtvo/e
czLN/kW/u8/bGM7WDWBGNx/tqmVeiCBeh/7bgfXhC3wfjoJD9GS30hDKICmrhmI6WYG/40ka6CXQ
CDJsprMOUps8s60RnmUgP9a/BQWoK/EoLdxKFLqkCurlYRZ48DpZeU4ft+KzmUSEUn4eZ7/41E/0
SI/322K77fEj4kR05QjMKCIwyd52/h7cF0Y8Np5G22zNwnI2tw8vngquJNHu5LLp9TvjoxiMoKOc
j/tq4I3tTt5XUOKuu4Bhduy+8t5vIGZKIhlt4HJO3ctXwqp7PTHATDWEPuEaFLTFrAJdtKb9KNnI
qDhUZjKTIc/Wdzd2cJ2YW+OXDtj2p/eXSarWfp8NE+k9SQ3E1Ukgc7zylskATJAd/M7NuEqmMBO4
aHFxFGw6SGWgAZAlnSGc8VMek/mzvcyOZ0zSYhkgjMRnmu1qcMSRNgBDs/7dKCLHv4GEBrpBborc
3XtgvIdjqX1ZcJKYXdJL7XVm3yRR75qiOmKP3pqWQ37WCfPnpIDmdTVtUBfK6O43DNVvn99hsSl4
bWgLV/IMKyCrdpVQOt3RFLhipctym96rzjTwuEFa4lWyUVszl2AVpxWPDpmdvDnXnSsVjifYr4pf
V4Bf4H2gMLUlosqZhSPV8AeZPD+1X6MWwlVj/nRJ9psm+17qi4eg4mo+nwMcHpNk2ev27jQ8xSBm
Sh2ZReeqeg9pyLkdxTSgREoG1MChRqYS+SdWveQiE2CdiUXmS1Nt+NO/M1TPNl0MYynbrUsD45Sg
gvGjSnll5dC6ly2hvzowUU4YsQMrZphLJOJ5qbarH9tpcnGCtQ+nHjka3oJSXgkPX4SoU29pVRyC
avm5RqsO79HqYjncaWs+BENbs7K8A07uS/r6JgNManfF15yl8KN7WAmsUB2og4jnvwVev6yKqwD6
GjvKaBkuGYFN1Mppyo/dOjUK8dCpRk/Mm3J8y1e+82RCwrfe2stYC6RWqW+yZKWNltGwj2XzXUmF
l9vB4xkZr90NKcWhny8D3bil+lzx2+/BjSLcAXy9zZ8BG6kzeyoVa/R5lma973aAkNyYqY7TCYDH
xLetCWR5pryGKPatqrbV+aHUFIlkSR8Nxr9TI1rDr7x3nZgxxYmvdMAb721M8oghUVXnWXNHwzoC
9sg2aJfpZnYuUceojo/luxo1fGnjS2zwm+hK9ITex/olVBCxcfi/K4XD+W55DtZkZ8EHAgeUqY82
Zgucgx6LRltYawCM/zn7QgyeVL74qGAEqfYBbspeT2M6DQsJ73j1se+1oUse8FakWrgEprw58Jrl
llhrXD/W3PDY3cYC+tb0BM3E+eVn90xnivQvMEwYkVhQTV9rFyjJ4oB1S14i9l4czk4p5kqUQPIm
jA/VJb8mzA13AJflM/bEi5Tq3EZmrcUBrCTK6j0V3azT+iobss+WuawU6sMbXcDuBG8mdTOgIEpo
Cit9xI1p72p3I1LAdtT5nXkcQ63ZGY6YEzkWRDQu+d+3YKIDHcIdKU9lZv8CC5Wdru5v7WYXY2vK
KhAApeIez4w/Ywn1B40iWE3p7S1JJSbKANs/V66/rrq+oXrpB8POQiYfVlfPXQZwM4izyiKfpVto
bL8YDUYTj7GRsq7IkF959OmDOpoILw31xPscP9vik9xd6UQ8VdlKeSxWKU3YhMuRKxOBwOKgDNcP
y18y0jR8eJ+3H2ei1zqlcBUbVXckkWpqWe0cxHGlCJseyyoW0XfQvuz0vbNAJBe7shWB3G2BfVE1
a/eGzSr/FX7MEDmtqJg8tDWjSn17Auv4aidMbg12vCOKUIJjahZhE2toQMyFV2n0yiJKSStU5Yr1
YN49mGCvvmNjywlRDbV6Y6lPzizFU0JQ2wo/58N0uAEtFJ9+NCAxNC7rW8kFi0xk7nQzltUovIvj
ZniH0B4IpPD4eeJiHL4ndqeIZoztTuZjPgkKofWkUd06E/bNvWl+SLMWF6ZfAh9dBh5hPLtymd+i
ZTbDl2VgclxN9Yww5TsKk9Jm2AvKJveMysP+3RhCX0vCVzmR0/1Ma3c+YXG9Ys91Z5emhun5Ruv4
MIVAXaFHWLjsAZxqfDbW7P1vIHZucmxlJVb6pALNAAEsRdDl7U8LyWIjkAz+CKymFH9iU1MJE4Wx
iCTzVuobobm7M6jNIhuJQBF1rUp5rVHv2Ixs4hh4nKNyG1oqXF0wk6s9AFLjLXDzh2V5TWRhYOpy
qnfJVchSS08Xvrhr87Trb2oldUaIBYx58twqcgmXOsBk4orht2vcJFF6n0AulPrPvJu1I0/X3A12
4bUJfDqwzdvU23iaebXxiRm8ClDe2aVzoYr3JHENUG6/8YbmCTjT1JgNXGUWpMCu4uKo2dtk/HWf
jZvjb4444qaZBh/pualZci4yXMgHJAV6JVnjAOMJsamTdbui1X3LfyxnIvsrs5RRnBtfttypu6GW
SJ8p3az0/yxmUSObL8oWkhbGva0ob5QH0NTZ36KxoZ8eXR8JLY4p/izJSxPK5OVSNgLVqBD4Y96x
GM5R3obGGqVRIYBqmCVv/Yrixa2wHrgoRczYZLXpodN0Cnah/+0aEueFBHVGb8inbchyGYTd/P2Z
id3io4t3GXENSKqUkTU3W3w3OQtj+Z8fGQgNLeAN9Y/YapFkBH6laoRxbQxK6apvLzJo+kNxSLde
YTAhaXE+WI6/Sl8DMrBDzLYDVPj0/KMy0eadQ1pkKsrXA9p++eIlEBJV5c4azB1Ul7UN0VigBie9
SuSvrt70/7Fk3S0y51xq9ynUbdjKJiwta3cQ9Bm5cZnz5wQeE1+u1LKaUuHxhX9XYKKkFmTXjTOT
HyIIwtUmSGmH0SCDs2/d2+YnQcG9hJO9mU/czJ5LOT9Kc6WiJjpj/jgSZdCIo2GWV+m4H9v5vq/b
Xfcl5AYkCzEcCURHjuehSwMMmBpSXPaSarcChfFQ5aGHQnK5nW7JpXm3DUe36eMio3U+O5nRiS3m
vXzLkkv6+c23Y3VDFnMnyoNSsyY5R1gDviUO/hxRO3tyVVvFDMxEkCzq/k2Nk6DfWGGc7UsqGiNX
ig4RViiLnXckZnx5ZVtIde1kyVZ/F/XXqivH8NdlQAzfKtaJNyFVtoZ/P8cTNI38lzWfWPourPba
+H0lD08y7LCE0OQJrw8pAJm12WG8PcrvX5vQNKzZp/Of/4J7PWKpwybU/nCs6sTEoWTdh34zJgR5
UDfgi/aOgUG+GcYvbgqKp1+wEtl7ndia1MPbzOdFtweD1hUBWPM7DbNnJX25TCgXuxJWDbug3d3B
8P9xohopR6BKWpkzZygbG3hfCb70HVStnYVdAcDPnQbN/6MJG7DuT/XnysqtdPRn6CK5a40yvi+f
pSfjHhdJwJ0gGCydGBd4fDaMl0aICYEJfpEx1b1VqktAy7LHmrOw7act/6+sMKuQgz/QI4Zt6vx0
s3PJdJLhpRxigUJGAqJf1sLZjk1aCgvEBOH8x4DrrAPWoU4cKJAgg9Czi1eXKNCH/Hx7ZC7O0y+D
4YWneSF+1MbooZQVxgqyu/0nYbWvsZm38jC9jek/4fjRvduBOxY+l6tB33A9rWZf3MufvD9xKFUp
dD0G0P31frNvZAFL341fpg0Oh6A+e9lD3wF6+Z3sQSOPDVm1NWlU6zTqrWWk5Q7adsgfey988kBn
yZPQdI17lYeb85YpsotQ0LpnKrT4NVuaiIhtVf4Y17w2sc0gQJUXjG88j6xjln/a7XZyilzTYxVL
JK4BOXfP5saKLnKU/NMiVnAwoJsH2wUwLbTrX9YQw31XvtyC49UVbr+FTgmCwfqT6xh47UnuOqYO
bvsj4/3ibuivWNRgbX54H7Eq9e1nc9rmebSypb5ccmyE9ET0NxIDqt8t1oGRfgPYsb2TCUZtDb6k
XmXf7e5uR0ZYAQrbpKtSBDPBgOITpV+TXYHdbdPc/fDB5WI5OxnJ9UDgf4dGXdb+gAYnirav2nxP
K1l1KYcPr1X33CWHYz4cJGMyEGx9bzrmpRmsbjOhBtd45mk2QFXp/ox+ZtJ4fzS3P1uoXIaSVMk/
mW1bU46opgITpCpWA64Pm7ZKzd/1fgQTYQthRNNqPAh8Gdp/Xpm9HiF/vx8OGXPdzIHwcqQ75FFL
mMX8rSFdWrrJ1GHW/tv1Xd7iT9Lp7E/9uWctKTpAhmpzSyaXcSW8oT7B/SQi9DdwlhKEaRyKFA3p
GxbRh7nT8TLh9vmTdGT4xVVX6I9BpFiBzjO6ZnaG2gazGjC+bHXnn+GC1Qt5aTh0REaanmHrbOWB
3wPi268YUxjXA4nkZ0xlJE4KXXf8RYKmULb/YSowsrD704LoVO/TPNXl1rLayi8B8CJAsYcslLq+
o23n7F+sM7C1jeLTUiKKATuJlAsaXvBbgF2gunakKFVHuXUCmkuVXszj+SKDgpOP/1E/Yb2v4fr2
ylRmgj/92/XH/Re5if5kFeQNlTT9w/Aw8uIXya5MDI7daqoRm1q5WMAhBZg8EspU84xoxd2FCjwt
3xS6ta6P/nSm6/xtyLAPvoimg3h837XGhTU51VmtAluE0ShSwS1czz0bNbIUIJf13HllyW+VxpZW
7n0F6NA/Bvz5isQYXlFADLBJMbx6zAVvAu006GJMKTa1cxxztCsfeLJCiOG/IGikNmHdOgDkzaRa
bjmpocN9UWTjBMVnGZLYi98whZnZzvbE34Hn5Jv1RSp1Pu4AbjszTmBqOY4bZfuy/Vh2rVHk7hdZ
7FhLWkb0EhBGm/G7cxgVC7hWGQKYfwoGzEkrcwvaQkl/BDx/IYyelZ24w0mS3uJDiA/Ls1hTz6GY
umHNszSOmx+jJu/NDWsQpFlNf1cz2CJBDJtvOue2asVN3bDiCByyE3D9WFF2LokqabjTzKBxPZ0x
zq8sk1hYHyrxGxtprCUaMg1Cn8SaTTqycylHwnLJKSInZjYeKN/ezsUx5FBAFLXHDeqCCIlvgIWt
LBXV2NJv2bUMpEkSJs/QTg9EaU04YUfpPHbp2xteoUBcAuEzoc6gu2RSNGOgs+Xea5CTArg7KgUo
egVYruZ0n8QAUsVTKQ2ItJPEW+FmLf0LCqWVSlTpwrOEg2FNx5TKWClmmE2wkgD77/zYxYnV/qUb
ZeoQQYnGN5G3xDHvQ5kdGFRW0Y+E9Q9asAaxG88AzjBR3kKQV0E90HhsxjOhCHtHFENP/5LI9TG/
5BW8x1+GXKATUOCjBTzQPzOoE4wLVr39Cvu59dTfWpk7lwzttocz7qApd6yym1HlaUyLShUnFlEL
vKOA7sXRU/fGS8Cz9dtJtXPcjdwOKWKBwBQZOaxb2klqXUEpfAXXz11pUf8Y505S+8q8SHqBFCf6
4br79qlsSAr/BOtR2cdSYrvVdN3Ieu2AM0yt28/PUKBnaE94S5Hby+Wo4+xE7B7hw3rik9ghPoUm
77RWVOF5I9+V9CyrMHSWCa1j71grfQMRfdCjcfNslcTpdoh04sTdAFR6QfhSKUZuzih27Lpmy8Mn
ikfEY2MmPVY2WZWD6OreHni2QYj9vm2dSX7VIB+CjnN2rGYJFhx9KHRsiiA2kB28Ddd6hnzpAA4T
92fgV8Q0bbXIcJyDzollE9G4BJMXDlfHcVBPwTgz4YzyHBM4cmIsEFjwAHJtFangAqS0/2tlXpOt
PNR6cOAJhd3GaZhdsqx95eCrfE1XFDLBQ+MCt171pvo3I+C+UmKioIn9ziG7lrEjLKmPZNOZMTmK
Oxo7hGzLagZQIE4bmt6Ze1ijPcYQ3/R6N8vg9XxwBa7Yt+PwpOQAq/YiQfUf4LwkKERsQSw4Mkdv
DoOw/85g2LaYEH+5svTBdRZ5pwZuQ0mjADz8kvuxdWwEk/8H/UYZP9zDUhCr+Ys/FBqSDPe061Kz
b8n/HTbS1073OLdmul9wimY/NAAEtsNE97096kacrXWomyHZwMrvnk/5UgWg9XgP/B7PHRubMw1x
OZUOK3aFHsy9Mjnd2lvIEJ/uE5jQ4afJ7tnn+YCRsK1Gfd7CXhzL7H5HFVspkNmTUB8I9S4QMGGF
azW2MdRGhckls873vGIGLvh7tM7yK9TMJeiOP5qjucv4dYDX7Jv1rqbg4cPpoljh+Ul8pikdIBlq
ZCsaaovet2GjFsmLAz4lcP+tYBC5+Xv7y4FCjHpuElEqhMF2wvFWp6KHztFlEfHPVkDrDk9yEjSo
4zli6Nc7a1LSFcuCKCpjznSDk4/oSPtNMI8DqRIUjid70EGVISWTXa8p5GpfDpbNBHrSaz4NjY1G
gILADyRo90cUA1IdDRKZ1jydJtuW4hXaynxuNHLqlPA/m6omGAPhL7ljqpEXtYn0L3xu84dT6mGc
/ZFu002HdhEhjVLKmI5aVdMhkOOQQUjJ0m9PdJn4odiaGr9gDYFeNLk2S86ZmubiOO8g6ueXufu9
DzvnbNhFOw56a3eDEllR4/Q3dTgf5f2H4N3b/0+C+7XuWsz/HKw6wZmMo6tNA5OrtCF16xmMIYzd
DtDlztvz2XfS7aDzreSrlqGkmDfiuY+XBIy4e1s40S/B3BKYmR9UPvR02dyBgANRik4Y3a8o+hW5
BrZoTdMy8J9+A07TbK5lHwGeNyyXgXnst/EXCgHUb695mAeTv5tBhTqVoudr9RI9Ov9CJWaq+Fki
bnvX+9jK0g/cLpDKD6fb4E1yiuOTzMl2u9UrEnmmhsrbx5ewOLssmj9vw7tyh6ZQl1KYxlczdQ8P
KCbFO6FiWhyiuxUhTA4O7AP96XcbtwQnioPYm1NOqPZkJJXLxOgitjNhSGP/i5jRcOcQNsaAWg/s
5jhuRqgF0P+NSW0uxWarW4GjwQc0jyNxmIO36mUk/Ka0Z2ZvTXHLun0b6shY9PYnAyePb4Qbirp6
U+V/u/q0l1wiV7H84FBkA1oCj4hIFRR0xd7QAJ8XIzLWCVVcLf4xNxGmE3NIRYn4B7+oWSLkrBbJ
799nhWPEK5S5rUo7+T9NZwv4kxIvy3ERxHvgYai9rABmWg0bIYZYm1UImWjIvWPHgJYyeQPpeVPR
s4UUBa4gdizffDhvDKFnP5Yon/rIy5F4Uvf9M6C5uYqcIq/g1guqFEJUXwVgL38ICyaDod5RbNec
MAwyzLDe5ulQcyba8mqeB9b8OrK7gdypbs5SdZMAEE7It/bOmnmN6wCd36K9xT6IcsB5Rp/iJ5w7
AMOQSml1w5FaxdZKeO/TYSkoeRSqB37vff+RKcyX/XjXyQ0Y8YKqhcFucLElTKhWHShfyu/iCGsF
MpeJT3QOeeH2JX5pTNdDcdmVR0MN5XREaP92LfAXlnoanHqvAP2V0684EDgsfVnXkngaoGfhSAB0
Qv7VGinW8vN8xBnWuriU8bpf6oSk1YKcZex8LFeCoaGjuD9LKe3qSFHcqNm6jVxuxaHnvrRJDLi0
eSFKBbM4xx0yKEiINvy9q7huqe1OYeoLxO7pXftq8WrnTIss88pdOCCB4r+AVwAspIVymRKuNhxT
aQu9HtbWAJby/MT3HkDsrHGrG7HtmWCX3t0L6zjcIxWtgQNaVQZy3wmlc/2KwTUUDdbba0VzvPLb
jQdwqxE/Hm2FnlQjJ/dxGZrQCIlkIqmopPw+jhrJTl35do05NubVP+clRQE8xBQI0YkpDgDhCggD
nqrFC7pr/W7Opksm5kHys6g6FUMWM5zaDUNrzrvkI1OU7hRgod+ln3KXsF8tUfVAkl00aRubjmVc
92VWTgv0C/rAR9R+o8B4tz3I8Q57BfPNQpZuRZiQ41+Btv16ucJdW3RnUNTHy68Gc/H5twGhHB45
IN8t4dqtciVtRwbVnwhLgv77v5Emb6fg3mp1SICzZNmiIk0Jk4hWIaByi66XMucAJd+73mLyvqVJ
kP/OYlORmywVAo18re+9zcomdy6WlC4bDvwdcf0yPy+YaJISsq+4LMAz8lFkWzY22ViX38OKdSiW
9clVZJ061g7ees9Z+qpWrnnE47HrFedIXi9k7+2BQTENwOA66VLi65kBF7R0kb0IhDt7zipb9Bn9
PrMwjZFSpo4FFah6ci0rAJAECIQMDdiw8kfI4qtrhnFO0SUZj/QWWZK0EpDJECAqK+qsNUXO18h9
okef+vbLKwrPTxMfTb50RHht7ro8pS+XYR4/PeEWHqYwtr7VU4sKJoqNcUXhJxOJLLK6Jp8sW5QY
13KFzS0tQqv1xsjdVcTSmp86WpTERzPbms1ExZgDeWUDajHLNskhvxrmWxa0DbCV9MYpjttjopHa
wiJQz0nKAf1U7m+iu1HWLlq2B6wD0pZLfCs0yOeCtvDIuRUVTqTCcIHyaxc6u1qm5m3Adhv2HCwv
NmFtWCIv7IHkvs9vEgAD0CE1J3DxT5imQxbESAkgdVQ7FsaMtf3mHzR1MongZvVXoKdlBVQ+UCYa
mhXqhZd03dTVxnrt/8nl3hbvGweMjaV94B/oDUWL4a97sk2mLynOrY3reZ1B24dasS+P6pBxbge/
fEP3YHccO1FkkSLsG3Q3N1+QEeFqhpDOVjLSfIJzhKrxA5XgDC/S6hFjpps+1c6bdSqtNfLwi22C
vJIM41dEe3y/YalUQsJGd5wMCCDLDN6NrJpgVNK7OgYSGkpRiCKW6y7SDFKSt0HCP3+QepjbSxCz
er1TJ+HNhJPwewF0xmGBb8/t/9PgjMpbKGgJ7vI5rEi8WbFrIARPWlhDX58hUlPXpjMkeR2zRz0i
7DbIbINERePkt4rc06D77rGBSc2uxaXOUI36b5uHRrfyWqMO8rOF+wfxWMSEcD1uQhjRWAkJx0fV
O2Bptn+FNkT8lYZ0ukQ0VGoCho6WG0k+X9eWQh5i1CkwFvrq1bcGmF6DKnJt6f5bvLLjujvoZFQZ
Gtn7KIJgk3lcXr5Ee/qdFIimU+ehDe4BmTYz9TqbbJNTP03bGnSbfm66luKtne+UiLtlKWrJYysk
pHFeMIdVMrS1bmp/IfUf9daSHxpAp5hFP0VqJTik35BVyoXku9pT8RfqSFg9GT4p50YPgXb9oo5i
tC3Ebxuy8b2IplA456tMUGwjsMRYc1Hc5LXabXq6G+e2KsvZq+iqdUJ79w853c1Bik3dVR64uYmP
h7BL58wZ2Ku+E9AOJq1dBCxuzlgbfMGOjtaw+E8kx8G4oE3XrnuIJhG9MJFFoArLufblz2JYTpND
UknLdt1lox4Nw5pXrp4HcJnQIRapfV9EiF80uljB0/baST4L1Im8U7o6ItM0yhtxpsOpMpueLfy8
iklOG3/si9UVCSpt+DpmUB1AN0MmY+rfBFMqKbypXFh9vIjb0TyN1xxcXtmekqfQYgUUBVvH4Oss
P+RrS6tE/s3mrrkFiA5Au0KRDqtDzGBT0jPieh5UUtFL+zfIYrSr7CWy1axbxrHWdJg+qut62D24
a6nitG7uhLCGYkyAf7I3jVPnMJQ9qeMVRT6taSXDi0bIOhItGew7tYzjPglpFTlQzvtzCs7co230
xLY6YOaQgZD9DNykmLezdbO5ZfgfYbGXV9fM77MTcjO51dxBJ4Q9MjpVALkzW/ISHEPOIzlMhO9H
mc8GnqfdwMsEpJ/FzCuxce2Oqqq2aEzla1MOCxLVY03RTwKcToS4MBvdY0uBe9NRrK9lZgoTfnRu
AOjzJAi1tjueIk8ITSIdJ1C7zBLgF5tyISDu3Jaal3Z29pr7ZZtpdULzvPKXPWGTLp5KzpFa/fGS
QfD2bfkUkAkH7EdaJiI7wyh4eCkFjqcKKa6WeMbkzlZpaOEIy3BpeR4e2EyNSM8syaxpOcNfbNQ/
Qtuq6i5gppWUP3mOxf0P3CQXUh/q1SNAWjGldAWl8bhj0yNNiGKwiawdN7iEWa1uqgjz13nsujUG
BEQpvKxHrzHcczTjh9l2lZdE6wiROy85h9Hk2t6dA0SG+OLEpp7jzCgpWm2t3Ryz0QYmSP+LKO0s
Ztin64fwOm73wxyN3lqM8sO2ElsQ9kNQj+VBaNzAulQoAmhWL/kXoHwtsVhs1qjAhvH4ng1nQ4Wa
e+Qsd9wm+CqYYoQqiMG2gFjTJWHJjRP4XIXkezxUEcYXNIu7k4IPAqt8eVZwb8alP6j2h5Oyub1e
fAdlAVPje1lmU5r8KJ/UcbV9Uo3kVWyRMfsAuvae1rdr/uMdwVlmbLeGQeTEEUAKN3FTfmG0ebTk
ZZFCXfQZ8U5EECB0QJvproEaXG8+w3APR8l+WrNbOr6wp6dcWIDXBftXSWYzz0JRJOfHVelpkF4O
JYCcj+qdINb+mALtlkwCYwGsC7y2Anf3xPv2LOQzgpoSUSBT40yGEGKZBQjTKQkFxFHVKibJ0gIy
n5x6sN3/67R0yaRndJA2kKUrDeIHsOvubi+lrchR66qOEbu4I4yBvgGq2pY8wWr1Stj7hMlDu+Op
BfeNPH2bwIerIvxhbRv+B52P6HgKF9F1b4nqgE3F34Q8EIqL5jX7OqibcuULnWi7It7zOHOkBpZY
nUpmQaJBTVBXpyKykV5h+pKgR141WWg9/hOlixgLEy1ElF+4waR3RsWSZtbR3TK30XbRbr/mfGMt
EVBULnZC+wMu5CfPS1WzPbHf3S1DBimaoTFlSRU2m4wVdsjCGxvOwMDWL22eIZrzshCNDeDpq335
dpcbHH4WnW3b393SKT2e/M6D5KgcRBTPDQ4kH3gFkzHD0XZDRx6ig7eafbkpWU3+X9tLaqgXMcz0
8LJIvQRkgTLUhJKBgxxojyux9xqPlv79qt6sYtaBEMq9pGWGymV9x+TP32Wu9fa/GBeSc6CLxoLh
BNdyLsA1NYNffeOFdJQath91g7xR3uzDyzrcNLoB6PdCRJ9Wlc+zKhlVW2thg9AV0Fs5YKkSkboa
9nbzKUdIKySXX1+7yqm21LUQQs+7UmlLdZFW+B6lGW5/VP2uawMcpOtGjVhZhlkuDG4i2HcDWWUh
EHaryO/czl2migv1wdqhZgQ7YQnz1Ok7Q4XYq5n6sj5a6GbjcoHV7B6kfqdyBbqDVHmRxqczlieB
skeYic0tZJ4by50mTq8FJUp4WjwdluFBeOyU/bMRZ6XuB2F4W6MF6aO2a7TM2IJT7RH39uu4NOrX
rsjjMUBTwDDV+45F2MwYgsQTfywHb8isNxv1kzS0nx7zBr7z2rU11iA+8peMkz/lYMxqDECYTb42
rocuUXDpsBTJy9MXNiLhvylY1VzCAGtmHld0k8l7CavuP/wQ3DOinzc0QFrDtCRpKZPQ7C+gh0yC
E81d7G7V5dRrVq6Hh8BbTS6wzDGiPSbP55LJexbBRUn/yJ5j/av/3OdcijkYjaHB1eqHMeiO/ZAt
OLT/zRXYTWrgvAp1Xvpy22i8pjX7lmdP61dd9Kvi82BVsKybmKWS3M6xN7/2A9j/EEYWeaNyp0YE
jaOXaF4lgFSgnNDZ+xTRQSQU5j97ZOTjGRDpvyUvsG0RMWhkXzVb6wvCQbeZPenT/Tu4EIcU7S5B
B3rPb0FqQrheHyAS3qS/LR+oEzbggzYBG/j5RcCtOHUyVKdrlelIXJ9qUYGGrIKB139ee0//18Rn
JKvF4BVs0f/Pe3T/XCjartA0CzFEWnYDi/nF1HICTSP4K2WZZ048ZUT38qBWPj2grnRBDb2mcylP
Yng2sNFqwVOnhTGGznvItyx9s6QktSUhaPaG0Afq0XkFe2TwygzzTstU4MQaVhFugA6ReeZOoiPp
CcIsKKquSrTDU75PBHF2oLxfk9Ndiv+DOK0OSAeAJx/USF5Be2/xhfzkqkaLwd52HQwShixYbJVo
GSNe5iBvllAqcbjaO1T5O7QQxwV2WA15kXqG+3O7OcAG+fyH9n7zFvhJqQn3Pl7UyergeHpGrqdN
jxJSX6T3dP6qtPCa0czYbJTRHsVlxT+CAZC7+ya+wpxohNUEbvIT09d9QT6NaqY3g/oROZ7lJQJs
f+JKzQkR/08qRkHFKBkSfswQWMUYq6mE2D3dC/6YtE3Z84TVmL4iyEHXQydTe7AJzXBCWr4/qC7P
QmwPQLVmeoyhLwi4SfRoeZU9zL6gAIxbWdHyNFXyb/eGrYSTP+ac/uu5M/81lg60x1HB2RI4TGEx
dax95gacB0oD6ovGPfgmgH7A5anTTtjobRN+HNMWq402oJ15lhm3NlutYsTuNWPuQTtgrjJjLj8Q
HlHIPD1fV01ZwiWB/R96NUot1vDUhjjB2s7dZdizLNi3e/Tk1TozyJxCPs9pXWDE2IxkQE6osvdf
/jrqAxuIQ+6mCGr3RSjPAUIw2dDLKTmNJef/y2DRIgHiIPiepDDK8iR/xluXll+ClzHZLNABc1Sj
mrHM4CMFvdprav4GtI0LIQW9nb3ew4j0hoBWEl7n8NpUV20LGWKp2oqi3QOGcc4N4lYs3IMwYgqv
growHWEV5Iysktn4IWEpfu+w72PzAIET0Sl54MVLgwGthvAw+YcGWzDkMxbXhfUkE0t7iP6v+Q6I
oLD+17vfVXmluL5eQmeuHEw4r3eX6GK1IOo9dfhl8Kl/68q0b5wmrTKqp7JNZEgxDNZIoZks7Da3
MFXuBxttaXynau0isQNscZhSsru4GATZexggvBnL0FCIv4fyIzpVGh+eizAg+FyQygp3T4goX9BW
uCum4B/WaQAJQclLl+U4pb9JpvPLU203rQqNENQ3EYu0idM9H+B0gXiccR5sbVeTDJzH6khwz4ko
/7bTrtf1PkGAFehSSMOTw+Z0XhO65KuMxaLfGFLCsSyWJJ/zNoZvkhj9m2bkkJiYGjHAlh2I1WGR
MxDQJSyRS9YV4fXKsLH5cHTRNxCUL3htAywl609MgaGn8m/1Na8+ZqiKv00Ff0y+pM7QwlXNq3Ld
D2b3Vjzf9yJmV8Gy5vRY+etMi6PYnqdayPrpiHKzHEHpp7PanaQYBA3iqML3spfrpvvNa6F587/d
XNTmN+IMbAWXGRTbp04+hyBnXPkizb0ytCnD5zSoddsgF9kr4/b+wKv5+17nmi7BNGG/NoHncI5U
pk5Qm85ufHB1cnY2BuFz9K+AJEJBmT3WcAq2hFdUL0IlvkDc++nKz5tB/I9MIMoenIz7yqAq9+Ep
CB8a1bLWlwlxtUvVv+04rakSh7HZkjCJOJLdc1lcHSvXxcyCY1OLDFaFiSSvjwqksbFHViSx3qQ+
WBZG0aALjbbkc0tlnVAdWhBjihe2iuz46u++vUA6UoNkjcz1qfQTt0r8GdR1eFXCMeKjYn38INdV
jLpHuyOZS12+lhHzodQyPoWHQdnsi41EV+AoNZVT5pfcFNT/pqbt4SXedsz8IuAuB4dZsFVn40WL
j8Jax4AnNjUNZk3DIsi7oTzWLaJjK8ch1qC2Dqa4btAnkKqHbS4jthIC0r0CUAxgf5lOmCT7mx1p
vD/iHEixEer3sh1IUAY+7vpv+F13PbLoz45of6RDLqusvD8IxHDRU9SIJ98OWCMlaR9lH9K2mhMh
T/E3FDWd0OjOkEAjYgjWC/q9uPArBu2g9l97ZaX+cgwAqsufzNlbstPURiEeUxj2I6MUitLqH6Z+
KT8LxGoSzcgVeF0oJWpF2FESrcF2FbFHRECCWk0JHNUb8z1wa7vFjJnFHeJNdIX/ESoTyzd/Cqae
5S+ALzmCQ0ExwXdSQbzV94a/51joQAeAUldp2Z6zCx2b12hArLv3M8MrjfICfvovNJDEi8bMxIzX
r2KsdFh5ufwRIP3PsKSJKjDhN2Pc3HI37JK4KehqreDKzVBrQcTfiTdB8dUg5ScVSx1yyAaB/6JW
rQ1oxYZDq6whLhEJ/9QEjCoviY61ZyF2l6G++Uil460MnzWBCCYbQTTOz6uJrsBr617OhbGE3NMr
RBTB+yBUD9LjPhXtZeIc+EjCyO6JsloIMk+JsnW2pRRS2Zq+04YFUGZlh2Ih7p79MKpblwv+5mNL
ZoW26E+15ZCN1JLpoN7XsRf/ne6G7GBx7aeFlHmKATjGoTJ7AW9bAN0ci5vVHLMmAAW1jBUWGuGw
MeSoDLwUVG9pdS8lUVJkuLnuqvvo2h6tDW6VCbXw/FRtZPijGb5O2U/68UBuIbPT8iGh2IXcyhGP
yFinQaq8hnsTy2EUeWm93kTzPqUFPrwT2TSACVM7Bg/y3soyDlN7x3TiSbjxpDSibmV+HugOFSvV
mHeihrlJcKR01W5l8Ulr5RLqurgd+Wpzzqor04tcaTbFjHIN2Nb66XFti3TcBr3S93xm5MO8c5Zl
dguKFfwcRr90a8Cw21jU1F3Oi/AkOILYTco0BXzGwmS89I9YzmmeqJUhqifLWh08gbdabqSjBEhk
DCeg2A7TNNbnhXw9i15SFVkVoG3jKQmScqg+9NUHcVTOQwDWzTmxghEJ8Si0No8cqTTs+QKIFjML
xi3KNm0/E+vGHtev08EV/C540bB9azRWga4EtFjH5/RdZNMwm1Iu81Gdbw5XillEHyUx4YMVXbyj
kgLs0ZGokUcI/UVqqyyDOxDO+EOa64MqRvQkLj3VWzkGnMb/l9CvNmaSTXcKaXiNh5QKUm4M48J2
G5iWk/IpnJx5Cm5ajhRAMmqzteZJ4sS5KjlJTeWwfWTWnjEEanxNmhOJ9auE76rDKOAvgJ6BlKFQ
pSEF6/J0rmKZEJZWB/sUQUeuuLH5FLYe4uWY2vcT4Btn+V7UW0Bt06spCBJ3FvQaKFHcbUlgv0WE
oryLudN3ZqzzqIibRJXWI+n5YT66rEiPC72WJmyXYivuWN87x73MdhkrfOZL8pkPGyD/b1AX/gVv
O2VUST5CgOG8S7f9EFswUzyuRB4+n4AD82GifsY8HeLPDPgqk12xyWMDzE2SfpjkHsieQCT/icFj
qxTva16BaY1B7lbu1J2GsL3agsmz3Gan2hLEKs74H9tPdoU4evFjj/olqbuit3wjhaGkJPcCHLmz
UkhTSF4QvqfJdgnfRKUNNJBPDM31ZtK2yJwUWaWmokDJ3O67LHONFhpDnxqGtgqeuqkfkuEBqieB
3rIb6WImBjL8N2CVom6HkfNtpR5Q21+UufGpdcGkqI6eLhI7yIiFlDjNhI3Q3BboCGUKIxwF1nN9
EpV8uyySN/hRQAl09Hek9my8Rw037ku2bSC4AOXoWXrDXGcqxoF/+i5trl4BnPkBySysXW6pDOyf
Z2BX4g3UOzJsu1zVJooWqhQjnXxwJJFNpKlgyFmJlPp2ia1r41ouZdQdeMDZ42O85Rr8Cqc/LToe
KgFczCEwoWf26v6Q3EHhIS+OpNoC5gLrO0QoxoW/cEJvFI/noW5sLwCgnOHP1JxyEktS8QC/a3Hc
jeu8kCUNS9fEAK43MWNfYPVcCHgflFrxnpYwyRvaoUwHZCKhm22qB5rGdQRWXXcqX17Huu2nZrTM
SOwYBKkT0KvEhonM0SnIVOsE3TAPcE1H3025jIprBLTcq9oyXcIe7c1sxG/tbQDoVU0APClQpgWy
kVJYQ8mSk5lEjdXzmpJuwx+w2nhPn/Fc2fctlCiQBKBmyvxu0Lau9pDaITA1DMPvvUdwkeb6BwRk
Eej9TZRbZFdRNeFSAHQu/fl/2lifiLxXXDCpTzXCcu+heGBAX+5LVAFcEld04JV8TpCylpnsmLrW
X1e5MHM/DKmGPx9gaYIjLJL/ihc6PGYkKOmWkKR/dqkuiECpXy7o5RqbNgv/hfYn9q2Hd7xZrZ1Y
E624kF7j3/9QbpltQdUDrskYfZXJnyGDddF4ZxupAy1K80sgewpS+ERYAQ2lKnSml8lnmFR15kWh
D0/b2kf22ipQUxcSBjanRiHxzQf8sif8bR7fM8Xz1JzzEPZj2UH8nrMyBugBCdhBHtEo8siq3o3x
OmKGHzjbTUzK+r6Zs5tNMpClTBD6+S5WsYxaVRY4LqiWyVL5+i4UbVBpSnG8d8ZGSF8jUNSLkLzo
0+CFXCEfU9mLCM2G4jCYFbKXiOI2YzmY+RRZo8GwAfXNPNxCaDkIswL4Klm6wBhozLD+A3f9Nevx
B7gCDXZTeVUR8qQvAtGLMquZzY07lmF8ifXqzJTkRZhOB6Wo22LQHB3Vl1ToYpmoBccyzTnSPOlz
cO92tCfgUMuvZ/J0BYTNKNb5Nabh+JGUjocOlk8Ge7a2Ry5F7tB4IC12oy2UuX2q9I19VGqzZn6P
hCtiNDZd3cH+OyWPmm5VsStvx/E1pqQEoaG35JYrLSBPl1QNGDjVc9JaJWwVsm82oS4hjPzR3pvi
G0hhg8JfduTdeckwVJe94QqBc1ry7hPynX15DnbC51H183NCdlMcqUjSmw7WNaP9CRS7ZHnhRGcX
q10C5fB/9DcqL/6exLjrDuaa7m035bEEQHxQp3DTajgFd0bxdtmPdkiHhc79/I6YAOsQcmtHoIUx
CQuHOKlFc8Muop6Ii2Dq9YNrfUHf+b3o3VhAc+lZvd8n8fxqRThokyWHTRB7JPVDgXhr2o/INLVD
Sy52aGH+8c7TzIBknudrOLsAHiIDPNPaEwbviNcNXjyiGbkXAByyMM0R2n/9CZcg6cmpGWcWd7S4
sXJA7zfgcLR/r70944pJ7BL2GMQQzMyipPTfAcnnTkmG8srjOHgROBFdWDs2Q+XONv0/DZWDaqwb
bqj+RWre/qr5dg/Lv0alIZ/g7QFEJdkuh8RadgJ7vnrjEbZ/M/+6/6NOi6OqDgkYTcYWVCp0bD+m
fYNLvmL2yrMqECZ4awTZAsqp6Y2rhTHY4vTxdXNVzVbLzO+gNC64OZHNKtjt+Xq8aWWSsszMXRVv
Jh171JAxduW93sK+5izJPBDHz/6ttdOH4p104hePVfxlXmr99Dbz1hhfQj1RH7yeKb81emECSEnq
dNHNvwHn+ZFot7TCG9oJNLxE3OZinW9IoEa+34PYzlGxdgffoYWn+RYIgLiXv9zj6iEMHznA9tBT
yqFVH2gyc2JAlmWXhETVPVcT+mN0bCZIxuh7u6mb9xQoZxqgB7Ioekeat6kqCnNy/VZON9ITI8BI
PM9O03V98WJoGLoWi1i7k5o57p/qwATciCn8kntmDUYoqsC/1Fg4/+SyAsqGba7T7PesLYlBKNLp
Ct+e+zoQ6XrFalTawj/a3mkN1mkyVWgWk8UE6VIGrz5jzkHTZmLvY7+es6/ilVvsw0GOhcyT/SGc
fWKPsS0r3BtmsMKlsuj34B7pGekGU6sLCbph2T5Tv7uwHUmoGhhSDPS9wi9qVSaDIWSyOkrvB2cR
Mu5rmpHcyxrl5TFY8rdgghQlVYNdRpo7UOv+P4wHMBPfpNjA3STdqhcSNZGu/kJJ7JR1fwyKQzVA
X1zQB4wE/or8ZI8SoJ860LusHs2uHXiwUd256gDLS6nkUw0am3B2wRD0uhlimCJFgbnEZaWR9pLJ
c0tYWuIw1g8QpHg75/CUmV+TsbgNpPmpA5fL8opmzVeURGtQuwG4MIn56hw07vFUvUoNVtlIHY+E
wLwFe2JrcGya8Esb1aaLFxdNw6NAAG0l06fXb/XoZXE8bjcDRci3K9BYErCjhPJGyUw7i+8UdOUF
wRZelw0RIF2U7hqiLyZlZ3D3rlUVVXpAtmF3Dbujzv/IRDFOi8+NyGFFCOP9Q8uuH03JCFB5wZj4
rZNgA8GoN/wZzC2c0V2XvnWLuzFqHNCBdKwLmQ9GLiPwWHytDarWAC8zjJofvEMPQ3rZ0MQMK3nK
abybpaTHA0KR/GyKC2WwRDiayIfO7C0ciolxrXP+N7zxTpE+UrJaJ3Wc7WEDnBw8ZKjwvJdzGogO
0koQUL3KV3rWIJX53Wm+w9oYbBqnvPL5pgxlO5lu/rDcm2qbLrMhmCnJ6FKinJ1bAiwYCiIP7fdv
0T9lZ5qg8avqrURcTjYqkSe1eaGmsPD/hWNYSym866AxKuq6OCSra5aDyjn0su22z3xocRYtRKqg
fLsQMcDVmF6cGEYgQ2LzGE+/a9CyWpMA4sjKll0dwoE+70JE+uCpF92qQHHyWgpxlUPE95lPjIGF
q6F5VBHRqVj11mFLmxEZn6oj0+ZY0MSq5WjIeS0OHqvXbkC9p/Y4vUpeoTNzoKNaQiOMMLRGBQ9V
U+Q2n67Rl+Upw0te/NrkqgncnrMmzGJ8r16hEc3ivUcwI4GyRFiqfWTP20UmMF8Q2jnV0ZpKd3jY
sjwqelPEVBDrb/VZoxUbX7rUXCMDJ3q1ZOvnG8c+arikVjgcFmKW6Jmhb9EUREnxgY/2MDPZD+3y
EcLDN7KtCwr4+fXfq1Ua0gaP++ciPHH8qQw4pyhGCjM74ToMOMgvVm66nhlRupizwn8MS36wX4s2
xSXJAdIcHqbIp8TSl7fyKXpw0IR3MF81Nqye7dPv9my3VKbu5m8XQN1cgLWVP4Yix6SwvQMThwQd
B8OGcIGwMJx9M2MiojP4vBU3KkkcsPqwpddhe/bY8MRGatbAHcCLqGzHXWBURbkR6oRfYD97Tfbt
KzkCEF7KsGxcLYOkBErNjEmcLvgHqEqkY7dNBAgJzE32t5OPQxh+EPa7HqQxSxwdg0RrSrpUmp9M
dECtTta8cO1gyActWwd7dfuOZSJcr4BpZ/bEoiHhkxgsDURPboWpM8QnWvPRpSY33PxdLDFn7Ipq
f9U0x5i5Ri3FvRa1yWC6MYpoKSamZH3VbJhfNcyCm3SZxgydOFVUu+xs6CqpoBQMiuKWJb4D7jHY
o57JoYjnov8UMaX3/V0h0wFjXKi8Akbx/bRcbfoCvEVQX6U5qGdsvGxDSSkW8sfQagYNLPpYUiSC
DhvT9TjuzcymUkoDujBcrL9xLvplrYSJFWcRRn0X4lSsxA3uSALdAQBPeX0gFliLhHrJDgyPkCZ2
+WbvFI49/9cDuKh7vmz0xeVz/sDz1dFSMCdAHxPKjNOJntqKDE0TG8nSeqxpil5h6cXulosBELYA
6FcotdObUk4WB0XF7cKBV1dzpXOY0urU2qb9lIuwig4J+YsB52tCfkS9nt2RBhYLAUK6lY8Z2LeB
0Af0I77ASufGcxidWb4r4GaJWtF7x8JXTikRE81W3ESuFvMeuj37xFdIM8WO/fooYzhnBX6usjt4
hoEd+OCx6gtPXxbh4UrpWC64HkCbwl6d8v0xOlW95kEUNoEtwGZ9xk7wzU9OF1R+1x93OymSo6c2
9UTSxk9qKkEX1AyhbcoXMnwUZOG6mA8v5O+0vDsnNh+FlLXbY4akd5+BW1SvNrCEsUNzxND8Uwn9
VqcYh8Q09mPdPOtF+P/AYEEwp2TchGbDR3FgOOwObfLbw7LOHD8GIbG9p51oAlKmn84wJXYmonaC
ihtIDN5KyalLVyeD2rzKwJ7aC+6vqPhfcGe3ty8vzBhQQAXOa7fe4lVNCVDmMRi7wwcNoZEXbYzV
n9M1ViZb5ejd/exyp0FpR6Y44cwjEJVZbSPantrPZwh0gA2nWIwUVIt0u/Ostmy6KQdcVXyv2kgb
yKjWevL6IE9KlUequVaJbyE7g9pu8008mY/9r10oIPqxB11G30mouCF+6j+TrpXZqfL9axg1A2eh
YKxCGIW1Yyp17NiC3g3CoeCfUhkrBluBrD6/Z/AdlfpCQA0eb+jG6izLasZ6drlGrCuSS6ktFcxX
fXr6tnmvwWvdkddXvq4J5bhQWzffJ705oJjFUXfnd+B7a6uAxrgIiiUlg18P19az8huJ3gQXXkLK
6Utc+ZXs+yzn9TM41UGkGeE3dFE0K2jKihmwL+p0GRGjL4i7ankl4q6hluC+XwHlgT+HKtZYMGYG
jiXTDi0O2+REfyrIRNeAtWsdogbHBKxvfwVc78ye4aU/LnkOBcC8iCiEZs2nwWpw/Hf/buhJVeWP
sG7HkUmMi8Z9tsIGDakgsBXGLNLlJ8ihiBgD7kTOyjHhk+/c4yZCGuEKk5YNdfg/mnmvdekG8299
YX0YDSv0C2MkvyEGXGtkSpwx9ksyFIKt9e8X8TcoIW9AhiineOpG59JM4J8ZTRuXwkSJED6NfgDY
lqGcdgV6ARsb/JGr3NoTv9AzcaZrfkVssRIHKmJGfCyw0Zrpw7RtkaSFaX6rJ0yUrw48Kifepdne
LZSpeU8J9+zKR3hSI4cFWWob5D8l+jg/D11VezppXihziUt5QzIlCs4rUxERQpfZWnwl4ds0kt+4
K15H+FzELfgmnCXaeu9PLg55dWvP1mv/8Humfn8MHR/H1bGxOcJejRICw3vbH6T6as9AhY8/aBCD
WdH3i/mZkXibBwOEGsuDiQC4zaP9nSbEXS5IWeoEC5nLabnYoiWd+BZ/1PVGchck3X0od7x2SgOS
WKt8VOYv4tKFjHMstp7QX439nnUBJ6uCc0sCcJ0hhNa8pgjYrbgludNo4hOMNSYcEMR1nb5xqj1w
eLbRtxRscH9t44OnZeoXiBCdZOmFD12kxNnm5rL1YfKh3Co75mm0KWWG1w1p55OYSx8CFbIy5rkG
JCJrVmHVGhiSPD+9YhrlYkM+BZWfBc6htfY5sgle53tfF99YKBpKWFWfSJlfOFXPraEeh6K3eseU
pZRI5C5n80T7X/9lV9FuuM2tupbNsJ89Raas7xbWCmT33UF/rcApQuw0hDF5IkRC76hYVZ6vYSf6
SzQ4+kCUXRzI97wReN65FDYMLdam+DlMn381bXUuB6JeNX3eduEkPq7W2LjGvjxhSywRfsSmwA2Q
K2pP9wfC3MxHzua4K1LayDTwzSeH/lgN6mWLBx5KIApUIVhiWhuPGhcUs9CISF4zpR1IxKdM4lDQ
g6cCoFPq3Po1admv+ujqEDp8IIzulf2fnRWausk0iDwEm/nHzzG+s80FxoashE2MOrQ1Fd+OcK1Z
uav+Plf/k+rdFHA/1W3pVO1MKiktRVuh9S51WIjAaVbwmPiZsyW1Ckt8VE4FGbOHAi2YZ1hSlOmc
veqD7iUUV8nAoCdeLg44KUcJWuEsPcLTbpHSdGEo3kpVZTZ+vpVJBUGQOB5Sgqhu3zxSDbBml1eX
jN8U9FUECVguCkj/SeJaIEhci32cG/nqzs9SFkgADCEuNytZHh+njOxqoesFNKR906mCEuOFvOf6
4M1F2dYqp+SuNjb7YKDUqRDLioKzw0kUMYehI9CL/6CULIJj0l+LrDMiQHWN69IQ4SmV9FR+hXam
/xNHgLOWfnDHvhmtL8/eCRDSu+0VAG+utoIVgYM/44w3DbNT9S1D4K7G5qE5yE5/+f2r5cM+b3p/
D4gFRFuQ7gs5MDmdgyXCJeKguhG0RMp440PqpzrC6KZJBP1CJg8wuo3Wpaae+gkEc64f4jHLuAnO
HfuG5AknSV70y9wtJeXjQmqtqxw+hY+BX5R3wGCa4Vxg1begHakC7NOnbKUQk5PJgTLnSOjOWEUv
DBB5oxkkZ6sEnLCZsWbXeZQFgqaFfNXVS12arxjI5555bk9Iv6Xk1vukc5fHsFvMxcGfdb1/tCIq
RiAuEpk6deRMBQKJay7XwovpRCTkrLqwqFn8yYkCGjn5icTUEHs54WnLlbWv80KpYTUPoIDRW31o
YdZAIqv0EBesFUbVkPGsKV7uo4Lv0htUoit342DpbAC+WAErSsWTwIe8a5xQ1HRBN1UBbFGPP3vr
SFBburLeKzH83OTuP3uU8knBaztxDLJeL8lMeFQta/AayTltWWeKOZds/3dxIfyZVpyA/DKMp5mT
1j71za5kW3x+Sl3uTLLOanRXGzGW3CaCr46ZCS8+1MZkHV+eqV7VhoBgZthScIU5tvgY4t18b+kU
UFu9l8V8pCXhJVo342rMsnZVFYQb7ndTzD+GodWGSQYQDfzWuU8EMiPmFsmUzbqWGS0vauctcUFi
eMnoYPxQlCwG0QaMP+x15cjRWRM0ocrn37qgfoVXckUt+VYf3h6eI8ltnD8rbvo9N0Ogprws0ChU
b17BBNa/zbJB8pAxn6wUaa5TzzClE0B+GkXRPDPKpeH3cP+dNRnV/cvjiDq8fsrm1YWJ68QOkq+B
TNAayA4x9lFQMS05aHYxrPzncdCYAfTxZpurA86HiYkCMgS91kJvcXDl7I8m6lvWaUdPHiqXl/aD
AsbXkeUNOXEbPwqlyFpZpvOikLtDVPYPZVKESWRuPDiomPWLGqwaSIDpFM3Z3UiWDpVg8KoPMlB8
NEijtHz7laKOp1hyVaTV7hAaMDuZdLmWoqJrIF/UBi7rRe9A26nGn0izssd5zFyDqdTbvwyobtE0
0brmD67cYv/JZb1pJWZZUtPY7bsDP4pIGCZuLcGGVaQnnRqqpx89qYBiFrII6tuX4ZQdYWwpSDww
h8O9kBzf80BvxAbmB90yyXin9uOid7MhtPL8JUHyxdEQggwoU3qgYry4ORRFS0TwLJEVKHBb/xvS
WIOnluYWfyfk1UvYgzYgcv40rCJgv429mrETXskW3NENRuEEEfAmYKv4Om2QE0YDvhM5cZtW4nq0
tvd/0ukeRft+CvRe9MXuWBRWsw9NQhoMqyj5jZ5AFmtFVQuj0SKs1tO5BNbKQ3FJy125ws1VXRpc
bfsJ82vOiHaohO3oGueI2b/U94eQcFRsj3X0xrf7E+WrtNv0t7AxVM4GFFq04HzRLkIcuRQKKiqF
CSLZPHQMvLNhYUAl5bf1q01aOHBBQPBFcVvbpGKcGOO19KsKS5Y/UFT/8wiu51JPxmOBGu/gZP3x
ttWLyqqPiQ704x72sX02Njd8UzCfFxlNMr4apW7jw0s5iuAaPqVR6wLpUXMxO8+ZnYkuMbpORs2y
PFlkaWp46SiuKG7l+J8+CrRZ7ehpz70viG75RejdMu/pQVKLTqJAuUH7nX/mgH+4FS9MbtP921jM
aiHjhh5B+SAWS8LWohTyT+E1AV0hPqnghf914Nwqczj+n4U8qiL9f2Y2TloLIkGpMnkyrGtgoSDU
qzoJPrp4hmrnRywD/FvmJFvs3mvyyJ1gmpePavG2x8vt3BsUnoipjE5tnScWhimyudV/rGfgeZnz
8FFGaIWvs6fY/IrdWFumkuUWWYFIhKywI+HO+avOKpnVONMBHdil4YEcka+lPlpH/yArEinBgsoy
mCfahkt2cW4SrqaVn/3pSVD1HpWC5HmI+9YudGy/px/F0g3I61uE4cWt2lIOSu/g4tO5STn8c+sS
F2WA/j2CzqcduQKUcr4mO5XNT1IoAIcli+UF8DSL3XE6ZOuEm50cPlTDWMYDMj1Lza2FTaFRmyi4
aj94/rFhWoxzDt1rnBVnKrZBrFp6yIXv63i46iYzYJsSe2yWNRGkJa6rr1hrishvbUgEfuUNAytK
/i5GgRoDG9LtLZKjQ/US9i95o+ENZtJZW93WLMJr0lJYzg7FrAW9MrgdRvp+bU4S75seVaakqonH
I0EsqMcLYszVf+RAXHTfZRpCbBG1n3mn/IDAN5wOX3UKEYDXwP74fAeP1sKLpDo0Y/dPfe9HkQw9
glocGKzkTu5mTi7j2jN1wByYHuF0C7+CHlMdFa/tPyj1HDK8bWvxNCsDKmR4YLtKYT07EtR0Ut5+
XQBq+8fbUyQ6cmfnsL1MbgX7sSrArG5tbH5FtDwDaexLIgjxudNB6g8YcaYE9XADGpvRKQp2unO6
yENAib5mnbeh3Fb6A5yg7dCdKG7yWM2LNAuzi+GpuRktO/udpJTjj0ywWxkdbZHJl4SKYMWOMA5T
AtgHPVp/o+7qMXD++97/5gs+cOzlSBLNsTD3JyXLC03alWTXCrtkRWpFfhsvyyaKF2FzJUhSc2n4
JjhneCG63or5tK/OTZANRNaKSSFfxZh5l4ehetJew/xiRzkUUUsw4cU5jB2wMb/3HjsZKRnV5IO2
abQCkwurc9Cai3CSc2YELKHqRKKaDtUvTO1VOWWezJkRvm7xggNU+5R64C3yXbA1H8WupzEEHTQo
YIoPBVCsVOSORn/4WMI0LqTDG97rY3L+48mWHdTOX/2S2HaFNS/oeJoCNLY6/sNoWb9sdhNCfpI6
2hvXW9Gbw4F9vmPKRxh2dSm8UJhmssX6AA30O2TmJMfQYB80KSfgzJ8a3v+Eqhy3rPDYeZsM4xaY
8ArDDYnlnxLOx170AiEUuZHdwclVdSuY7uhY9OYirSqxYVGrsTJUv7HPeG1/Wdo8SVpHZdImwV8a
e1HNM7l1i8pQef2fTmaewefRw8i+8UjFjV43VY/wYU/58bIG5DfAkJ/Mqp507ZzEVCd8U7JcX3aL
cdtRHGh+2hRur/WBHnEn9eS4IxejtURSaGiZncj+7joHggAefuFQtoMs0yOBo9BMHW0PZXZSAqGU
UrIk+s/WRW1ff1EYu2hjZ5MGQr7/vbFyIqeKMt3xpmqEiF/3QmtiHsd/tsGuiwuFrojXSurRQdKF
Ff9oscZVmvPsTsUQwSb769IBYrkhd2QHnDLJv9wp7ixRcdmFfbkqKgSPvr0K2/HB4gA/MVW4egIf
+FFDH3G/HMwMCFLUGCkk1g8bYIcXQoySkq7NOIqEy5N4WX6vWbyq4Zj1J9IffKfjZEyYFgKW3iOG
4U3VL8CROaL1aopzv4ovVdHaRM/8KwA5hEJMH7GO+WKG4ytfOJ8yz9lwWfL/hGttQ7bVj/JmiAZ+
dN+2AUgkxc4W5v+NKrvbCbV6ESmitRJbEsBYcAXdPwuXI0FpDif1utVV+Lriv1yjOvMEAWspzAhh
WiSezXwBakS0J03b8xPaeXltnkORfFawi8pRP+Vr/0xmuiABK0AGovq7alyavB1is/5+Xl4gVJzP
pZzaywVRcBdHhZRTOvqLT/NaKVksLIMBOALCamXqkYjE4DEAqGtVuB+r6IEKDKbkOxdDdql7+nwm
IB//HlOYek3hINgcYgtx8s/RFHyB4a7mKHw7p7jgRI3HRJFqlQ3BvdpWcyfM1n4RceRGu77KxIL6
alBZ6DxiN7pktvH0YmfILXzTx1oeGN5/WtRDG6GQypVBgZAYEG3tIVTqOsUfpH0QkpS4cTLwpnBA
siu0Kt+Bvuhh5xOmbwhRMl45rdV5c9zyVMK5n4xRbaSrqEzyut1PgWSDwdpoFlUgA9aJEW4qVFcB
JQSGQa/Uz0G3eHEEFBWGs+bH/1/nQVgdZ70pce5rZiWGSUz8zYFpV5Bcue0K8Gik0R4c4yzvc43O
FgjXp0vK8Yo3rf8HJcH+YXsBS8DsTApjODQWb8OoupoGlDg9k/BS71pIH05ZGuhCsjTOHQS9ZS/J
1zDiu8NTblIWb++dKy43X1senwg7RSN0gL0R6aWnRW1dUAPh1ppw5JVL+5nIweBRrlK1th6EHcEH
xkOC/CTzh28X5NsfGnFEAODYgnpvYUna2sKiJjCbpl5Wv+ek62gytdEDI1Kya1pfW/D0RJi64UKs
pnW+Jmlq7dNlEdGOCmwHEJUZYUAm/cXMttVevs2nY5bpZPBJBveYFmhKQQVMvEdwqep4ww5Fzt87
x9H4ypfmidCpo5aSV3ZF2jRYJBnAzwAjU6ceOIrwcco4QTEwi76+2OqN20dyzR6WYqrfrLhjKcs5
L6qO1oXLfdQ/UTdFzqxrYlss086VDZ8A3KFzFBDyCQWt5ipdkOCG/w7F6UcHRjoD/Z2Ufyv4A1wP
pnMvZTwXXWQ3y8g1fCvH9M8tUt1voQbmmkoIrsJutXj6kB9QpHszhhH2TcfamjwbTavrhnTU/xSu
942Kq3q6m3qhZ9AdsfV9QTKmRa1jAdD5a/mB5ik3VQGTnU4SdC47S6iWwZU/RM8L6mOGX8jxKH1B
AUUC+18XEhHe8VvWYIyY2ptRaeJHv96n9UCm50e2mVGa/OZLmcqszr/Mon/KUVQ39JGuNUdIE1j4
HUgFiFcjGDRv9a77GjyLG5n6J7L1DlWAuzjaMb3wVZ16y1nepGN8/C+GYGo1a77DzfitL29CCIG4
CjdoBczVTjcEL9nd/yFpbh+/cjlitLZApM2hJHb9RKMHCEfRMyWKrn6VduPbFUReSb1bgS5mlchb
qyeviGvF0Eld9XHt5aRv3pipPWfYPG0oQYBEbM2/4QhGq2ezdb7feBo6MdfnzRNhopIBjbVc73Th
9OTGYxWAGhYw/HhwfWhYpsfl8n2Gerw0D5SWURP1GdLT3D56k4UW3aELxvi8jYMck+1QDcYAZM0/
gLZrf8ArXNX7j+h5cDOmRZYK90J8Ob8rKi25BJdfWD531FF0cQg/Mx0vOvk50TJ1m1fa7w0B6hke
WuNhlL880Lxv3HKaYPaJVCe11rsykhaBmqKf1CHIK5R+JI41zeUrHQ/YlgezQvhkMiHllF23yR17
AWPEMxcfMvwxPUlYPOlvKxVlbFNUIwK10oPChp7a+QbwxpiRqNC1Qx+9u1aW9EOyH+aU7MdyFFEt
yp/mNLyPTwc+l/UQnVEKcMPgVa4QUbYI3ekh3fOYmCG1aidO/0pyZsbi1NLvwW71GhLtG7eDO5Bu
HoEoI/745ciYzz+dyw2sQ3ViHd9fxJD+noNwoHjWOtHyKvDkOC925DMCMfl7UXrOyhPD8gkvjje8
Hh6GZfzMSrIdAf11r/JpWxD0wUvyWc1lEB2VO7JT33PwTBlco0MxM2lzeePPp6fo8/hlfpPeL2ci
471piLM/k+XqG4OpBaPvh3eXnW9/pCH3oA6JTtfPnfZccQTGpDJ9l4et2uNgc9IniDmIhrNUSwh1
R+hJE1mwE2JZToISNOgZSKEGwMzDoz7Iwtcq+n+nVoS67hmRg2qVlgXlGUKb+7kGc612o6CjDQRs
se5B+qfMOHwTRDyn4R9wBRQ/XgLkfqIX300B671qHzGK0bZCeFMlK/BnE5tDgMPqqkrWgv5xPRCp
wxQ6DgU8Ui0aV/yIskQp/Gj+1G4y/uDPBS7/044+NBwGlpjMyV857djaamz/qy/iYBRxStetpcma
aRmJMog0iCbNNfFLc7ESAPaD48yCNnM3rNKWpk2QmAV6KZkVK3K57YDOx/EhV0+Ron//FMpaFaOv
IDXmGwncE8RmYbAEv6qkhtvv4lSsy4tx3s35AxTErXv+BO3uIeguQuAfWeTWra4iLnRJhnFx4IbP
vSUjQCV9IZiwRNPbxYcGQcvIaAEJkXeWUrOBvA7uW8McWc2CySEuag5iB8ZxNX1nbDHQoQSVXGy2
CLt3cQMc7hQoBNnuZaLl/YJsXGYUES2ZhzYz0gHMmzP5JlXw1KaGHW0wxPjt2Z7v6JVe4OHPxPFM
KcRU0MXv+FMwl382Oxb2I7IIyheYkwxgM/3XRmgrYs+JzhO9TnQA0ottrnx/nJC16MAaOI1bK73u
NxjGp2uD08EoNNnX7F6atXrdYFOghcz42S1/2IdLJAEcT8G60wtqcNcyxSqJnTqoNIH+sgJi1ONa
h+4yTJmvZ5wpaX1mAv+yjf0Z20O+ZdCNeTN+mMex9td9VGah4wz2EV2WoRMMIDalzZe43oHeGl6U
OHVDhg/T+kASuhGw9Rkxgp4y7QdF76J+ROQUn2MYmeCNcf50q+67Cyz5cPjSrafqLZREpjGr37if
CDjxm1lvpjb53xJ9An1/Zyc8IIl1p8mmy0Ui4/l5+veIpIl7dD8UvXw/BjJSVaSsJcfFgGUaaqVy
BKv27pJ2xp2/CSV9leBrTwkS7UtrLcuY/YwNNJVptWKw7R2/xPPSOM3SPtIgD21n8veU2MgBH54U
EdLRjK3QeOTMTutFca5CVSjHsayTkKMHQXfikx3lwAZ7VayYEGrZCr7QKt1QToogYCkNaKD4SUOV
eqfoqTw0Xg9ECtyyUKP4RmlUeKGHw7XnbiRvKyutJxVz7+TXYdbChsCwl+xa5yi9DILmG8YbFhI5
1hBz/otGsIqS/QFf9b6qim7vmPovbGCr+CoASbuNEjPU8qaikq21FkGp+mNiu3CSMbpxbS01YEFV
00iefyKlv/whl+g44Cy5e0FZgMpjBPrMgJDqY1Czf5CEQsVSx5GEhPeIuP8dn0ECODf1NYr3VV8j
w+K7KV5M0q6RTDlTw8wyw72nhpx2RYq0wS+7JTxdlvNfqRUbGc+TvLL+b4HxwwiFISxxMcchrYwP
1wb3c+fMF7d1TA4gxAqT5AMtZvbAUgwCjI/cWTiMquv4w/j2vGlu9+IelfJM8JCU01B3G9Q5ARCu
06R3kLM8v3VUc4tf7NxhBTgCyV4XEQUSuM3B8+CUghGMaVnNXXNoNZ8v6MmXYXcTM+kW+LH2PERr
DfgBg42zJ/j7Xh2Q7rsU7wM8+KGClCSfAq2mfD3ggS5Vg7ST5AbvHQ2GimnPNEaU+nQvzWeoBZTh
QUYzRXKzEjoj4RId++G2VbUL3jL1DrkKIsHrNwWaIL1R0kacurAqug7C3dSsghLogy1cLZ0WntV+
rdJVgnx0XnoOJPHneSocH3DJYioY98jc+QBXA8ZFyivhUna2G7hhG3YGv1OzNjprnf04jFABMn4P
EFNM//SbK3US9lgQhM8KO1/1zcRC1xgWRgpgcI0prNsYk9mUCtpFxR5BYyamV7QvigeybO4vcsNC
vP77zr0lbqJiAAM9N+7FpNKxI6eUHkJb0zzWOcxUftreF9d3WW4ivBkEXWsvryXfjanoOmAVdop9
Lyq1UHbUL+DmGN2Uelqv/xlJ5HoBzIb3fTaDwaPGt5iXDu50xqs04OlFmaHT48Zkc7cM/IZNf8hr
5aOPOjLdTGuOMwDvzjWsiM3g8sznMWPuP0C2KmrYbBC3XuJJ/CliZmnDmZvUD80FIvrG2iY2PpLm
Bim9zBcfM3kaw4FW79p+1ACp29m/+TClenf4vdAR6t2bbeeYxZrIJhzAA3MsY47Y/b2YSEMU7J9L
JNnjPyAohSqVsY3C2BBI8kHVqgegmGJfanuiRbG+xEeSupPWPzm0v/hBlBIMV/1/ztsTD/TA0FGk
LhGKXxMSjjk4XerYClIWPrMxPTRSN+5KZmwzU7BRvIaCu8rMzbv9Q108/I1J9711D6oO7um1R/XE
Re3E0EDU+T65wr+hOF/A1sKLigCqgPiwKm3/9z7EOfhXnG/i9SIyLKfdJyHrqeRtGAkb9ZX/KuuB
O9kh0Wl5JIwSXj0A4cfLcav6ThK4hNSsZDNbU3s2kdKkp+YZPxI+nlxKkFLQJCdETohusxEB73Z8
FmURjhC4fAxQke6o++0DmorJfj28nKAq2+yIyPlwhmxsVwPF8yvhEGG3Oe7l7oovW2Fr70pXodOw
tqYPW3Ub2xtkqMwOKLVOGYWya/afmu2ge3Ylw4NfAFKufewPg33Gr8XgNO5e78KUSnE7kGdpJnG3
gLEgfv5HvurS184yMM2ffLpVZrNb0+LaJ8AH4/ZpQHc1wDwg6DJ7X+RNBcbA6IGeanPsJ5eVcddR
3jWVoKcQfdwsB1/9FBjFvorSB52d8S9aPPbo9jz9ru3jsRH3c7YMfPf4ZTbdSDpWgTpzDWbRbCuk
7hb8s6O/7A8kOgMwUtYeG40n1aqT+iq7IOFUQnq8WvkE7bNqHfjakRqu14NR/w+0u8hfkLKmKb+i
QEZu9waalzxcc5XT1q6aaur8jYlkcv4HReVRzANJagCNLYyDq7yegvDaiLuL78CkjW7AaG/H9GuC
uEOYPAghDE+MHNC68UhBgHGPT5rjKalnUIMWz7Wb/IwZcfj0mLMaYGL2UjjeMWAOGYRH2mLL1lba
1srRzbJFfVwqiZfPVmB1LvJXIbt1E16zjXsNeWtEOpvVc59NCCY7F3LIfthcbpvBCeHuSHOoI/2W
PkqUeEogRz11XlmbrIUrmX6byQ1oJiJQ4TvtSKOmVEjVxV8p51T+nhBtHRIjTHyHvwx9fHwWpzAw
uZbMDYGGZa0xhL1CTmDVHFq5kW+E03VUiXCSf9E8lJmuUMbo+d5NjiIxn+knMd6aOwXgk5l7Hn1Z
MqA8/l544vMcx6jx+uKZXN8+kLsDCFCjCUsFm//ZjJ68T/oLsUY6TwZ6wiRmVam+U/XEbOp0xxaf
DNG+z7rkotsuKXw1309OEOG8fDAHTZHUDXWZJF7WQXY2gXDYP5VAXYRalF5KujCUokH60kXbbUWU
hU2eBHKNhRuaOzo7JJZ1soCLP0W9qzkYEacyFkoH9K8HbC+fQp2E8u67lDcQFhAAQyje2ay69/ZQ
8kWPlFEEnz7tuOxd0IEG6DcGk6Uw3cesam5d0sxUag+t71TeVfvUc/G0RSLkiiDB8YdgWD21lzGD
DlgzWyUIvPTerbDvcMvIweFLQryD0qPvCTH579uhRzi2Uz9iKraYbH4q6YkjPEYaaeW2RxylqCFS
o7GXFaeymEhgjJzO+385F9AFg+0PclY3lpnEtG1Q8b25d/0PUYaWCEPDMoRcYVaK9HFHTDR8y7Y9
H3iMzCxh81PTxYVHdcaVdCKzZ1YJTZvmQQBj6N2GOs7sUpen3LTqV63SLsFwrAtmM0xc+SSxiaDy
UTa7c+lZ4xdAycsep3goD6tqm0y2JsgoKw295y0WSmwJoIrZOZ2Eswihw0G9PfrUEEuTcgXPuu+D
sEbydXoDGRXcQn+8igerYYGgKDQ4Tk//FyhL5KDN/6uJ1ZLSsQ9TNfab6q+5+uFbzwAgM2M1PrSR
A6VHDVKnNwgRAbGeL7urPWANTSDIYzwPSKXlhh+A+HoVIkUdtLtf+F/Q8L2iaZdS6RPgPPwWQJ2i
62oaHeehqkeDXUgiGdI4C/dn7sUp4tO07RUzu6CYnjIKiQf0SDl/JaiLLlJmafQSDZwD5P49p6o2
qJa3cmb9VVipEL+8Jy0U/aw2nKT94qtHh8EKSf0RarwRyVqsB3loS4a4A+gQOGd/Hlho9uDnCzFa
MtIiZ9PhGgrJEVmDY5b73gf/nvmsLLgY03WgmC4Y0ri8uPPe/fEPYiLCeWg4NbD0ZkcI9ozbrd4k
nJD60/tXdwXVZEuMZVCATCZW42Ld1M18dZDnxC3O0EyiFuqjTVO3yc8UmuDi7Xa/uvfo7aFtSSdU
oPSRloX9vVH7CaNNAlg5Y42VEnZt/3OPdk4PsdLkMyq5MrnTcPyFeKfojfCNhCVwBPYcUhDbKILi
4QkdSYPcbZSa++PPfdBr/zlMOrdoNOGgQu09kTFoI2xcSaxWMrM1URZBe6lQK6Q3/TBKDunVJKZs
c1JjH6aUtQbwBxgi2b0r/K9bbJMnGW5XAXF4lx/r6IpQDKF9a1WLl9gLj7TfIk1fmfe/cP5V+uAH
GOkeeAqjFFLYX7q/NKMoZPxK25OS7mYbkJgFnmWGJcQQy8OFdkEtGKKG8FOYqhBkMfg7N1YLWSZF
kZIPnR4tm/tM1MKFaVilw0mh45BJXOpPfEsWqoEpDJw/FlhFyUZ8UrJ95rcvnntF+okaZARF3YOZ
bLhlEoKQIm84k/EE2nKzd6hphNWdW+WACVQoAcgW10jC9FCY9C+ayKr6M/9bAEzfZwG7S7a2K2vm
6Mbbqe8kSP3aDzTvTD5oE2cboXcWq/2osZYd5CuwaJ3KvK1717lCpwtvS1Rr+Vph5CmfuYAK33kw
iJCF/l+uNRH8toGB6/PCsyFA4hNN7kwbXw2E5r4pJ91DK/kqA4rYI8uahNTk18+WaBSSD5POWa6L
DPIJFhvk0yB7P0IKXCtA3jEPd3c8OFUtexaxOuxGzdFipvp7BRYAENGw96F3Zjo3IKK05U+d/4vm
o6wKxtbo93Hp+QPubPsr8wZuL7ygMZGg2OvnaGm+4B6LDHwA53uO4C1LGF6JgnuWIjgBSPS3CbZo
Qg4fEvzETidSt2GjpaXLjA1Et/7RNgn+7nrBFOZqpVbUf3mjlNQsqNktP4fVEtLGutaGUlK2oiL4
CvnWKS4A6c/MV+phvETNQ9JjzwTNz5KFHmRuT8mIiZg27H10fo66nj5yURppXKHR31+Wh5uF1VHT
JhJXo2l1sMWioSz90dNur6QIF327d9yssoY5YRle2A+Xzx+hqne+mybz0aenKzmPOj4BEcI4clrJ
/MElGug4CMvD8mxsxMeUqASDK4Z6VgLGR0E4Ir2nKwedHUVcWn+Spplm5sboSlwI0BhIcQ0xzrfv
pohtOqr2pUKHVUhwVSCjaKBeuQ08M6zunrjeg5Tic5W0C/UHXG/xQalTg5AG+GDCCCo0hj6wiJ0Z
FuFX6HoMfvZIwO7i26767cbnixXWk6/aRxWGNCrY9+Lur/C17FVqsiOLXKIbVyqDHujiKqk/oKu9
XIwM/zI5KKSMEAN7cSa+v6re2FEq1bxUDyJ3SG/oEAzc9HAunQQn53OjpOQlPUQioB8Z8wgS6IdC
bWAA5vN3lTuNXoPrf9WblCBN1fqEACd3ksbGe2uocDT5o5QWUVBaL5iuKyTpgFVdIvbWeQtUkLwS
0EYWawyGW7DeNG6e/mwp0dg+oBK2nby1Xa+0WnQT+JZLP2Y1em2Vy2KqRB0b4v9r6Wgu+og9rOOw
aIpSomMfJKxcRrhLe5MqGvRXvHBkzI51qE1NRYAbOkLupIJZ/W0p4rlYS1dx2FwCyEzGJfva8JAM
TudHy8tGUaOf97GAAL7PWOIDT5xtpRSYZgxP5cF089GfxPGsX5vHKnSgvzRdkbBMcyf0vMaZYyUh
I+uM4tUIHPD+w/t0rNvs6btNIBIyeRz3L45mU5qWnmyxCoyam3DGcyS70tq4r/FmhLWJL27QvZnX
Kio8jbVXrJjSzcBKKRUEePrClqpsaSYciTAXBRphyR1H66dd0V8QIrZhJMwzQeMX7Re+6t1DUqv6
rn+VGqjLVKJzpU8Vb7IWECkDj4JUehwMya/5GgBidmuo4/wWRCO+UoIICqGFG2P+6OhcmeGl46K1
2FoRMPrGZZmaX5+rtt2Aca8PQLspIT4HbNOlW8UrYRqWJyjAlZCIX78IkpV8P+uNcaC8bZi57jpz
LJ4bmercoE7pyNZBG3hdJGiWZHc94m49t8j0CVIzyLjSWyWO5z+2GTrM92y5n97zIlj7K8ah73sO
3S74lj2ow974IteNJQ05Q8IGCTxXHRKJ48yF1BNwbZjpaqt12CTwoBYxFL3jCE6XXQypotaxej2D
FGUfvFjcByHwOllp9M5hbiQOYQRtimOoYMgoJZJMEc6KxOWWMEyLdYkVZnqPh2Fy5/taXoQ9GenR
Lete+jedm61yTfeFWEy463DFr/TYRH5zyl4DBmIgNqjsE8j2fXIbH+ASggRcVQfp5VjeIX4qRPw0
xKwvduBt63ug24rtyOXjI8JKBr+Dc+soXpfVB8BWTf+SJ3Pq6LOV1K2DuPXx6vZHkF8mCsjtnYKR
IKnfOru0SIjSbCCDcaFtsEWdqjGl1XZkeEhgOX/cogN709zsemTjjhW0e+NQha/6LDuxnIP2X6vs
KUOEli/96W3Y6J5oAGHkI1gpLhQ4hJbha666/quQg5yntV9xmQVK2TXvkL4sEfvxEFi2WGp0GFKJ
hPxqgbCiHbwmDBLVjRQzggw95yrV+gLM6I5RVYr4O0olWoyvv6br+B1A6DW/nw2vkqrpjvA90sLs
VrV8pXp4Vjnv+g7gvaq5yp/rdcfxULKEPw+y9hH0WpUg7Oz6uQbaD+AMmbwdMJLT/i4bCuootk2L
Zrd5tiWH3W5ayPhAiH4mAmEmBlkq/7UE5LCqAuUhufluRHQrTZNPWiWddQAEYmCwSU0mDTpHaXCp
NbSc8Lb4cYoBx1HVpJdMZ+PtNqZiDBz11z5OCTunxUl0vniqeeFwr33hrg2jwGIPF5jzUXRepxm7
M97jMCMJFpiOsSwkwdta556E6zAWItIQApNtXshLNeo4iTZyrRARZ64K8bKOElKy+0qIxBsxJwnL
fFVYkoLj8egZR8UdJYXNy6QEpAwIg5h9nu+H6RaLVMfec/NGItT6jLm4AaOdPVWHY9sHipZwjrKd
xS4gP3MADGzQ0MMWDsg9XiJuzqRKEq/BR6Up1EKeGjU5bbg7KhVfF9y4KqNQBIp6Fh/C4rcJOo6n
CRAfR5A49EYfj9re2xzFHp96kIfFUWGCatj7f8+wuTxTQtCtgI7on+dqxsnzNcVqM4ggC/f/EvJQ
mw2Ig5qKtFbf5H8yUbXDnvNxMBrKfrPRxndqgqUBSHSzYpuUfxj07UGjAWVlqaCEm+v8mSnaR1XK
9dJq4gQIS58G43pRoioW1FuwGf+FMB8HcECBM5tJCB5GVZgkR3lmmXAIUTTFyPTl39/iHguVtNfy
K7Slja4KGOj/HKlDnVMxeyUr2z7biCSDb3yAlUJ1P4eqxoZn82Fs+EqgaCCmmzkf5UVN3dJWjCwK
As4M6APmbXQAMhdrfiPT2xtcL7vyoA01wFTTn9Ga0cb006oEnTxr1CxGVYTMICO9zXEZu5m0XF7s
kJOaHusOkJ/H/SocLlybWdS9g0aGLd3sRuGT10CT/97Yk20RZphiU+eG944pTQSvd79VdayKwhKY
MukXLwDM65Af1t1BcJlbFYpuXKQmbiRLya0k7GNBHZxVZ8gty0DN6pRPaZvZhIA6PHOycn1zQapp
UQgSpviqrsAJE0JCJ65uxZJqPKdb3XPTqJNFu/TmP1eSJfbVP07Igyn5wnVIRj0Q5if57iMti5rx
NItqaSFMKw+o0BCrefUD+xiwulnDzPXnN09J+RDdGaUEC1nZeXOutqTQb6W3lhMRQ+feZeZBRPHw
rVZQVjC0w/79fevtRk/BAadA1ZBcXQNpARj/HEP9H6F6BT8S70oGdWqYLCAL326ulPPh/nhbpjgE
NAJ8uKdKRyRevr6KGn02URC7e4j29LQQa6TayFELJfDmEPzWvxGzRBZwxHJrkouuMhdcNVwDpl3q
ERplugbpL0bXF3RLJ32VqkKb6NSGtmmjvP4Et5ix6xIm62B3CKFEmA3oI0u1SzADdVovPz12veZl
w+4nJ+5BTb/+Ojepvhio7PssYboGIqcfkC0U472U5S1NHivSDKt9h27YFzbXlCmL29qVdU7FuXz8
pz13dutKDh58Powy4LRd6yjd4MWrbVaZnTX40sTYXdM0DSPIj2PApRdNMjc/9fCmIuBwuBoKrwl0
igtZ/vearQFLEciguMBCFsmEZLH+SxTP2kj5gXK4o7omse2ajqIFV3VXp/OtBCpZRVQa7gMMEuiH
SW0r8JPBa7ZSa4UlcO2oLnuk2jcMM9bG1ZkBNSYA5k2tv/Z+BKdZxSuq4j6rCPBXu+f7aaUWmgZu
gpj1HgjD2WwXUB2u1ablbnPgoSFYFGh29hLU1Ir8UUBpS0qzRl9xbugOP4HIflh5UWdNK0QpeGMA
fRTKhwZS/mmiHyRjZY/XS4tyuhyMCHHX8h39SG1VIBfSTBh3FKZ6eEcBE6yqRQAti3q+v4zruMLu
bOT6/EHEhJPxmpe6V6+RWNe1ijRzS9SHevu6c94zua8oa1yRS1X3feXeDvCb0T3mSFGThcY0TUoE
7euR+HiOlsXpYzf7m5i97SzAy/dGIQFZSXPvFy8DgxQNgjlMScjFWpKPUEhV3EiaFv/W7woTuO3x
mjeYDezZCtEDS0K65TQGIC19kDCep0Lh7E/KheMZBjfz7+iwT/+/yPss2F+jhDHvF5mdqqmcpwpq
6TqVnRRtcB9Th2WaGo8QG2smCnXjV1rqQq98I/01gPO3NHsWwNsubTyJmOXe4IlqD/g+lgCaY1w3
ydXksS1Ac9GkJH6s/K12Hi5mBL9z7EpcSP05XP2nIiW+QVslG4vYJ2Me2cQl+KBWLtP6xXhXpjG9
2Udw96/8j8Qf6lMvj0ZulPbIBh4b0iVw068IwS9FExyNLkAONABSeJFtxFsyKmF9N5JokhBADNg6
bM2QejVPWQo8t3YGPmqpWgFopHl130owI0YrVUhrcKion/4wfSU5fuvcHYxKXjcDsRkVD7o9y54E
f68nYAhsS3LBSpWngMMHR+kgFPEeJ4NWZa3A9QKT3f/nEa/D/Pmtn5PF3MTYJIOIxXOV6/vrkaz8
CE8IyUW6Etn+ZFf+zoM6NsEQg+zC6bNscIbkQqF4UtdF4OuMeNQuvCKLnXzyZ6yDmtHuANX6yt12
wNp+5viQjzluyvTpRhT8xILHW/v9jDPMfS34sbk+LCwLT8AuqBGRYk3KnTS2TE8jzKRSVp1D0tFl
5xx2762g2jiDZOJHYpMEzVDqsu//VO7r9E6cfMPsixKLugtc5hVxfcQ9hIrIRdkoch2R71zj2IJa
dos5rKnh7Wq1ZTTGQ5ynpKhs2SevgBprhc8GIxXUH0WTxcaCArWlGHTPWpVRKGn4mqrUXmQy7TR4
IB0O+sjm6L0F/xOZcO4DEhHpdRMv2fVUW98t7yG8w4gD5UpQ7Jyp6/pPdKBTDKKHxl8Wus2+MjH8
bvZ38tciOHY7UoJ8tV5XQvWd0iah1UD1qVfllXq8JbJW+dsu2cNqjpPcLmuPxHcRkmsf9cNqSG3b
OwGq4qId7JDQ0LuXHU6GE/Jl1epludj/yRMXQoax5UolhSkU+H2KMwUsZKFt74ftSmt2l+mvw0pX
T27NAiNCS5HS42Ylr/uKQM4QyRx6RdJ/Qh9IKo5PXEjeO8FwCtK3ZPzcdSuKZgRQOyp10dpAr7N6
nSW9JbfQfON5EdvlvakJPdVE8yQmtYo+UEMpG2A7z2ECgbEZDuLR30GgcJ7HaxpwyFR5X/6Exb9e
8kReDTrD3VQeXA3NKashtu4jOiR4RHZkkXNs0LVk/AXof6+8T2RsD6+6Lwa9TgAXzxAO4R35Bbez
QoBkVhcgvL152rW6urIyqj9oMJVcI4SfWUuuQsKusrBT2Y4VKO7+cu8N+R3f3ANBZiR9B4LP0DOr
iiYW58C1wMhZwRNGjmh+mgiZaRumQH/etPZ2xxR1sgNFsDgUNiKqaYSDAUJBLYHFEfxuWcVzwJXb
UBDEwXahck6ZVjPG2S9uxnqYz1PoWlvCu3fA1EUtFU8x0uVn8DKmK9K5qeVmOzsrsJi6yIWvcs1Q
4SW6r1hkkEvSOHv38yvKEwIighvSnAIJa5bUv6Sj7/+hJrBOFuOjH1N0z9kb1Z/r2uJXiYl/e429
Zf3BD5Yboa5Irf64pTUYsVoKDOu8rCq6Y2AlkgtnyXhEKjrI8SdtHIAY7IXlyhuhrzC6XXut3RTR
VVwJWccjZNarMqHi0c7RtxDyWSgYkoyZ0NoZmrkClaoGnvt5u5c4yF2B1gYduLjK4X9FxfWe+N3v
enFQAZTAwyOcj42jQKqGvbPsig6WA67j7ZJU+HFy/7lVX5V/K9I5iOXLju7rvVwBkDsPB8hMpSnc
y7aC+RdBYsN4ibTQcVZJAFY76s24btvhdK9DhcVpUEjIiMfFO25ldJthaqeuqGK2osfmRzDg2MyU
LzYZTHffoVH9I/dIymr5VgkrzioxUtqYi2YScG2G4CMRFr0qEYngZMLHHnEPKplZ2WjSau+b/iWq
qc4wKD7CjnZXY8BoIw22BCwoj33+GILmTwy7N2iXFcfWu2wfkqT9hzUPMTXGxtc8DOv1WNO0411t
pKp+Yhz61PDnC0gjoabEueeroSF4AsFRMG5pgAFxeF3KvE0jL1xVPVmYIRBWPbp97+ZWdhBkGLh3
yhiAqwk63DnasoVaPdu2Dl1xBQG6J0Ns2d7Gn1cwsIfUKm+yzT8vxbLLSGgjR/Ri+qzAllmdjb+A
WMTB1qYzBN3cVWxR/OwyVH0Nr3nGJzfcw1Kl573V2bLJ9RLMT9OTcuPnC2uKW5fargB/9xVmixdt
gDSnZ9Ij567gGizAIU3FbnulYnwtqRBLB6ZxuygYRdIiEVGV9VKTuj85T52wonNbBwtzt4XzVVOe
LEvO02CTbqiFcksGZcBpSkhzRMwYxcuGy9BOwUDa4bZPDCN9N0MNWJAQWMXdVnfjbrtcyAnNXEvc
+TpJWc2mC5KSnQeZuhtP6I2UFcDACRcjmpAzycPmJrhWtCCtNtilG0Ppu4tjO1Fus7jYWIJta1s/
d1YqUSVuYeeR+ze6CA+x9tgkZ6NZKPBSfEUZPnWduEgcHUYMMh3PRYb4AWYzy+ZrEpe5zEo5QgEH
mjzYIBsSdZRKjKicZ4saVizU48YUmNhbjzIhT+5qVgQ6bp/q4Hio+tOLM8eO8qJyX9t4JZ9WGXrm
fwVFPZ43YCRFTxqa7GHlbCyHyzegP7bp6lGnvN547czI9I/tb6GYvpSaYN5odgP8WYoT5dZI8erk
Mu3FiqejiCqexDfE4STwJaLwPiCfHWMERmyXu/73CeEbn2v/MQq+YNkNdEy9qswGh0vJQIi3F+IQ
d1Xjrin0PTalgv+93HYSAIzxq0JT1wcaR1sBvti8BcfPiiv7NbX7ge+kIGIXSj9Cs9YRZORuJ+0z
1Rdqw4/4sfPVbgHDp4hRfPsQ5E0xHrktRfWo4p6+1uHGOd1wF54ZS6w2gm6lTTnBKE7MRHlBWh+x
ABubcIq5fSSm8+nbg68mXWAt4fGdV7YrQ/B6hf/Qi5KdgSeWzrFuihft0s5KXl/jqsrdbKo6xig5
9thT6I5MNS1rcPPc/sP5mLdYA2R8xmxw4ajNFmAsfxKm7Eh2LvQRKeJ6GKQyjFqCTp0b7NGr+jhj
iaeevsfs7X3OYd7bevsFhq//w+afbMhGBlER2wJ4Y0FDKYKKm0L2q2Ymd0aJwf3qvr24Qw7GDmBZ
GHXR4DYe/oaL8/QUK3REfp91P+N197wqsyUXV7+2vdzA4o8nyjOmhCI8Ekf8HUDZElJ+vhtTs1mM
tGIFu86S400Jg6HZh1sR6rBgtX9PSUObDMO+0TjlXb06GJTmdmpGRLFkLgoHSD9505dWQNRk34WO
i4/uCytidRrndUy+WTiX0pUoGL27jIBh5GTNs+KJf5JUkaMwppxjWoHj4Sg4H5eWA33xuMyyTMut
7M5ruJ9Z9T+jut9myDiRdJ1BZdpzPjJUuQVLFO+jF3eLApCMD9xSH1DLm0wCNNiNRQJDhLkD3Ijn
Y9vaoszajb4+apeHINLrLOTYBAQfyrE9EDpFWu3k0SK3xm+Fynyw235k0hj1JrYuB+QUvgN+RSjC
Z8jydDlAP8QHtNfIDX73knF40Q96lYqGJcyZIWCV3nYHGAaExq9YtuDukfpL5N+Tg0ue/bEdWTlY
A/fsU01FZM85BXcRrtz7mYSaDfeWTMC14dQdakRdqeZom5XZe1psGkt+xm0ya5k5rm4viPCAKJGO
RHl2ay5/SFR3tZPBGi8jkw88aN9WgNBqpuUP4e8cIat/dXkB/bhJqeZQSY9JxmA4x6xH89gfhfYN
ffyLJ+iCeaD4HKNIVTgGoSl2WtJd1MjXOGzbclnBvDHfKppz+mBwUpytM7Qzn1XggltCVlZJEPWZ
BZprXwNSA66LU2KsC8FOojozDkRtgl+UXSwH4c3WVYl3+tkwJVro+BWadEW9+k7Q0IPfydERZAeO
t2nG2FEI98Zc7GflMwd6hOJ7XeRp3NA1dz2vPeuzENDx4V0XgnaVlrZtXoZbQu/4nZCmYti6fgx7
tS2ge02HYqNeuHZ/lOFkdVpyYHJGHkfM9ZjSzJS0V3BKvBGgZHxsqLm5ew2j6OuqvT+PsoUvYM2B
B48+kJwos3krgTtmt3gFcmp+74+McoOVXWa5UoTymdbxgfr41alYWzp0nzvPMamdsSPiFdh893ga
wKQliWnHUeTmNPUalFNFdQjuob4JxgwcYibIEYnCYt8Sised5BzYxDiyaiB8UERjtyFBk3N0PIyB
Oc27rl7AB/bS0skoouQ0pogxIwyVYcfXxlLVQgwUC9UE9L62DF3Wx5F9SG+Ad5wyYWh5I4H646K2
OJb+6tT4It+DWzyGaawjrFOCvTBedH9rq4a0NZSuJ65oKvhbjIDYRwN/B9wSR0cYz6CP76i4urjf
BCFhydjLnT1THZNVirmCGDukTJ3Kz02RHQV5mm9XtGHP4Nld1fht4eUHBgriRRRVrzS0x6qhnzqZ
WvCbXM/iLcAd9kkJWUqvtMqDXeRMXrQudO3bYhum+qWhxHAgY3AhT2FUW/5wlcuBfvb5expGEq+t
b4xjW+vAwf25WbT8iBc0Chvpp+9R1SYnN2myugOELzwVGMbw3jVfTzw7RB4sl9SriXAXhtnQ7a6E
6RYzIAAtoagAq57QKAQKvvh5GNQMBvxi/JvWVGZQmgg+knafWr5Lst2Xsuk4Pu66nOaPPKXiLCG7
bdJ7QdQbABLpVjST/4+4vig2jfKFuq5tz4mvYL8P45exW1PFMRxMoYzejEEFyIyrnKUfedp75dFL
6SAjNZ3yj71atJKTQD3UWpzAyNSOXAIFuSu31AOZyIMbqmH7rfSoVMrYuiwMDaYNIBSM7SUmMvLz
GPy+pFmTYNlfaPVrQ8o/8DGaWddo88g2DFJJjLvOhjfOqfL/mYPse5VpTuh+nc4BA7Ruh/jHc4rt
q25ynraOjeSP1EIb0mdltv2tEGD7e16PYvK8MPcL0s9P5RHpQwdX3alv8r3rFYfeWvSdXQt1m31N
WiQdjd3g4uuLO/S7L00t4btmWPGqElZTo6/u89cuh2wzZ9hw0w0zIWdFA3OXNrslfJyhF4CP0xt9
YvRfb9Ok1AQ82ptBfMCwvRgmBD6uyQRRwfiXC8FxLHkAQXTpeSXHuA/zAs/LQnm7BllovghZ/wUT
O987n1NJnqR+JA2lvxjBEiXFDDzTWdpcbG7QbmWfVVsTudBaMbCJRX3TAnILMYLXQLi8EP4e+4cW
xbOBL3PHd70b4B3+6zKoGjoWsliYRHsC+AGRvf6LCer7atIbZ1xc8t4RbpIoQRmRakC22BDwj/ZY
ams/pCktHUbx+RwfCpyhtBJJ2u4UQJEVZuJWE1w0hhj5r9XLqOg5UDecpnHF3QpFc/3qDrOZAbYy
EalZdaZq3zMWM76gJ7kTntbKpKHWyayG9qbfM+2kdddzF9TjoaPr5DLTPiXZ938dBgxDDyVOLU7m
RnjrHBGAcjElN2kpJ4TcouizwCAhnjAuUFU+vJoQcV/LGpcdTR9gCBS5CPxtUwllMjk9kul9XFYH
K59av3JQS6voM05NaDHrPv+QO+7qQhaX4zV21OsPBpCwGL5lNv7d57fR3cfOIdf/uIGrF24zvWuq
XyazPMX212XMgw74+Krufw9lLg5M4MxiTUHTSz2Ss8Rc7i4bewqiIPqUxk5ayMyK3iPO4QIUw3pO
/LQ3EXYgwqvbnemgjNYunbAOocKl43zeTIWLNqgF11WZAggFzWCMtI2av9I6MaBfApiD6UqQLc55
RuQZHSGMu/ugg59/nTpmUhYxHWxf5j4IrSVOBdyb1hBWZwYyh+HLv/gXc4wdcPdmw2Ue/VvW7W+y
HZhY5gwb2HwnPq1sg1OiBLqguIkupnFp5ya1zWwcWVdNRAjPukdOCUOM8Q/ud/7/NKsTdwnNqjg3
Vb+OI8PVU8yzPuRleW357MqDE0zGwlMHxECjcoFUWAH7W+4YAgmtiRUK54pWpuBXEFV/J4HV+Kwu
GYx8LJq6EGfNZ7WKeTr7V79vLUweTL/yOYdsAI3D2p82JRjDOTi57WIBkUmQIJHbk4InvT55PGCx
XJLOJ4zLVSnUYVM89zuJTpIfaoiosVLAq+dxQQeIfbNcsep4ZhdinPw1FRt1HJBwhN0nQ56EpZe8
s7a2om3mmPHVngvXaW0HlWH8o73MajFdyXHty/6bIHiT6eYnFHze+8Ihomjt/Ek/Rs1yTi+uoH0+
jGoUcTDzCiyZ+gC4imWoWrHCuDGTaYXUhHed4JLqg8ygtchDpKdikbCUXxiUyyyVBpLVvrs89BII
HG9ViSnpycuVapoVl7ajJZqzWo/imHJldG9fA/WoV9Yp2vYSKXOUIhyy3OsR+iUNAeIXHElqmtm4
XEI+hfUfpZC1VXWzr6rz3i0K4pKZ1ro/ySh42aKK02RITMUdZOlgC4avXFOzJRla0NaXuWanuBcx
Y9wr6tgQQXvGIzRy9zEbdccEaGr0Uty8laGldBbYicDD6/LeJq5mmP9p+FDO7WmprdWwTWCqT7b9
PdyAmCGfkWenmfydfmMDxVpzEWyEYvBiu70mx3g/eIUTPuAPIc8g9UYBjjB/7zriBP9ZhIT4TPpt
HEkftQdPCG8M6r44WyyZ628vGfMBjL/Nu3SDFGfIz9sMmyO0Nu7XSOQulnwApCYhfNMFfDQxrQEd
jOBw7TGuDFp7fojADAZ7B62MypPx66/sA0qn5OtZzkyMGR79WPLBeChTgAZwygVXd8iDV6F9m79A
Lj+NAPkbby8uJjBkJZPi4A9hE0s2V1TtSV130G7WYOB6b0vWhK+WW4y10kuG8XjMslXo81JVbvjo
NApbscOJeOAzII2BDOUnLn5xenDCrGtnat5BRWB42ldlN6jYhMxUsQ6GX3SRNDx6779K3SQABplg
+X9VlKpCXsBOwKLdYEnshu2qn4vStqS+8vH15mWBj6D+c622NdkbdZ8sD6yhP1dDT0uloR9H1+0z
kK4dlNEktw0QUmNzOOKQ1d14LL9Ovw8K6ruSXs6jRnCBwe6yjukUdv9nEfx51aVE3u1nINMng5Kk
mq7sLxqAjSYY3joee2nHZlJraK71bEiRDWBLzxWpBhQkdf1ZG77OAA0vO91Ns1Lt9h6gEP3i5zLc
tBr8UCreDSwAQuBGKqPY2X9Dwrt9ExQTGZLal+LTLPS4EUcCKDgG8Ei+hjlxh2Nmt7KfgH3Bh+yM
Jx8PdA5EZRqjsvKsV6POskrrdf115KCnWpH326UjxsLJfsjU4Q9qVrAVrvLRThKj+Ss/0Bq9wTHW
RyR/kDZ8MAWWPjFEyU40zdCJGvhAdhuV3GnJ0e10rAsiJozu8VC3/4F/LqkFNp2r3xx3UxJp79hc
8A5YraZ35/Du89ApSn19H4TkM9WL1vmJoYnizkOZ/eqwqESsYFLz8TXJ99NjoaQRCrzvfmhezW/E
91Oho2utN/CRTrAFuCD9rAbW24JqYSeoW9KdLsGLnx9UNOYa0gfeDn3Mtm2Zzdx7cazByZ3HLpZp
w0K2IcM4RovMqrPSu6pGuoIhYBr+EzmgIlcpH5vVcewhQkFCLCnii57dexaK333Fs99CLJNJhalt
oZOd/VRVbZK+UXUjiMr3sNJTDqVUpSgHN5dt4swns0WPhT8U4YmwLOOWYZwCCC7KwSqm5Z27KlOv
piABejRcxQZde5a/+TAgRznpf1tL0Ogg6xBZSSlXoeXfPulinLaQVbZQsDCrlMf8fz91NJWYlHDw
20lBqoPOYTwnP7uvPb6OJTZL9Q/8EQl4bP4NCvjgvksqfCFVqS8KEpUB1dejsf3K/Cjrp/aW4LQJ
y5Ezkm2mLOzCc6vswmE5fyrffBh2oevRMcIIxWwk1ZnCj8k6N3zyUOaAxsvI86hBB6VWfaRC8EQf
8CE9m2higSSnptQNvMSyl3zAQuEaoDGFBccHB1Qr2UGhheRWBppb9UAtrEVLKZ8Q8MkzdFgYJ2A/
of39i5OA32XFPiwj1Hrw2J9eOEwAU6F/Fc3nrpCBeGhOZsT4YuIB3B2tafthYrdi8tJz6UjEiRPK
RoK/2Yz9+dawP8Em4ljYQlr6AQ5RX2xb0Su9LQSZkk5qPufWRS5C+76gwEOlwWKWef4yAjPzfa+u
989Z0KfESf07Z7F6o9hcHPwnRS6mQ8OITdsl1F0cGs0uTkVs+sDPyRMEm+gOUCGogPB0fgYzHvOx
EM0WOAzIO0O1x5ZAVkwNqOunBWwmVl3rjfnApf0Yra5AQnbcgchvqwEuI593bcSJSKKUUsdxTkII
s/ENeFxgsIrUkV2em3cgX7vRrgxXC6rFqba+nu2OZDP2eeL8H4OcXiNHH9JzW9bhN05C0Gk8Aj0L
Q629b1ZPrtczV0bcfKS+AVq7kvKkSLUnd9gp10EkztNT4gXx3a2JZnw/5ccLEMGu28dGFT45Sd+z
JAzazYVRplzmOs00sk8/g+NZwpSY5elMem8tbaJ1nUPtmx/fW+2iti1ZSAAPHn07rPVpYr+eOBlH
9N/gklkAUVss8LaPPeD+Y+w6DMLJIi8vkInEbSy8t+2O8pS5doxCjOHLQPb1L8hY76JXUjKupyJR
mMwkzNQKqse7N1xScoAUG4e6GkBOBfg6kOkg9TArDOtoEXm0vRyv6Bvl1qoMsd86MdW/srJpjwBV
muJFSWokkxSLrPaRYGESqn64sjQmEh9lT68ee5E63UewmZ9pqVis9OqULJNdOXxaYTUK56mPhDe2
0TX8p2nyYT5gmqAkYeSk52dX4a00ON/shkCysGN0Y7GTq/LTzHpVkYFOTURfoayBLVXwnPOwibxq
bdVN9M17M3SvcKXjYNCgc9oVNo+KgWRpfC38Jy/tP322tphwtbj1eWi6dzYxFo1MllJaAk0x28Uj
MqE/KSzHJS+cKv+q675+zECwGGqES28afev1P9PaTABojYBQBUVrCKKQxY5P9UKfNgQzNDfNayRO
TZrt1TXKDmF2aX82lTPFfBaIJ0fWSoCD4nImb8UnmIA3lkT/j7sl7YF+wH/NaCL0rBlEigJgLQBK
+3/jo1IVfBYAYTZuqRaf6fAaPqCLixRDTHQThpCngRwerCXfEb4jcRsVn8u++GnOJlcuIpeiIxU9
fD63Dn2O4JKcA7aSr/n1/3Sz8TRV3W0zulaH4qtXhlC+Fm06h5lWr3DVjqjPiAFMuPklCbLrIaJ5
OvkSvOVA7l2if5c+ha+bZDVMU5QGqZxq0NzOJ07HzoCpIOGA3CZQru8C8ReVurvHGpwLqeAGON+C
BtDzWX4/TjG3hl0f/KDSERdwRAZZVz6K4QpngTpAVTQ4DKdcX/cbQkDUIquT9YmNn7lHqRrkcZ6N
LW8Iv+CAeGrxtlZoN9So87pbInNeSXpQmCWvVQYw/d12X/6qEkmmSeUtKTMe3LKdtNNVdHtTvgUu
pjZFXHn/HfkhjIwScRAkjaFhzWtI6T63T/rOrLdVUMQ3LJ9NAWaE5dDM27vpO0Bgvzby/es/9O3R
xljBxV6ljwUZF3r4iHTjzFYeU1lkOkwdyWU3Ehnmd3zUq478IXX3OQXtr/qOz4Z5x2HHbNu7cKWp
k90atmM2es69VWwO2o1qKIsUY1AUFg36ia37FachlXnbeQeKktynilahKqptfxxILxe1vxpQjqG3
LGwn4kfUvxHyYPDAnt3CCXeYbvSIt2ZJLiZsvoxkwiKCeIeGBoUvxB6XRU9zcyrVJ8ksHLisq09A
bttmVtMJ8CZ5wROAP3zpdUz4c3BOfGsDQLlULZC0MlKJx3ahJLgvsn8lx8klGIItaLFCJVweLhoO
8fTjrSl7o5ZW9epPBE9Pj7WCylOSO8M0ojuV36JvbAUXl7fouwDmhamAcPho+NxusRIik+g+sumb
rtGwxLPga9Q3goGU800J5nE5Fc7xfj1FD7uyRN2OxfloqOLo65QgGj+v0XhELPs+ziuNVwmfjIRH
iUcHWcUhkBPzKT9gCh+YUQXvDEjqkH+IZArYCsur71rLEM+Vs60vhdLHnjK/3H2br/chj0bjdKUR
A9g9NKlI0xfdrWL0OZbwT1vMovJ9fzEgsXZbsaTzQCT6bzkp5dJronbF+DFctwUiCW2d8naUpAi3
dy3dW+x+2ZemIaJFgTMNkYhoZfPwOyGKsSXY823rJzI/T1TPP8UAqlifBt9LIiX9xGeVccWXY8qx
lr8UWTCyGrls9P4MkUVmMTeeNccA1PqqAskYv0Dk9MKsQxQ80HDsUHPXCoGfBdjnb5YyabIh2pY1
a5szjZRq/tWQBbpoWvrSO+GwHFfYFWDNeNxYaIm3Gr5SXAUoH9Q2XgkRZ0vmrbs9lt2rzPo6GjUZ
/hqu2VIHwln0BfZVWy19swB4kkeBNkVwh/n8NR+nLjamvElyswqjIO5rTta5ie6+Ab29zC7U1hdE
0hlLUEOo3yIbWWS6TVVX3L4fLZUnsR3dIfOwJKQiBumC9eZOOQ5Bb50y5skH3/NJ7/WjyP7+SeL0
AGGWOC4z1AfQUP+qiJgt9/blL44UdZvwdK1mU3fs/67rUIY1oqBYu0LaUE4enlOzWnxtgxkxCwLw
1uzs2SYJcskvsf9SUS3oxLY6kp3tJ23sN4csszOXvtmuGkSSYuKjT/BVhtVGj9oHX2+4PP9WAP5H
beB4jsBhW/01XbYHsgjwFNq0YVCxb5rY90z8xSHWFi0GDccLkyE8GktCqjqloDCY6dQ7FMRAnv2T
2ToyF/NZYzhRv/apopa4Htq+jNvUL3B1RjdHtUswkUscQmZJRjSqRRYtDpPdK1XBoJazSdWygV5a
0F4On3+fUWlAY7UTFeiamJV4IH989dp3UUlfMPpkZ8Hcqs0TBVKX68RJVwKQgpIKGimP6ufKjDgC
yBd/E5Qb33Kee9d9PclFX9eebMohM20PHXLFhqIBJqOVbA3/yX20Aaebcxhx7Lc7UP0/U5zQXC9S
a0/vAIeN49OajGmgPzr9YvvWXdGsdNqNssjuS6JTop3CBJrIvTJ64oZSzXDqDFNfkBMJxHzjwZ4U
ntHMBZcMWeOuhTJs33AaBrQxmtePr6eY5oP23Wpbs8160NLJB33Hpe95L2VRVY/wBpf5PLpSpy+n
iyawC2nU8IuXuB9iwNNRpggRYQP7JLcWRz4fUUmxLSQdgaY6LUYm14hqWSCDse57VSvPbZVDBH99
lZaiTlGwRjMK11tY9c1dYF9HfUZP9gYCZMqwqYl8nQTVqTeCppDcJG3ja+OP9eCcSqdZmc+xX+K/
UUHBPkKxLVC5Tu4+UGknS1GnGnN0SWvJZbglrLZ5tnBF9uaZULjS4h68mNfQaFgKMg8pe2ekBAfW
J07//MwJjwE6co9IA+0coQbD9lwonnwGaRrX/QnxYQXkLOd4U5s20p2PZh2jX/OUuRIqCsf6Ex4u
X4swdPWv/4LmSwJ9Wk+hmvj0p1YuJkYDC6Dm3wlnH2LyajnzPVprizFSq5sVhQ/9/Vt7jDtqM2ud
x/B42ulsqZnuzQ1daj49UBiRphTymj1y4osXCYxnlh+WsMGMcXUqZJSNEagCCGdH7mWJatnd9mXJ
fv7X9byZtUDZ2lpX/Xc0YKpaXgp6lApt+b6ChktTYWBdw8LANOn6AT2AXuQ8zTSNZWxGJ20zAUNF
RMASlH0OtG7M6qpJBupXNX8zuBP7fudFzNgVZNaYOv7YOYLLzLPycVYpheKN8YAizsZ4D2irxHf8
cPUgGEh08/hNMEhJT8P1medzvcFoczSdv7gq1COZeFS3m6ViF8najx6AEhJ6g3ralHGtGqWctXq7
KE25RG0Mnrxh0oLef87d7gFhOxtkdUY8t++aFVPqG/SuBcQumNNid2bMe3QKYcpsIZwWTCHMbddn
Z+U0WeQC2wXPzQ+tp9iw71Qb9AG6Zjrh97q6aZeptNS704y/10MwDRRoIDUBKgbPe9sBn3uv7Mff
QfQfdX/6YzU7SESe2lG6TylnE8v1rwdwZLFeCfoGb2JFGdzC7Nh6/14QyNwod6JESl1RNxFZ650m
ZySJB+2jssMjt+sfmFer56qvgpcD8NIUF2MGe8/TIUIMH+rOmBAZvAhINxrzmWDtgDz3XUNeHho/
5X/6DgD9TI1NlXrNZddptiwIQ8BcdVdTds0OfNMA5x6UxDeA2cZseW5KRms7qYK5hfKCArCbO1vM
L0Tj/5xOcgH5WoQfFfj0abCsf/mfLWvG2OFrZhiO51lgSxoE0v7cwHQiZUfk8nkd+x4Vwakkv+Yh
2eYBcT5qkYWhJivyHh3AqyzBhQ0WqwjI5CbFyaM7FGg5L1RB4WwGSpk06pfIb6pq87LRaCLJgB+v
wNUUzXPio1BiURVZ0NUSrDJRuOX0BWDWvkvROlrIbyzztVmelDy2/VkIlGONG/QhS8pUqynmIgoV
ZVSBJoegjytW5nBWMAJu3F9EhuLCmuxZLJqWxSFvgCRuGlrwWmq+UFrodkMWvNC2/TZEwQILRGsX
fN8i608Cj3+Btxvida8HQlngdsfj+4JHr7CW5Y0EK/1aO3vSgO900uPCAe6AGUvX2up+QMt1jcV5
Q8/TEnlRnG0a2pGZQ7HBZmT02jS4ztxZIgdGPH7IQ1oRpIDZjMwGl/o4WUmmCPdSIwU3JKR6c72z
hbXKBMTI7///Qdpww4F1++/NtVEcCXcmgl9udvlBLGseetTOmFBpvz/udKFyh11Zzt3BGahswJ7k
TtW7lQpDqnHFMn8SQTJG/fSjDXqGsURPHn6CbpO2ICAOJz8UYvHHpdkJS77jSkffNQjSlPSqu1fz
OumhmvUKyBt/56ktdTfszO1rYbP1ezrdvZyW1Jks/vzSV1K5Esn5ycQ1Lfm4qp4nssZY5qF8lqo7
FdOmsK6WVD5uwezJyl1h8wuLT1SdUteYhzPzkIIOEu0YX557M0LGsqJ39LeTZ25xFwWleXRflurk
O41Ye4EAqeAC9agZIdssjNndRzStkHO+GSXHoF5IEWFcTTujaGZVjxUHHqN+K3ABSctHUMTtiG7N
jIrEg2wbE3qfZDox6hhMrFhGUoXqpU63ER1hw9mdUtd05cFFz62IdrZvKq6Pt++QC25+UXNNS6fh
ZdoW7/yfhCksoMbpraWbvODRywhzQsbOMuXRHalGmb2jkgOWhmJOrSU2Rh46uclBgFEQsskheSIV
XPSfAnfcZ7vGvXqQIC1TXG6l/F58kdYxV1roL7/24GwQANy9k49qYYq4TwNJutUdym0zrW7EFmVJ
F6pVxehdqFaqHi1TMOwMv7zBpAmhxsuE2h0qSWOYHZZMS3joNGIA25vhDFDJnCsNCFYteQGAjdHl
hyX3snxUSAMxhoaPgs8APNUbTNa+twM/0cC0YJZ+7n/1Y5FXl8jeyc9oaFbt0Ho17TlU4LfSnDP+
mxrT2bctfB21fIjTfDmy/2risqBNrayd88Qu6DiMWwM15VZbQtY8keCW+fm5koUgl1yK5V88cT0W
SRTYRoHInt/gvIkGRgVU4nRuxDUBWgynbsY9nIkmqYuS+LLL43IDv48mN2Jb0NxxeuZYEYlWrm4z
8jTJBIdlCjrkfM1UPWNaQQ9Q1qd0zqu+efm7tvbZG9sQ2YfQ2U7YKbwTLmxPSxMwkfuPwLardPpI
gUKsVbzM56XRCbW1tkokQdVhuj/0TL5YVoJZ9bCPt3Yj2WcWng2EGIqfERj+/Az7p5DDqisUtda2
ldjGJCfJ1bcPICImX/dsnCvwCHWnVwnEbUoVzDoi1lmsF+OIWc0k38phjDmAblAM73/zLa+NJVHN
2zM/IMyQG9GMZ2h026qgniSeGWIDBcQgFiVFDGS99t3HiIfH5yiwvleCr4DcVqIZhUFoC5dUrdan
gXPBH8UV83gP/qEVxTwC0Y71QkE0AqIP93dRRB6ufVsu+obGQ21Gh+KtYYDk4c9vOEgcFFLWj/32
n0Os9fNf7ekfcquJi/VBfbSMHsPmvUnaTdHQLLkAjLf3KA+EcglGtSzx9DqqyNx13UAgpt7Zy3QS
GctHKNejFZGHZrRzD0diJA82Rq407z43SSvs00RaKn7WsgAG1C+UkGcF9URBokWXKHHBYbrjXMwd
kXKidPkJf6Ys/j83c9kynxlaGRZXkg/tX0Ygi0ra/xBrPadsMXwPZhFBVv/10TAT7Y0akzQfBxr2
Vhsr2xjyF4WVq09E9W5ir2ZUNponswVAMn7xLsX7didL+rxz1n127/JBh2x0zpMKtpzcRP9ruh4W
tWn//R3NCVMR159ndjl88odzMOIvrKp9+c7KEDrJXTQEJuDju/kfRjXZhNlMK5XvNc9X1ruDlAee
B56POg9kD//eQUNPLWHJI6LJzdFSJ+I+yAcnP+bvwbiAgThZMZ33+x40bZYN26K+JDhGWGIE38sc
Z+SZLIrWhfiQPHbs5fBz6QuPph7QH+IR5sGJZ0FpieEhEsp6Gjq/svVDo27UoUKxQoRlJL11JIag
GSKVTCOA00h57Wa9AjdXPAOizHCYKg0n5vfEA0alI3aTlvYMKfX68rEJ8GZifZxu+QhEp3pQMOEI
U8Paanks7T8+PIitzFKdWcfNQntlY7Yfavbhv5dIunul3FdjM15xgm5+Q7/HGlJAGZXD8agPjswl
HekyX34vNucdrTC8L2AZYhjvR5lSlVMNujNBrNnVa5uCjJEQN2WdD9c/NyCnbPNuC7RERg41a30j
lL5gaoghYvIbimmUZWEqijyOqMN/gsEQmkaI+X8KGJ5fFLF0zWeXUkQIwrHdqlOcGPT1UyjJVPCM
QJGD+fUTiNvdqwSbvCjFnKJS/H0yCImb0vStKqk/RGW3XoRFMCmJ2lUHStBczXQgvukX3MCBPrkh
hsI3ZI8pJYAhVLDqLVNkXFRbieVJDsKrQQQiuGgh+yP1i8Uq5IyuJwLllwJyg2b5LjUDAqhnUmxl
Wmvn1Xwi5UxUPgVbWynHzhrmE1DOWJaqWtogDGz3DsHkINkNLn5cHKjgpzD+H/R9RcXIR7o7Aog3
cYei1hzEUI6K066NaF8FM8Bb55hHUYwc6brNOhNZrgOTB4UwWgnQGFlqk20eRfEbEMN7DGr+3jNk
o7q3f9IRDoAk8FlEQcED2EYJk4yecuOiFFt0vlkz+FDZhFbqMomK9miK644mV46QS2fAQaUWabSB
zLeDGImZNzeAYWMfBoMWq/H53DcIEAuMiyb4mCtTj0GLz1+gElL7EviDL3yGEHgf7pqVQRzoKmHk
DH1Yh2PXE/hjZCU1MirN5Iy1jHKHkAXjMQ8o15/HKc22AAl1nKhbLU1Ln+95nt3Dx9/hbkjjcs4P
XylBHfO70P15Y5KRcZ33FlZcn3lydn5RZDBshnAuSIb5spMCnx7VoGmbMFGWXIFB7yggSzGiaS7z
blAWnjvnBS4tBljQhIj2T5uyn5zoy6b/zyii15EgqYSyJCcHLzMiqUk7dxLfBGeF4HloUtg8UPAm
0LZIWy9QVfKUOYV647WxFCHWAcSRUe3HAtmuGAuNu1HCkfUeiOn9fe5anj8+we2togqM/1Rev+9c
vnBUsL4bktz0WJQ+IZw5ZknovZuaIrNSJgORCaUQt4tH8y6zHWs7XKqPlNSOO0vSz8mQPlefrZcQ
hQRhyTbL5+t3R9/TVqRL9gBmCfSUH+qc3TmjqSJiQ2QCBejIqDaOc66UiP0j94x5B1epuIU9zd3R
jztClkknJ0gq8/WphzoWEYLS+43eyMWYk4SSNjNhfOT9c0QfiPgNwNLkBwNPJlgTu5MA8EYgDv0g
uYPiDfSmLJVq7E0Sg9t34MJDQWL1bhEZ9qQTgfAxDkhXt2yUb2G8zhFRnIKNGCQj3aP6dYFn0FBg
thVMbd72u++BNzUIVAVsExyRIDfTCeizNU9u9/aWCkXYPPwsBk15lwget69agcSzHnm+gwLpQgBn
Pm4Zpqlr06cmkYhXfdXLWHXySb0oIqKyOAgo17eG77OXoxp1eR27HS6IdENK+WWbyhwKiEiPNRL7
dsohs32j7JEEdf5IaqXPCNR96Phc7kxsC/CBE5OCawmHz/ZLnFfWFJMh+M8ov2V36gM1wW6G1CzI
znSc1B/pAdPHFtUvD/wOwqqz35pL54ugoGZhW8RwiqbghUSWVr8RHMjNClV7Z6002RijeK9EFzYL
Lh+NJCE3DAvIr0VYzhGj34CfM62YfOC+/cuxwxqqozI8yn6vloRpBri7lK/x6uUba/MNzrH+mXCq
cxURP69jsLo7pbv1TrGn034eDf2naISzAfZR3fu87GNMoldPxjmXaDI8DAC7ar70999pX9lMQHDS
V12RC8/ScYMOFZTvfxaW3heDuWZhWhk9Wp97WJ1CrmJMCObqvnzggJ9x/IdGF6cMmtm1kYDuQ8nO
/c5tpTOl9vGh7HeUqmnPPmmTBdHB6dQHY9cy90kudYcbjEM76MnQtagUNEXvxDKeEcarnLFV6Yp9
yg0y8KSfJ4ceQU0bkrEnKZqKInkE/QiPeyYvOPsT52aZ9MaYeTJKz8NsJwAZn+Hxx7Gz3oYg70Zs
llxsqnvNc5jbDPUO/wYzOAn1vsB3Clvucv7JhVKWSPz7HqTEIZ2+plK6cEqaNR4yf25XV7ugSYrf
Oz2oeTzncVKoR8wWvioTGfeH4p0/37nl2+UmlpUhjZOBswzvlNmsF+Uvbce7hGpwhtx+zJ0WjE2X
TRKdpcEJQ1pPYNQUg50H3KRXNdeAB/1ognBSohwu6iWPfkPALQ0WjMg/VIilvGAqpkvNXG+YQ4lI
IVZSeKsWY+OJfNwTRt1dGy5OWkNmfDiWeRi1mGxO5LWV7OS0IUXZ+XC6/tnxy5iJlmQWh2x3HVon
vTPA2PRTX+DjvWDm5faXV/xuz0KFe+UQmXX5lfln0PlnNlL+yH6YyOmxqQjxUrvac7E3oljBzUWa
cxbOuaoKW3D7l1Zf0Y8pu2jjbJL23qkP8H7Xq9re+aFWZzs6c+Yu/+iAvFjFtTVH37RuMob65nJY
SFt7LmeqxktvhI1bz4lWoY6KKK85zEpx9se9QO6E6+I2ejXUmlRMf63vwXn2xUbqoruNC1jESCoN
NKrS9yBq+EIYZAHy5E2LCzCgO993+uml6Lcb54RGQ8cwTAtciLDQpPWS7YL+sKx2MibwbUPG8HZN
M1caO87X1INmoPmWqZRH2AG5vevAlsD158GkNyRpoLCex8TUnF1Y3v59KIPJ29mvVP6MEylj2RYW
M0ZJiW+j/vyaa8aFIROt1hgZNbRJeqePBvZiRzjLt0xarwiF7UVLmMTMnmSFrux2lsgjBmw1Pd0g
xUfA4h5Babb94wYCzoR6Lm12XCPs6fB+ctKpo62MJo+L/7F91fHQ1BxbnKPJ8uNbthtAQ+jvElT8
TZMw6mqNLlSMJeaShCUpjXnx6D0Qn8uwPiKksgCEbX5uvGSMI9PWoCFZJNHF/kDWDuMds7UoY/0S
0tyCXRQkFTCydCVlxndM0eaC3TmMibFZNP2Ezlraoi2Z7p4NHt3MtPtkMoF/haAK+TqWZJDDD4QJ
prBQnkWVtPZmFdIKo+XNvFyytQgH9FFHIEPKAMJ66O6z5vtil3MUKObISCDSXuWYqNvy/ZPHouKx
W1zgGqewrJT69ZoWBAObBXsNUrfsC928rmwcy9bgLYOHHkwnbOmHFVM6t5TBdPLMIGhVeKxandOu
US2HlwLo1LqK+Q0y/Rq67sNnL7FUpy5PQWr/nOYOSwxof7fBFJ+OYJnRXuvkDdEdifazwl3jakuD
/NyssOEhqpg4+SBf1xSJ6lR4Xnc8Jla+Xo0DsltGmBw5Xa5P/leRiOwfyCIjA5MOt+lPF7Yah0p9
GmlCvXrskAJ7yc/PDwTKJwI+1SkqtW4RetseYvImsRK2B4d1ac5D6mJkbVEO02oB4+UEeWIXuCai
7p/AaY3O52o1Epyhfy0J+fPodXoAfB4SQ+8/PC9hY4SEskNOLWzDxcDr6LDt5fiuXTcPDwOQeSey
xoCAmzhTg36Tl3x7KZ45JI0IjZwe65pxQIQ19LIzA2kPnuJvML6dEbwyxYznjwDWoifN4+1cPId4
5EtNdTsgzMu4gu7dcoLUq0meu4ElQz7dgnbUlJBVnwY0ATDxcgqLcCCHg/zCoO59OBMOETbJ9lAK
thNB5x2rK2Y6DwGgdp/O6EzziheX6fFuAqsLOcpC18xnDQT6GigQwabb/AtUt44wbKasgjBuNEAI
VyxE8uLnyk61eynBKA0n/0oQUBzZ9e5BQD6Pd9j+XTB4VO8NmCRcNEMHzHmQ7PvAs7FnJ3JiqOdu
Le2T7nusT4+3I4H3MMeVK05xqmmRNOmGxKG8qt5/OAWO4hxPzIko8dPyJ1WaZ6jeF1g2z7/hWLLZ
fo/yCk8H18BRRiTzu2tDmOBgexyCx5BALjSKAywcADr0fTZvES+kwMXi6ZMvYLRGlTFCMvMkzihh
oZqyTTrJTQpiwkxi3jx4pffdwOjvRfho8UIn0U/f7AF4sRmvEw4kZpk0y9YV+DA0V4CIH8PJGeZX
MGOkoEKwNNFrygu+kKM8FAohwZjyt2tcG6khXxmLP4poJRMm4shADb0B1zH8/PbTwGsDBUJn085F
E6C2+MD/muKLP23thScWX9k6zf1ETBJlC2Hj3A0p1hg1WEWv4NJ178DbpxMzsrcosyTrzSDUZXx5
C1X1ASZwbpvpvxHNzfaFuWnvnNuSswx97MqTd9WGcGPlqkk+x+mlTX/mWS2tdtlfIy8Z+SgJCs8I
1o/Xjp4fpKPgRljOG0PF4aPgK5wlkCQIUU/+4FyvilkQAaVVNrBCNu4SStnv9JGh3A2wbunYTg3/
e5JkrAaeHRbQptvWEvS/rqlQr6eTM+zUu16Ct78gSsI12b1pynLT4250HkQtJHVSlDA9eaVp9Jzf
i1RNZGqgCHQsWKhIk66ICyqVLgeMXJxlaOlJWiuHsRMYdsYLhQTIurwkwsVsQjDCGcXJ3bDP4Zxd
3M9LVtZ8Z5dxjMQFpjkKD/1TCXV80TrdE3bPb8MblO5fXDLWTNX3pt0kQaYTziBx2fxF5EiB9d4X
4zpOpmho0oQvWmOb+Yt40/EAS2sQ7AYPzLkoc/tkJredTYX5nRMn+FNLeWrbfCQHxTS/5we/3bwG
A+dUZoYgwtBScIvxZJ44AR9Hd6bey0C+xeABWSIpbrhnK2SDh5hTFMtYDuG8+6JrqBQRIfaed7yY
DbGmqkjjQCegJoeujyJdaH/q8adWPIy8u1OF6OeH+wZvINZAD/nG4X9J3ftJF+4/GMhO9UMYoj/p
Jb7KiqC32W9YJ4g21ur1z9wdUDMKZ57OVwGhZidy+hq7pdAdLwpCq2oPh/JFmOI4VF9eZ+nZy5BT
Nxg/cxPsthQB+bar6liylkak6BRzpd6bR6tevC1vNBBhVo+9cYphi4Uf25d0PFivCKVKjwsmoO61
tCuLSjqqFcvQbu793RY6fLwmAOJxVMxKlm0Ku/+pUjRSl1BdWIWrha+FnZwzTVNcqIIxFIkXXJsf
68gsfaKEuY2WaaZqSHD9CgO0kKytBGzVxhBUT8RiWKhokmTFCI9hEQo4qCrwMhPv2Sv26GSxO/dj
s+i453au8Z0BmIxQ8T68NyRlrLu1x0EiatwnVtiLXmbaqqztx3NPDBz16j+Jte9M0rjJP5icYbSe
6+awuuEHt70eubKQyh15vugdERKiqFmLMLmxyVQR5tjOHlJaGmlljYt/AA6IKo5VsCW04DECUxUD
OrdiTP0AzMo9GyhF+JO2OKqyvfV/Uf/haEgANYwP3zlXLQypGGz00DgH9xGVjBGY/Xi1fIcGScc8
hTMaZYE0NWb5sxBieH4Wmm1RfNEX6Jw+CMNbdzUMOHLjWbzPdSP9OdIB5thHanjoSLm4aHIDRFq3
lDKVVY9r/CiWSpIWQPjG81FJdLx+/vDRGSx8VA8MYKn5XFY09SssSt4B6Dhzypv2ZgwvH1CkmqWn
QlDCSMmGO5d/SbVo6RkiaPWP8F8G85ZWXphkIAv/X+J25sxS4PCMchmRUqZAgZp7DFV1lcSnhomv
A7QXtL0HlGs+1MlxuHlrxpVOPz/v7VWS7wVtuLwDtKOF+KP1dUxVLNBH5b++aF9/3rh6r/t8lJWJ
pMry8QqabcH4fXCd99tuFnKvpNInRdx9uJsik7+KuvKwpZag94iKh5ffqRxteZhNz7vHKRWxTqTA
gvdvrxR90GZ4Zf/ffnuptf3Tk6n1I1br/fylSVtXipTBDVEPZ9lkTkaYl8AgZ5mNd3rhsVb+fzTz
7WsTWDkrW0q6uieGXZB3Bg3+C1CT0kj4qZ9E0DfrBiymQuC9HAPH8OCfDO5XuQ+9FAgt48eEOZNL
N1KOiFJNK6g8IhirV8N5A+Nlg5CUTBFi/RK8lhZrjwZAVEE10szBbymU7vZ1S5qMlgS6SwntQZXM
a0XJuoSRw3sYjTxJ7M32m0ReG/HFZE6rPcrXFOtA17jS8dzHf784+IUJOr7DRkHQ+4WoQYwcST8O
DbWvESllXT9Kiy+/rMTigQ0xuib5Tj4gPyv9wwLTL9J0xSSrDSoXhjt82Fyos9xS5uh5QzCNUbTA
X3UoIVJRIcMxtfEUAL9wp/LvyVitl70HIEpjGv7R9oVOI2AQJtKne8nDN7U/CGSFBg3nKS9AjH63
cI2LBEiHTnAImJbUDG7s9XQGxmdqXqgFL+QPC5kAbavEcu5IrvsxSGTeD6ArNi2IJ09gCiR9nOPt
Sah8Lh6e9Rn2Z8Q8r0aNRLn7ifXfu3NYQ7TemWWicVj70U9GW1dsjQ3eRe71ZJ/cGWsqD1y8CiOX
dGyXtTYQRogldj6yVegglGbQNjW9lx2x/viTNbS3YxCP/GMXAVOg9xHd06mgCyFRRJ2FfluNshA/
wlLYWjY/57YvdRK1llnJvqC631rNon8xOEVhExXMAoyyXtYSGEGEZ4ysjmigtAC6uUwm3AbgLG/h
TYEz4IHQ/Bb51F4m5NmAIg7nmARZ3M+6/tWV8JWEgPnOWiQFEAhdPEdjWKhecs4PW8JVgs+2zfRg
z3gCyz4dTezVUcz6QrVAkBJ4O4PqMja/n16nTrWCSBo4xRHvjnbtY3HmPdrjQVHjTgwJYOCQGfYo
RmyUtGg6i0i2EzOL4bAQrQUpzxPojwqd9HXrgZFgMbGfEBH6+k+2uZGX53C4Sp4YHFxj4+s2Asi4
NEZgjmDcV1LdukIAXbcnBn9GkqcQAPBvYiIfX2maX97D1XVbzAhQ/vzQ5bGLgGpL37tlgkXhxwi6
2MUpgk7X9JWN4ulWjLPUfSMVOYRF8kxHMsFCYgPU4J0vWlvvy22cdkDHvmHwp34hNmvExhuxmvJl
OC191L2atMRvDxH6B0tpPFZCP6zv1n+ryuioUgdEG408sB0+rT0R5aCHW+9UghQQfFZGVWGb2bSB
E+FIbe6AYmrhjzc8h4badDh/kORiW7ILVbtjiTA5PyoVKpRK2cfduPmeoZjDeZ/xTx5TlpcuwDCB
ZcIWRC8GViEatJnupahzTNeGJA2VxZYksMyWcmuhjUgUxAFna2EmhVYBc7vfo2q8YL8kpUhPQH4M
bJHuz+tqrGoLovjPrfXeHPfD6R2g0ZqlJ23uxNySIHf+Kcumg2MWJmelyuJALMS2vuCd7ZsXDcg4
uynzCMMTM6rI5kq1vTBb/QoaZ2WyTxSkc9CWrGK+Xp3pYo1YTW6IxuvwAerr+x3m3A1P1cqeFNVG
JD0jpzKUmfdy73+lvoD8OT6e/7dfoMxVCRW79G1FbeIE5+qivE8sDQ1bpvYpSyJ60DJtUv77BxB2
eemGlGNg6E6vptFz9jBOdgtFXbg73zY9Kxg8T4jI1HjKHQ5V0qgebzPnGesr/+UV7I5BtX2bwk29
BdA5J3Ik40ZpPhcgxpUSW3pjMicF6VXcZW1Uaym7IoOm0W6ole3B5IK3Bi7rqYOTL75F8Ib+Nt+5
uAfp+Zqsm0T7WDGGEbSlbU2MpDhSFv3Mtx+JcS+bHc9llAoEmwnang7r0gxwt1Ns5SI4hLPKYLhT
XoCPEMr0raDmjT8ygKzztEE+J8dv+X4yVZSN0BrqssuA3TFMDqYXUp50VuZqbxRd4+4u38iQiVev
DOhBvG3vM3DzrwChmBQ4CgKBiq1hODlPp9w+IwK6lkPMSL1D/pf1yL/SpQsac5GG74VXeByHf1In
7eFL2Josrf8iPGmkfTDkHdZdPLndTemfPOmyohuLV/dfHJkNe961sPipSjOYIoPmzWesHpfdvzSv
XbhA5ph99Ki2/BU8gX2GNJKCQwbuhgBGNmWhtTXR25lgAmge9Vyv+CHc3lUzcemgpbtxAQik4VpH
cSi/4d8b4zmh8uR0MjgLf5xUHwcjifWsMktpsHkO61WR9Gdzj4ljlUaAaGP6TAvpadIf3JEdz8D6
2cXOqlNYD/35NVcuD55C5t/AjDqNxKSU28ThMfd4XLZyQM3IjBmiHqopcTT95dTTfqs4ZFqlpUJp
RPpzhA1NPEKmyjHUImf9HT37NDBTATT/8ZMVlEjW93TTVJajR+AjVOIVNcgWz3jAg5R9xBlydpYy
e7UGdvsRsCjQ4a2MM24z+r3R+15to4qbO+012w9zLYU5WisewAW77SogbsqR6p8zqUTrpe91YO8T
La/npc3kawWuhKFlgrGOIJuJ5YJ0sSJ4sbydqJxCOX2Yiq/FtdfSaVEWclrHd2OnAvznHbVvOqoA
Dd1+dL26AF3NNhtTLNU4LVVBXa4dhCSKseAAGoVQ8IaAUU2BH81Smm/uLrbJbZcWKq3JERvVCfQk
c+8n9232G3dHVYXS9VMmHVG7YX4fKgLzw7osy5UNoMsYIc6BPP2eMu5lL19dIGW3T/x2x0lRuKSk
OC1ZgSqw6LTk2atVr0EINK1Xh7t8caZ6++Tjps/gE2gQzRJ5Qitdwy8xbIX82fCzmKglHqsXtFNI
+VNbsMm4c1iD4GI5TieCEdNrbF1aDPyrEFYRI+r1PqDgSTTLUcpA6vFl9WqOzw0evUjv5ZCHvUv2
u3fmTglVW0tSOVTcIF2fTRyp+0pZmlfDrUpr0VcJC47+VQGgmCKl0nfcKyPRJZ26BPRlHZkhbcRD
xQFUmYNvjrs7gmsRrc9uvT9+0ap5E6XzbKMcKunLEkTs8udpBDjGlVu0AiyraA82tUabtIfsyruz
v5SnFvevPabWaAsrKuIVKTR+dHqcsv76JI4aEtNYGs62/wkaE5Qr+XRlY+3p0N2b8xtz/pAnplA0
kZ+ouDZon+hJggYZyQT2Y1MUcL7h+I9wZlpImIIBlkXMVLTfq/pF2q3Im2+6AHC7rHmGcHWfb636
J+jR7dhxD8cg9wwbQdSYFkyVdsz2U4Dldf7sys8O9DnfXswpcCcx47fPc5Du1fBDWAx3ru9U7n0n
SrCTvXphfhEpK+ngCmK9O00xZweIGqm/SXL7+LwNghuFAi+avBtwoiuCz+BTWaxBntPfKbKzg6Qo
LtQTezm/rTUh0pfRp5kxKo3GMJaLBhbqDHBcGS8WPaONdzAF68CJxdziF24kaReJl0jbBkMQLUQz
rgLm+MUjUQdtjAXKFjRyA0DbWH6fGUOwpQiyE7O9cFyrA74o2INlC7OVWfRLMRhlse7vY7WusreU
h1fXpeXrgaycLtgalWfmPzD2YRGU/iYS4cGL5K++cUdJA8Je2cOK4TX+lmcL+MNeinWWgLmX8MC9
B1S8aTxzpOjGq1Q6vVdJ0kItg74Pi8FNwmkAl8a1XUNhuKPBpEdWEG9diWVBzMTG0JbmucOAj4tj
EDB3JzNg2XgdNkzJcBhfwWS5F+QbKBrAERIcaWRQQ2N8piuQVq8Sd5Xyo3q+puhPsZYaFDl2tG1M
QUwsJsZeLCVvLe/4nWXJsng2JhzYPUIBcfElCJk3KagdptUWmDtu+BogDU+ha19w+xyxJ0hzGa+9
YpUvKNcIu9gyOlT9dTpJHAsJ65l3Xs6jczBWfC/2pgKXyRwk/hklgEc3EncGVSbkDJ2ZQBhXpMvR
fp3HorxiR1KveSpdgRSvGNPmb0F9qBWiDWgZHdZKgswv85UzyCJKSED7tE/MLgUxeCUh6DNWRqlP
q1cWsW6qKFGBTXUM29YaXjlXeOTwBtKEYHZPSAg7b7G83YlVjSsaCzc00DPcoPNBHA8Xakt7Z84V
zGavAZwnBk91jo87O1AYB/Ob0VdU2HPXUBWp+fvFaaXqjucO/QnCPT6KM14x6fN9Gcp9ne4mYhHh
oexkKYV/+GhqvEO+0574olYzMUAMlGXJuXIVnbZH+wq2pzY0pInD9hVRnPG2Axm5IAj8z2eVjPTV
H74PjSTH/phlkzpSsLRTIH1QhSuHHfHpeoo3DJQRKIC4cYGl3/w9WQIVrLLlQ+u3rMVQV72VECiA
kGu+vqGk8PxkijWUv5jQ4dd2nInwlOVf7kOwKWBT56I3tgwpcJMk5QuaXf523/1ksMipnDTU3rgv
frjXUXSEax5tl+zqZqq2vJ2HL5CzFGUzzaNMSuKErTbQGXnDgYxgnoAPRR2ggRQgNGYCFYJ5iOlZ
LwCZJQtGL2aqVUzdbywox/Ig5X3rdSJe/hrViPRB4BUJ2DodSQQLUYh11naKGHgomobU7nPi4GY+
B9gRE3VqHX14ReZ2Kwd7dMyFs/Sye0QzsQ+bH2oan5T6SKhD0ppYMyvbJ1BsGuyakeBUAgfJGuBY
2Lk++JZ5sf5spUHzq848NeJmoI4MpOJa0QLvTnsXmxBTVXcmhEg9NnhXkJOaUHrDB0fCtJwNr/Dl
fUHpIscNI2RcR8qaq5NyJ/GcLHEULKBoG0EwHEBaiXhBWg1Le0kwXWlFAViq/mODQFAz3Em+b8M0
YgV6V0PRK/OgqRGhJRpJkq7uZPNp0DhXzF0H3YDeMJ90ENmMLGOEA9CrcdwcOTU6k6GOdS8J6Fht
uiBuot/ib+W4dhAH2U9K28/pNeYY53dybKebjdR+j5KC8ShFLIOv+26aKxjrL2jdmXaKcGWptmK4
Tnw718JTQuQBwqgO5EST79jS9nMXNIXtNwbKRBdwK5ffIzlUsmCrl7ILcM45SE3PWUY3woTeO/G/
4FkBur9OKKaSm+9LOug58YYWRvNqwnxRhhANaihNv7OMgDLOiXwxWyfL1vZ/5kMCx4IaH42Ooz3h
bPNY/b61xVnFal6+faPq+DbsJ+oQWjt0JzTDK5FvoL2hqibW+cLsO7guDwBaIPxygipMYKXtpd5u
mQqYOYZ+LIOXEi+i38Kwmt9J+AEMKvzOdvP1ozDhOAgbZQfbp3+D2ltIFanUNvO8568I6SYcT7bZ
NELII6HnHd1E5bZaZkTb7Raw1fK/2VobhMUkIr5IxloIUb7FnYgq6HDVPwyP1ZHfZ5H/YtBmFtou
AAcRdRzoTwmrf7yLfqVk0QTTQWe2hs9+6UVlIqFEzlGgdH3rJAySXj9U6V6mCMpw9vmipK8R5nAo
BV80g3qxuAO9LumAFtmStXkRYxraLEBPXva0aj+V4kWEy7zB/VCdtfzi7nKthG8gI1uVlDqKFzWV
pSbFPhoJ3snh4vr7v7pnOsBUhB3etSPfxUcfdqix0UVLR1Gckr0vqymmAf8G+V1Txc7Ju8GTVPA3
yotDwGcfpw7j5e7Zq3zB/OMLaQqDLar5GF0dYIlMqah3nudspTTTEuwB+tuXvj52bjucdg/gM0fc
/tyrwLc+KvAy8jlhj3LhHqinQ8h7AQ4tibSH2LuQidEYP0LNHCMcVsMivypvJP6M4LJfI54fgrVT
iWoCVYhL7rujAUdHjvLn9hFx4XaMDiSCuewKflmCoZZSd+KiBsKGHmmVEC3EqjQ49cb4XYLfpuV1
fbpue5AsSUeGnb+J4Ef0rOU+ploAlUYfv/niUbtQc+Fdi8R7geFBoRHTUkH99/pGPSQXbVCgfWP7
9UM5fqcxSz2HUCx+5Qcf5+w1VKQneaQvGqCQXqodNxHcikhyhoLqaToQVtCHtBazNAXxrGp++eES
gJfKHY2EBrR1E+jFhGqIBqcT7A7pMUTtDx7wSd3zgoifkVU2P1PKmeiKH3pxWBvj5qn1px/0lT7f
NMrP6i9fJ1Q6TGr5BcNYkRIHMbiotqsTvGitvBUwEIZdh78RW0OV6Ca+/8gavV4eevyqmFKAVlj6
Gc29VJBHyU+wbIExBzm/QU4S3EuvsvOeO4V0TADlOs/KSOg2TTj3dr8VQJrPnyvQe+ZnWkhQ+Bpz
LhmRWp1fHXqRP4mYYKrN6Ifcl7JzkjFxLl3v9WuuL62NB4mvn64e/+DGi+9tSQ6/4vlSfdkPmUW6
4beW75Wl9MHU9jGZAOYP/81euI2+n5J/Q9KuEWJKZ/SO6DSkdX0mbiVLSGoYaNBJCohZyJLVlASv
kC5i/ZR78GzGZ8QVeHtTf8XP6JYuV/Aw+NmMZE4XDmdh+DpFq0igr+/c82ok8TO/QxMlnbtvCSrP
fIow4kDZgq4ijaRm6QuN5xQeRd8EENzz0jxW4HeaPHBKLsfjgrwUE+82amNjQd8HGCE7aAH0Raez
Q1FrUnM6GUvQSXz4Hg6acbvMGLXb6lew4iXWmwDWhny83N8ltSC4cr+7QGoWLji91+Baoq3beW7q
cMqvRWfLjWSAt0YCLDXj9PIgiaYrWPqLYhc2uxAQ7cpRRFapxMuNYNxbnjMxIdfvCOaY9gVROxZX
i+YbzrUmKa/tC4+8biwWELz0DQB3QEJ9xkX3O8CSYwOlqkW5uqS3CHXSu9IL3KfeGPyMk1M2p7kT
zKm33XnYAfm8C99ExCxZTOJ4xU4rWMI9jweQF1aYFn0Inch1lUlWfWCj/k7Gi+nvZweJ28FMJFNJ
/c/OentBzq2Cc1J/hUHWLZPW6A5TfjniYSrZZGnT6Up5x+ymtwXQTs2R7XrZ5ErOBjRDMsUowi5p
i/sqkWv+RdQ2/BgDwlt/lc2lxeyRLD5mBpN3iyqGUTTKa4jdDQOi98EmfBWbNPpRczNx40cZDPW+
sTb4dl12ZcbYBr3XsMJQgCtTyWPGAiis+D6iGxEl4grBFPmuxd82ygLSIlUja9b7wg41ugW7/12R
aadWLJkp5lLQlnU9fzslS6Jkh+XfMISy2JaLbtryiS8Lgl3DLypVLeaIAP7yLoDTIFJNAhwgCaXi
mUFgfPzixuPhSM3YnRcY5XyGfxuBaIrnUVuCmSq6mliMPJFJizp4m9vAX9f4s7mlOqe130iFD09z
js9gYNnh/MYRSUTxvHxAFCRdPq5S4CAhOSF5i4MqHo8UCgKlibwoV3pMH1WBwvxGQncJBjTpQ1Mp
0W7Z6ej8AmaVIwspksXPuCzyaEVlSKSh7GTZ/Z0eOLKX7+MgdZf4HgN3yk6l5IqRjJjTgxxBRNhx
5l5KsHn23oCsJFTKFU8M3fBUUueh0I69IIRTSWw4RrPKnmT5VK7O2wyDGvsHfKHPA0J7HcKSJlnt
CRljGBRq3aY/izRyTAnaf8iSCL/mSWtyZVz3VOEg1aRzLauNinAwej3D2VmIn1rru8aZ2z/+/xUr
K2UbHB4Gy9mnHiNIFCwjRLu3ykXDcpoEllmaE/Kadfzns/d3qtyiyyxZny+u9D33mMvbp2Mqa/6t
yAS1fZxYPRn+R3hZm+R+qivZs1DT6HKUCSxaQHxomJbJ/4ASzqnunyubRSFPwMk4r9wUHWKob8/5
rfPBPwh3M9hesiPad29+4EIG/JVkoOKDiamKGXgfnXVRgffnnLGK11hOlkQjyQZj1VejOaoOEkYx
6bs0tTPpOknFVUN9IYvl/WsNwkRRn8eAA0RoXM7F3TElJmW6IREKXGnift/a3WJmEFRs0uR+9xZ7
qNy+K7hF1BfVPWQ1KVwoOCHsfmAMtLL69MlFcwGUwZ+eFDQ7vHCrGZAo59jJ5d19ETlRkSNOS93h
zD5VVMzAPsApDQy0p7j2/JPmIzApOvDo+r7CNHdO3jBXCaJ0W2ju9/2tQQh2Bj70ubTPyb7gTWfS
gsBc3+pyzfGJOhWSI550rx45JoOOf1eXM068hcIUSOoUZAT2Q8sNR913TXmxR/7IlhvDW+i8ydlx
2zb45A0Fk+bKFAX2IphR07RW8Xlqd51Pc2KKlU17IQmnKXlP1bwVNST55HHJA1fdi6wPjMNyf3Mk
k9N8dGRfGjSF3zALhPU04RE4sWn9PfKPWHDyDxtm+6DB699htvwR9oXu9hg6qxSMcidx0YaYsID6
0XMqQnoek8UQMlUJ6C5Shky5+PElIFWiaSC3OzEck7Y2LwToKzMXIaM1zcYJlFXA3uK5ihKGQuUG
Ww9TeBLJt4MAiHhcg4AYFhQM7KYugJ6ZPNng8/qKQ8arUMvxjnbTk9OK0Zb20A9ZQLR50P6TVAqm
iRHiO2xIcA7uFOTjzBpOqffTtOXpgk0FVKqAPQKL96dFEL/Vk6cdmMvg2PhI6Ogttc9km1lrr63B
uC3IMPZKrwKagXLwr7gMAbx5vfjykLwSpycyKm2Z+AqIvyDcXu8uOOFqehTTvICm5ZYV3QK5yIAX
JXPjF3g/GlrrFXdYHfTFM7RU9A5MD9OUCiJrWW1zPv1D58v2B5Sw1mxTfNfyxVWDITpiHMBm9PlB
hB9MnjcUBH6dL2Gtnazi/zT2DBj4/LiKuZ6+x8xrjwg29rG1FCyHjjT4xYwnZ315RCaA75ooS+S+
//o+maSKHScGQT6AEpAS/7dijI+fo7TiRXDOKQlaRAYRcxk7/WSDa8PzUYpOk9EKby5Rv3NbKmo8
tTgqegvpeBHpNp5I3jFUb0xvGS0MYg4vO1TzQsnAqS6/K0io3Kpzp4WfPWvBCf8/MPq7vgBhHoQT
8OHS5koWH0wHNZeuj6hTJASYwa4rRD/ruN7soyydbBnkUZxwQVnVYqdZdEPk8cq/Kn6d8MUqPFLM
Slg6tYIdhmbPrKrcXLp/x+NQ6mV/LvQh2q/1zXD2bcN7ELh33p7NJZoHf3FQT50AP5A2QfSWAfAL
Ev7zC3TRRXn5gk3QpsWCi2zVnmBEEDZMYbBEbt/xG0zR8TPQQvCCs+kS+6qk58I+tz4OJUin+FUI
j3zd2yG0Hg3FQ4Y1csTLEtHnq5vFoia5sBDVwEarOfwbIxttmpRULAXNzbk5Lnsd28PuJoMGEueo
w2+wXDeow0fpOOZyeVnQKe9D99jdB39Wl+90HAXYBX4RBirdb/VifoiVnsjrAhgAG20H4lVy9uAj
0jonGP+OEDZ5S/R32iRmGC84otmhLKjL/KExMHIQGGOcQlJXjhCd2wyl/3N9l9XHdhwCyiR5xBJX
Hs9Z2KO2zPG6A2V18Jhj52GgnYRweUpNCQP5dxMm+biNELbKdWVDk1DP6rl/nC9BL2iQ53KBmXpq
l0nlptZbbyQ9lnOI/Wfy77GtJQBEJfD/HG8nBNoKrKEConxiTMxqKabH4kpvykcCRG8UYJjQNl30
+8W9X21XKXILH13obh51r563WnrfVu274tWdqkZelQb3AHZcg1Ip2F229bFGRwKaFz/6VW3xdri3
nSPri53t21eZaeMIJ3+E9fQPrEc7mGd5l13A4TMFFydXNsZIJZ5H0inGamOadqz53aDULJ77+2Lz
vvk1hjNYok8mjI11K2DUdjBSp7zWcV/EgIyyoUXr8TU5s4uF87RM4aUCrZRwyz5NvhOI7oGAreF/
zN6iCv7i2FIZNNaidLgqzMHcXIt264L4J1/xAZeDqPZ8/vTN1XwjEkt/ZSrqeKfYYJu+D01p+TTP
jECKDy/zIS+Rjku7+hq/gioYxZ9VhSV3F0ZHQiYRkzGlLBKwhh9AEDeGh+EmyUBr8+V0eFcRWLef
a4x1cFQTKJJnTk/1xyDxzEdFy0fAYTKySN5w4Os97qgg6hWheHlk/An1Mc5uNg2dBJbPeNmpiyla
KeQSwzHxMZuBfyw9moBQliQqeCiCOB8x8ID8g7LII75IrvGUWrAaOYY0C0EBMXPogwuwubbiDLU8
Lsm/JdRBKxkpRxM+zxmqIKlOvbfYW+Q3oDmHyfFkNJ+UWCCpa1U/tgEL7QDjn5spZ+lAphpdkdQL
9kSaE2RA3ievmhL1DLgnpEscZkBp3xqVVAbpV4BE9DED2dT+GpJkNmIFOu0fBlhHc06vJYe4dM+1
iQrxlFbckCFZTBGYXjpS/eAdXJR/kVeIeJkP552bzbHIGjxiqvlaq+u8kwieqWyOqWRCQ+lYc7bj
MyCHlz1nfF28n4QOkddw1JhQauO8oZ69661sWUMTQUuekrBIUONHkNeYtEEM1+0UHK4rXj0HVbo2
W1ysh1gUCEJwavOE/ipmBqEOESk0LOYO7eWB+8p0B+jfCWV1iO5wq//4S0MpCQV5deKaf6oTCONP
mzf2c54aYQvUHIowNwFrTOWWloppUGJ9YbSeVjAxSaFusnQ0liQhwSqRmjfrHieW1daqn1nEDS1d
rs8iSqVw6h54/RQsXL+FrOXdfDcxsFL2KsUAOgqnWJH5mYmQXpJG0UhKT9uW1EyOVQTDu5LaVUBy
axu6r9dfFIaxujRc+zIEjph4Wc5LQg+i7ZTwprGTq9Uh3pLa2FX4nc00/qM5W6fhcbgCsr4ZV9xi
OWzUcqzD7nDNylo/Bt03Nr53/LVULCrtkCNRUJFA28UZ7A2gP9gUU1IolG4KktAEV6hWmWdwrsaL
YRJC/33m4yQHw5qJo15P8QlNbeZH4JSRmGR5l97XynSUdiHacvXMu5ic+GIh3f1LDPQu0QXfMr95
D5AooG0hTzMrB1EttDqSKw/OA5l7y7WOgDcIFpGXD6SHYC3GXh0P7mfFPIsnk6kEP8DnkCFKojOO
HnxAWActWP6hVavwtE2i2UyOAWPBOcCZsX99peCo4oSXjBbPPFIPM8Ymb+E/u/UmIROsYjiV5otp
wP+ExqKgI87Jx5ZWA0nPeGZY7LTP2JcEfpQCelQdKxYGTiwwlGbm94M1calpMCFbJGy2Me207E/I
zhvWA331fkwJeAUCFfaVEOt6xDJIhk2Pi0kBoB397V9It40/7V+t++Ch3r2oM3HTpLWt2VkEcH2N
RxIftLkj16RRW+QVjgQLfI4YMWxBRQKnvNK/gimhae0W+kyBOleRVPZkW0BWURsTDSVvNMAwngm7
299yJAs+r1u0zLEufjwgeTTgNJvTmsoepQnjZXW9kYOcgf7wxhSf9MrQ6hXgGw+lYMTCXMP3Rk5B
cOxvlYzrix1gTezncMy3OPGq5rOV9HToshtan1uvdeWkp2ZECh2HVHbHWXgW5VATy1Pp97XyMqNJ
H6+6XUwECN+NhqQ39NUV+izG2X6mjoxUDBDI1Oomxqj9zN+zqpgKYUQuBcLOTUH5DR6wDuQIdoM7
ZU2kPrkox8ZbDVdVjBZxcejGT3+E5w8h3a9koUS8DlDCgtVlFwrxvM73AoixGTVLPH3sDpDJZ1Od
eAw7n14CunPpYChYx0Jre0/EmiN8hias6kSPNNx3hbq9hP7V71C03Vu5pQSqJmXxQzBVKN8kaBM8
8fsQucEJ6RUFN/DBTJTj3RcPc3oJHertMvhKSq2yistPD1TRukmCkhoXGWYl8sdAqqnpr17ohWaQ
pc1So4R647wBS27/L4amRKx7XOz3U9WPPUPi7tgdfn3CApNy48jcuzyOqaBIfUG20QPQ+SGEt+ZF
ofLqRDZbRweCcph0hZ1wgotN2HnTrI0UlyX/2ewBziwR5zls2MrPRtQGRV1YKe5GwLqEbHWxN9cn
S+VEbYbzgcZQu50tWgEw/D8uPmrOgd/lG2NmP+9xawh5U8HciU8cWkmSD/nfJnOHrXZwrA2+hx6n
Ckpp6WCaRGT7aft+pwB4PzKF8kne8RO/GFwqFX5JP/tUE3K0xj87tskWqtbKQXWdVK+2nqNF9Div
qsEyAbsmpUgEsa6EhyDMP7VoXpkdHz6sFGE0NZXH7PCocdui3Ip5de3JgWZDYduSpaK9aTg2lcnV
1UWXJrjlrEDJnFw0JTocO0ulTYwIybXgh3Ec7mzcnIUYPkZNFExLQ/4HpQqPAjVtEWmv02AbXbDp
4Lzys8iFZB6YkQ+2iYZZCxwq1Ir/Up4XcCoZ+eWJ1AWQBbkha1ZhM1OQQzAyqu7JoBHWEcsYiwGV
kuQOFQ0kNO5s6+XyN+IDuAOx0hV9E7BLbiPcIgj7KZ2O5/riDc94AERKLktonOAQRjJGCGVfoP4R
6cNjbmv2pT1nehLriUz6L2wt9e5wtvgKxj0/VRDarcLiTlXnKfJJj4OCOPl8t66LC3N1oy5/e/lD
LvF2f0j0VXYaR3OKrD6PGYQy+NX4sN5QspwnRsyeso1nmQ+0SNj89VEPnuo/0AFVqt2EjnqHei3j
eBtuAMeUthGa602Bvg7CsVmJa41TPR8EPtDmUeRBLcmHPHT+ZNCicy+6xLyN+uf+dlu6fUWmc2eC
ruo8ZAJatj5EyqnQrMkH7pdW74FsvdRdsLndhe+aXHbXhnOBFPFzbEE0LoE4Dm78q+RvmaJNJTgZ
WadpvImcHCxmdJsZUvueWdxVF+Bw7AE5nd/Gucxe3JARsWSPYNSJuWs5kK8y9H/BhLfCmSawqFeo
DR5Y/ULHvdit2uIBgXiJjF8M0kbSmxQ/A22Jszt7UZRvudcdI76yftMu2eLZE2fxSLS7A3IwXhsP
dDlUebQ3xagqS6ABRSZBARLSRT084bOININatg0ML9EIDkVB84tp4AmJsZFS/IgUCT/L1cJpTZul
ftEECI+YOiX9XGrIlxwQwZ/C8iaHH16AbxM3LyDU5pbh8xKh8zAXj7BQnrwK9H8sqitlHMKbSFgX
0+EGUFGY2/oxSXiBYj+XRGF5DrAkaLmhx1XJiNTwseW2DQGG+FsEXOE1375kaJUdDvF0DRW0ys+4
AuwQyoO4vIergHFlz3Sen5KHFZZ6fuxkHno9GPmSyVZtsNoL7oqC5KlytkIa4rk1pKOnyzFvai10
g7jjqzBgi/GadqDeF1dbrDM8rwz6Wm0/kPxiJ8XBc90Touddoc0Z0eEbwoMvVLOZKNLS3X83UTot
SyEB834O2Hmv6nm/oOxBCcUcQtGYBV7TL7UFBtfIiErnTWyMp62dz820SgNbgmF7ZyI0ZnFbY75i
LoDChmtcu8snAL+yl49fd8O9JJ4w8coweg+A6IKWF3TYs07IRxoiGXe3RGXPnNIG6N3r8mr3Q39B
UPLKIupt1IAJF8EoVctSWOc3/2C9ojiCHflhaLt5AMJDqVh6THm4W0exExy4uhclHUi++kATL1io
2pQTWcxZz7n/KMf+3rd4XW/TpJsMZ/gMHUBOHJEfjzNB6usTTo2i1g70hpt42KaNMdEx0uyqjtG6
qtRXz8+yj3jjrf9vyIwn1Pa9o1dTrF6aRS5nojMXHlg2LLFWM/MmVvF9XRkiUbvc1lFjIUn2Eugr
dgQ7mWUCV0DcBNdhv1OIYBSNSmY3jJMLRCRqvj7USPoIOAEbC4VdhVLazlW3qIcwPmTU6y9b6d4S
sZKIggnT0eZA0I/b5UF8DfiQxcsMLz36M86bk/DJ2OTiB9N/2wIBgdch42VFSb+VKetjJX8/6Ibn
VGhj3hzBydJJJuSp1ePAFdfBTM5aSth1W06/Rpf/7/hWjzIO16FbbmgA3zX6CkFjsdk+Kns7FwEW
KCZd1ZDKrbERgNhS5iU1FB7ly72Ei4l0/OAxz2Zh7BJrsnxdStLtXB+BIIcgufTtnoGtzz3NrrLv
ul/0L1nCcDib6yY3WdwGvJpLC5E9MKe0v71b5qcVngwgsdTqUy7vxEUheEEwWIlTHg8Bn2X6kww3
A9OzO7G1s5/U/wUzeqzKjQSMuXaxkptmIcK4KySRlpKuSDnz4XuiYDSuY5CbRdNRs8XIBD6uXhKo
YZJs1SqFQw7fIxlIJAVuEOrnYKRgiyGaB73md9pRbQb+n8dRwDMfxkynrHx/dtMeOBmqk3Fl/hl0
KV3W/wwvk56rkRC63BCyOAqVA563ckFC0gWJn8PHkAEnJgPApSTTJq7ciSgczRclcDpHPchfyPg2
kXaWUIfrJ1ywGsieOqo121yHi6QSd8ggc/wcmUV1so5HE5UMgLmtjG8g3J0NVr6l831apejmsGb9
Bc9HOAVmBomS7SHVbOToQf3hEgMsXLraWK3/4uS0AzmJFSGkla3zWRIJLToGryUODEvcquThjuHi
uxVFBtOkjbRc0DuWjuuCypkUmfqB2UIkeoukSTwzyDjxGNb6KhkeBGbbvpHYgo1jUKql8rd89yk9
oSG2n6ho46Zdur1wdzl9HthWghB6J/9bwKUgFySAFYxNMyFL32IR8RPZqV0rZXGnz96X+4unO3xD
+1X0nxKUAzAqZmgYuOxvzyihk0uib6MhGPA1fw7gcCWLNzea0sAo3cscfV5UWBd4VnyK2zqliUpd
zXoyZUGbjTkEoGDzJey8/tlKfDvzzijNroVjjIP9jmS/A+DfEu79WpR9nYNy2CJbJme+lAQwAAY3
5FF1HvvIDqDgHVYhIqCOo7kHEInvhfnyX5Jlq4y2TVAvAzSQS9cpz4iTI2d0y7NkVpdJhCxqGoDu
nnLqwmEoL72+yUujsd+Wpv6v4O0nz3V/ErJAgcVcuhF7WBcQieLuiVkCdYFDhVadFLLbG3GxBe8c
G5b0av4LudEjDEg8mZ+s6DXZy4LJfVh69g10YPKdVJCt3m9WUpIeotx4zhtIRnoL1IKR630oSsI1
HN4DSgpyqIIrqoOYJTHJUtwarQk3r92D5SGYJhVW6kHq0tGvvHeTZBvBmMMvmAsVet8JMjHBvJ3/
je1Wu2wN5Bn2YDQ7BpCwJ8tzHE3V4CxpGy+vdP/90ZRDhe0mWrcwBcCv1lkdgshI488ZcEXRKulu
uKYXa+HPOXHV21nUnrdgrduW8/IYLT2ARfcqcdSm90J4k8oOC/t1j2baeSoGxxBjPVedPlzb7OkJ
3yK4aesrNYxhaCnIEBfw5/Rtr9syn3BDP6i3b44YhHU+cxXZQL6Kv5qrrURY0C0V4bSoMclaIT1n
fk/iAKBSNnkxe8bHqazYXYydA/Yzx8fxcH9F+edCWXrEIinFcHqCONof3hg7Dt1Ml8ReCcJNGBkH
a+0ZLoR8LzRS6QxcgN8f1yBR0aACRSJpwwtQnzKLpuTdgJ9aNSXSQ+keBAF6Xv1ACSVtevm3eUOI
oWOzr/MdZgSPqmvOMet8CfmTeGCDDM2G9hDRxPQQvZIsou0UAg2S2eoJwGQgp/OQIz7UIouRGwJf
ju40yyFiGs3AlRHzKOXo09zsElbz0dj3V8GFPSw6SLAjTANR0KlWy3bSVOGLSWMpDXIGIO2Fv8yw
tI14Hni2PiTO9BShpKrLFZIKbNcwEosZZuM7T/MfIaiD2nrQx1wQP240qSGJKDPUWwpV2mOmafVv
RpXlmOneCtB96Uhe/qd2JLFHQ1yLP4jPyIcEfXGFKJOsjKZb7auOWw5w6T9zRcsqJKjCHBG7XoFM
QAG0fNHNjEor/SyKXdq5HKKthH0VuT9t6zgLKpzdGZPhu0J97n2BI22kdZLrFHuzzSuquSpG2fIL
mV+jZJCTclt/bU/l1oErGJFgFneNnD/gjG0r7IpC99vfA+NvZ6XfSujL94Nqzk/FSDWlgFMgC/xj
8xDNP/xGg5tQe2852t5AVXW2smCsF1PBs4+KcvOAJOpeKQ+FHw4N1aayOn8NtkkreRTop6unn/a0
PvTmxGauhqe7tM28V7vkoBH5XaZJ7d25lqC6LQL+b4Qa2jOcYLbrBgVXNJLC5PqSm+sDUkHeufQx
YGueJbl9rvZJj9pMwoOmQgCKd49Q/afVlM48E3m19Co1jzQdz3qmJcHbUiLS297Kj6I0g8G8/Dat
mUrNAG3HyTiIXDqFxSBWdnQIJYbPm6JS5WhuIlCZBVvpQXVWRWpOnKJ/oUpmAIigbXkiazhtXu3C
ErH1E2F1n2iMvatnw0GJU6pKpnTZhWnymMsO0M651v+PX4P9M8zZsUrjyjQxd5WFpuf8oVMql/DQ
pQC/wc2Jz15GyrJvfeE+xkpQFaykkl80VfH+4gjdkY8F9qksDZV5s5E+bV3uruogjW3kZynnuZ12
2YpBi7Z2VHnvdZ0ihUVhwwSiC+PtJv+59eQZS+OeQwiocLM9KKo3HqyAYhkmc5cJ7310IJGwMJvA
V5GSx/9z3n72jmXTbO89REC1kCTQSobv9I77Y+cY50nBnj770v4zHtMmB1T4mWy7ZsOxbNUaMnFK
f3euiZb6vKZ1aT9HySqMVaD7MvZEoRd4gRkLKvLeih3kG/PaE1qD0JDrtzcOPDvF8Rz12SV2LKE2
rnBon/5+D7iSUD6KPEN6CdimiZ4aQs/CyBbvpY1fDIjQ3U83k+zaZLJgZccT+yRw9RrG87qn3FO0
nZoop16MWcZi5fop7VTmzhDMJPMvJQFEji1/v9qzGNKUTJ+y6zEvYjOY4tm9yzl/o1cbBCICWjZF
AbgHTyXIaOhcFXTMp8z86dtkdCzg4k9DneSafgn7P2Jzebe+TWSZTubLsBhUtI3SUsg8wqgMHH5k
iPfeIf6oIpxKV4j8+m7UQ989zMF72pbqaculpOqpuq+O6+8ZFBT717Qccmfghw1WjLLuWjAffrIj
IrQuWGKxVyFSmuBwj21bkPElcaN1NxC4lKX3vG+5B0e7/IyCnGbWXlR+3Brf2Fi6HDVC1eylkvqo
5+Eu6ktwFGNpH9yFEeeLKJAbEKm9p5EdnYlaV8szDA986GFNsWWGiTUDuCxmCWYf+duejbjioKSb
6MPEx4eMJJekNVbfQgYilDyARnl6SXJuootCBNhUddLlypAxc26q9XISh4OXLpgLzbeP8wRPp4tf
Q0ICrYpcCoSW62bBQnc48WGuun+ZIVxNCQdEiM7aoFPQKWqxXjmcNYjjfLpMdScCpx32jLO5ZgYN
x5sXU2s8Sb7kYW1Ti3cP2uRlRGWhLYo8Hb6aWwFMrDgtIgtU3ejEbLJ1kpGZ1C6ObY+rsGsfgvTI
fUxpnjruCKe0XzdExrGBQ2FK6yHhIS15BhA662cCvrf08D4QsQ/slzuwuUgaPlPhySzRD3z34CG8
xADCDtK7eKBIc2bgBYJj2pL9mLIxnMjSVxpOS+vRxPRAtjAQB9idhawMjpeXNK4HEQI3+4PJNDLC
srimsap3jScEnZG1xxxVKoxb1ozDO+mMzKMPSZ1lEzPCqur16kz8aEu46H0vIjph6Ju1xBYGgZQC
WNXFvAstN8DICWV9AWu5h7D/BN+ZiffHtnz2VoFYuCJQd4LldMK9h/poimjgY5G9wEbZQENBG/q8
chBFh3eCtaElBAp5O8lcOmMj5Z7sdypbyagt2swGy70/7qvp/4sAcz+H8MvdpJIKKTx7gFFmj5pf
syABHe0AA1BA9oJ7ghNEfCAQ/vlNBIYf2nEXdryII/gRECJPBu+Tu/G4xbWs+IGjOXJXsD7jO86m
sYuoMzPwD9rpPgRucF1dyxMDoryDPN7Xh+QlmJAzDUA7ubEsjSv4lkt1ElkRH4AkUJbEI94e+k4G
9J7qgmBoA576iwxThSGLXfqxKLvs3asBvsMvdhvHoTaVPTT520dqHNNa/YGVTHv/qryHrkC6La6o
LUUm8/vyjotSYVyj0IpWFnwFg8E04qoA+55Lc2TE2uCNXez5IG2panqDy1NHI0uhkjd8gowURvMx
aJoe4LKwZ0aKKYgZvQgU6rm5Ru0Is5F6mtPNnX5l4YbuhnCq8t/2JG6LTOQGLlI8f/0PjaW8r3h8
8wiyrPKInYPNb3J+qr5qOL4ocR8RctunqpKIBte866pzjeMX5izG+SDp2GdgXRCGrvptWTEBRtL2
F1VFOyD6w1qIT/7wfbWRnQjGrZTKe16kke54bH5yQ2WbIHqAcdC1LsNB3+2Qn2IeamqkjG8NzW+A
nfJIJTgpXS7gLp61N6LVeV5y1jU8pfIRV53CgLWrYW9sHvjRYAVGR7lP+vvfCMSWrkaU0yGZ6P4j
gA2ZJt9N9CALZtgJVl/9wXFra0m0hDoNyypj4XJTLy3nJ6DG0CYu/ixVkXcOz+kPJMFZQaGwxo2z
hVPVA6v3mO7h4LoSJ+qnsXC37uE002CJNbU80AYJYqWY9cuBeHkV0sH3JLZn7stGH1Vd8kTXk5Nf
Owj+Jdg/Kumwwdf4jJw7fruaBuBoc0ZsQQr/xZvyR2P7AN9fK7UPpeVsENn2zON2D89tL+LtaeJn
KHO5UPAjP3CX9qTiedArI3lwelKsvcbS/9mXtyhUHlLXVUxFwhquQizrgVbeqhykPD4iqTJR6i+5
qABVieHol2W0dE2t9wXh+QYU+f5KvYzqwe5Wu5yDTyXoDdsRNasxiwYd6kxC3kt5Z3k5dzQBWBW8
iizvrFnxARJiJOwrfFztUdq4pqAllHTFH/tUlpK9Harp2y7dUW5VCCStZLCfVpAtAuB+DTPRcfsQ
+9qntO+tZtxlXUaQ43TpLMS7sJ9EN/ytnVjo+Wy4u8AUKgoPNyDnn9bSjB+RDc37l4OB6Al7GO63
DGLG102+ggzWq67ifjGY1W/XAjlzNRjvaZTkSpmGgtvJNvyQZMJ0HjV7t6siyGvL6JmeXP9d6B/M
6PRr6UTSNilh7HO0Gf7iiwtakexFqbStajWvEgU+4H6z2Eeeax7i/ZA7gNrmjIYnKKXhrHhfcYHY
Wco186Be+nrEshFr2RELrMwbzZrvjA+qIRg2ETBNTCDkqhsHGt7WlUqbAmiuguI1e6Ki1JKwZWop
1DTly5Uq4zJfxHqK67LeGfv/eYYtUGjxnqdpYjiwtk4L9T7nDaNQl2YitmMIpMviKWuIXOiZMmR7
qfyeuM+CM6JW+uN1+QdgEXgbcwY1w5wh6g0Pz5lbJqpmtOtVtVFrjp33efdj8W24HCaIfLFCbmwj
xLpONOnx/wDHqi6uPmD/6EuocKFCkHaL022wDKMeyDgdukSnr2p8bcY3nw3oIJra9hK6m9y/WMpU
Sl3o3UxEWb3dmHzZXueJK33Bx6mg//G/VadaRMpt5jmjl/L7qeRDyNkCiMBJhrU5KdYlqCj7Vuq+
AtSAOKJm8Mi43HieckSga4dWmRxgwhhMnO5G5VjII8buZ3Y5NT02mJo9LhsabfJhEV9EJwFC/LKW
kKO40QN/1U8lPR8o15V/YYYnhfiX63NnQ8vQQAM3HwYJUY4HTnLDZ9ui1P6F0kHW+/3qOjwr4Nws
qUXwrLFMoSk3IcAY5gRM0X+7NRm3puNCNw7UGKcP+keZmGHXgHBO2yQeyVrxLdTS+J0uqSTadUix
yE6DJw3zI1amtlLGbD/K+lemJ12VA68UTQkkO+hisuO1RKVgemGx8fxhksMti4b9x+O6p/x3U5ae
f0yI9ikCYlod/JpJhAuC/itGHG3nGsps6g8DEeNb/PdlAbH3WW7WD/V20i191nVpUTtioILvxd0S
V4ytWuKiz06r1tVD1t68VyUt16hEaBeunYQKPnSRBfy6mEBYnrYxXoZRF8mFS4jyx71BOMU41115
X8c5wFO7pYLcCAoSnXJj5+iPJ49sy2QomGz0PIOSe5t95rhlcN3dGxAKmE9FfJnN0QKgGKFDYaQe
Yt525RMx7f9NLhR9J0u3A47Pf6nMzLHRrRYUmPC+N2rZzXcxAY9ra0kcQLnNjBiI8XuGfy22ZNAA
octnou3GKvVKdXQ/fx6/8j2hDHk7fAwGuRwWsiS8VwYkkjU9gBSvRerMxie4ytvtUGa7sSHp6Yva
DtfHae6fc+S/gjG2kh9vZezwNnJE/KXeTUyBPEdeLSNuM2gLxspqQJFStut7tLJgq1hMAXZ4SmSo
o9QJ7rZN7+ZAcH6Ur4mDVv0lLW2L8XU+ziCA7id4pCqTz8/j0V7IvI6HHsi7UQhpQkARaOZ4rdUC
8U3so0Mfx7ldxAK5mo/3kwNHS6ZugsQiydNPV+nT1FwRHRt5taoKHbyVUjBoKLQ5OnS1aDX1QyGY
+wVz37KR5EOQJpDyTVWlh6hi5K1tQqMGbYe3Vpfd4oragn1yFc7tZz/cISxHnjnMCzBX2zbrv2nu
jOoBxfOuYazHa6ey5w9sWJ0vixGQ6z2pM7/c0hHKA3wWOggV9gu/Le6y6BHgaGfNxHlnJlpVlbEh
u8MaY2E82qMP1fk7eUwskGIjCtj2JpjhVt0dONbpFSJQwM1IhF1b/ULg0BEuQvH0yRiuWQfH/Vu0
PZlOHJ5e2P0FWDKE4dgRIHm03z06FoYzaOgnoEexaYFtH3CIaKueDOF9VFSZrpk8ZQNCi/spvZ90
JlEGocjuZlzbPP6Vc6r4jQgvKQpN3b+0BvENFoN1W/ju0xGoDU1R15A81gMWvCTz1+i4jUBMlXM3
fS9JUCDWRJYxqcz1Dq2Ys0c1ddePhAy7sVPrp2NrRiHIlJPwzJI9NjSgNMo6oOY99jiZsd+jaeSx
Tr5Oy3q2m6+69r8hnz692ihVOXYVLm7aJFLzE52FJPr6zgU/PL8idx6PIAG3pbE42wWM4n0fjNmI
CH2vw/ocvorU3GcEQATKivl2dloVaDK+oRqVC0KCnNXZN50OQ304en6heh9wMNGPqKOMiZOPPnu2
yl/sH91uBGMy6YUJ2hfY711ufzXlflHoB0gqOcFDg4HTGTmecUEZOvzOXcKIUinH8GY7T39jWrRK
Abx3aitFyQ/9627z0dg94rj+P3Ni8YjAqHU5H9ymTNdw683xSnfom+GhGAohxwQbEoOPPBadkj09
6FdKWRmskJd8OIZf2f6bl0rlnrHkNpq0pboJrFQMDK/qVzYa5mlM5+Uz0eZCEw6XjINlnOOkqpie
0x0MVB+uZRNPK+h5Oezd6oPTIsdICjLdQLqTRERjLKSDJ9suDIDiHRijoU+Edbm4Rs/o50ieOUjB
SUT2P7P0K8z3tWytaXZjPNMxmNx4sUrNmhkhVXvBiwiLhx8IUpJNG30+4kDHj60v3Tj1l93Kue0M
KDwf5mjyOsT5A+j6dZmL7YFCfYnnVmD1Xb82DuJ3rjxTrUJ9IdsFfpRqoPEkPfxflXhn94lbufhs
rDCoroXsmVDpyoTcR8pkZGMj9B2/ZlcI/RWXk1cFRSAwC4IkU9wAlmhYqcVTxvB/Y0UiUU4yVfex
fXFk4Z1YnvEDAEOLkxd7dynCzrufZ08DwrJRTy2gSAXplbVulbv17NAH1/5JW1gUvqeTwlUJfgRv
Mpj9LpXloCHTx10SDFz10Id8oTRcjwsYbPXKQPr5lX/7no7eBuvcX9j6gm7mHVJJ7dPrsvOxG+IH
8PdUszsudMd+a/ELJD24cr+wH4QNKt1VFcUyr3cTNbKxHgI31KM3nk9baM+4jZUu8Ac7nnIqqGD8
kbT0c+MrQPktkm7ZLAzEqakFqibMefOqvfqZA4+HbgEB4hKBUUaRJyeZSg049Z6cj/Mbc5BYanIL
uwt8N58yUea6as09gG54kDKeje9CVOVTnYZVa7fcTrSN5QikYRTMvbUAASWahw05T5BUYcnm0EqR
MhZV30uA/hDEhTOyzaTapQgEiqaZCDAu6x6to8WqTlhnD09nJLfVQ4oD2ECD3d2ga8XYcf3ayIzI
k4yjsC77SelzX+tLfH1xbTwSd4vQEb8BFOdvjMf6WzsSR+pRgdu9vlMqZADfxoYtldH+KphOrQux
i69HdCD5c6KMU/F23fSzSP+AdqkGiYJoMk+gL3bWMS0BVniPznJ6Jnqd2+0L3aSVaGUQXcrwwNaD
BdyVhB2ELMeS8H5nAADZIPnJ7A8tJn9m0a8quvVQFVbQEFnNyWdOjl/BnbruYk6KI4ln6T9IewyO
EO6T8Tugcd5ZDXEyt2dJDImukwSn3/56pRQ9F7glAXzN+IUOIou1IaixGNtEa5NS8dfFn9Bx5pmc
JD9x4opUk8nHNgW4azzZmdNt4I+Qw9r+uoC10Yd/ZcI/qkUGZc5mZyii2JJiCmahv3t9vAiaQsLb
FJLzWP54IfASH+ETlSPQnH/dptJVqL0+WXhWRjw5v7JJechqFJuS4zHJQ3WqJLLvXJsu7MSRKG6e
kjqYJNmkvuivtIUFbmGPE45i4RajrlbROZUuKCM1GQEcwHANtZCgHCnfB5lmdHvak+oN6gfNUnIS
EYnxF1PY/siaY/QSNuZCAHbwQgr2E0qVz8eDV/PkFb9pIdnlEadoI9J4+iWt7solaDCCJVmYs/Yf
z/63J1cOCtpPbuEsJItxq7DTsJIt1+bpliz2p68vJI2NpyjVvWMfm7YWcoSujzgVpYDpZxbMrEIq
1nrWJ8iiQGrouPV58Xa314o0sxClr/5lP7tapxFfGer/BoUDpR3zVM2CKP+RXe8lfD6jxp9FtQEa
OpzCfzcVS9c0aKubG9FrO2gqLvm2y58dZm5YmkcxlHg84nJxaZeWFtrkszDZDsPdXN+6umInmdjj
D4c7BxO4oO5uldmhrV/LkFPQbuhzT7SoFye6a2f8guYRcZjTxgyfzW4UFib82tlusbR/uf6iH8iH
KhvU7UEwfzfy6ojc2/zY9dhoFlZVFRqjW6NFlT1FsaLxHHFyzszWOoMskZONG8CQlDrpCu6K/W+B
UvJXSt9dBoeOFWMv3vfYqY+p6qlappGERjWLWsnEEn5XRTZkJ8Ym/N/NMlTv9PPXca3Grfc/SiRS
QkRPzQVuDxGNVjh9ntkBV900bgkIXNUOFTdLkGOzV5eV3jAmNJC5pm4MDfLjNRdumT/s4XcIuJid
ph9XK/IVvNuYoysJiSq/zRus0ti+j7lJH2vi+Ag/kbTPuAY83QUofOTFN+/DZmmcdl+Y/69tq4tf
p+oxagUDS6zmApAOBQ5uN5zMtdvj3iopE4XluZyG4Q4HpyQYxfGrRn6dgqQO6h6N73xhqzLy+Kk4
tD2z8AAfY0MX8t0cZtuyo/NsV/OSkfbtid5NyuQ3CUWjuURX/vhE1/xTTBxhDDvtcJl3TyVnlrLD
esT/wzk4hzq4LMSOUIfv2O44h/IUPnyKMGJthO9UBMt1cW1QLxNqlNGAfk2w+gEllSavuiRZ6ui+
arEutzMJtgwXZWrjTen4HJYtmiKNBdepDfkHs6s6IDEmGw3nHvxjAtT9aHvGYA6NMYTjCIy4RGUP
ckGgf+cTBfOTW8ZVyA5UcsbTeye+QN/DIj/u6B/dPZSjRkukZsv9bJa3eudfY0FdOFtHR9R22z4N
K+haNJQ/LIeh5MQo/1moMfDgiZbomAaLenwzvGK2Z+n2cbC6UxvMY/7xwRTnVVWqaQCPY4PJqxJ3
TP08f6CDlS/mmknXLaWfkTiS9h/w0/CBJ9/rXMhNxILSN/gbWG/MHHIpgt5SJBDZfLdsAhjq4xM8
/M6q46KdQuhbG+yESzMn+kMS98cmS2bpBcF76zQB+CRW4k5vZQbnW7cEsGQQY0xp+Vts2D/rIgru
/y/f91Xja/8xvIu46d7C9XjQcl5to0MQaMtSm84dHn8adTBXn4Hm+OA3q8dr6V+UUZI4H8y/dH6A
q/zzGZFSA7QiqdOZC0dAbk3lYkos2z6XwQjCCr7FX3s6+eiPJ4fUsIu106UqFEeXOmfIjS1XTXdg
qzzd7aY1xp/yAm0reTt7JvQSTqootGW5gLl0UP8D50PVVgSu2IqxoQBJEsNprWk3ovEWvcSfvGyG
SzEhBFwkQ/BoYv8i6rhQAPiHEAz/aVDTHZ5Vsam26+EMXF6+TVtiSdIIwfvJonIUFxmOTx7DsijH
w+uRv7wTVSm6sWuPzlC9NxrU+S72CP3G6TaE2gxfR8Zgp/VWnLWMbv8ZMzFo1MudAB5bhrfJb2Kg
dmPE8jG2ztVWPy4oXJOde6KNiXA98r1a1vM/6vYFC7c436hBJAvNcSDcdKU8MMh/D9MwZnAmRYDp
kw3vMscYOe6LbRrQwklnRkoHzLmD3J47c9QdClq+TqyHRYudAdwbcoAlLF3cFQBuKLpc9l4sETL2
/7EYs1ci1MFmIVEk/5kRKvXPfbLyd6DuicdZouF3SWbVIQYRCMweUgvk4LPzLgBeRv/EFnPFbR2P
msXymXHNCupk7LTmDyvCmhZJR+QKC/vsBmvCRBW81jQR8mX44g3ZiZKq1L4mfhEXyaLU9dGQJ9Ft
nFavwxSpVA6RPMGkcLuMxmg5GRzhjgO8O38aZTceHyXhaNLaj9Xgp1oJdUmPAiTly55N+tc5hC25
28BycJFCuoidbO4b3rvaq/HAOQ/V1ot4FSFbHmiYY9WpNGgQWuxQePEvy7E6WXQGk/+969nr6CXP
cxvExcgY4rUeNI702lWdwauXyfOe4h0nWNLxwQkyeUrFd0Ljvl06wnc6L7VJ0lJe/qqkR7pHS/lZ
6flx3KH5/JPCqnQKlgWcASGH4iF9ILadcU0ROz83uwXap8yS3teSS/A5NpJ2Dp9h0XpOhA49VIaT
y4p4pX1+e1gz4/8Pc1Z8LeiRYXlkwN/vtO9AOln/7xdi4K+zdav9QgRTmeD7Vu+YPdDFFNkAQgLf
AUZorH0KJ96kLX6SKz8Jooy9WrBstryzyqcX5gQwBfk7tRmJRQFN005QkJOnp+vSqVS5k4R04scC
562ctApODMhPC1szq164GOHimNef1z2X/UhS5X7uyfF/EpaKgKhXbJADp9JoiH2B35EFxmKyBish
eRUkahtql9s+BqEFLKwkJMwlBnbsZyo2DxireQKy0tIqkNc9FNtGQouLqLxscLLxPPRDiQyMiw1i
1UQttqmR71M1R5F+uUE7dyhieT5dBd6C8TVo5TIf5u6R/HMlQJllNmrtYNfOr5xvSr8IpCHpopBQ
65wn1CwMR+H7e3F2xN9LFK5f8uu1UM0UjDgypYGpm0G1Y9ap/2bA8Z0Psr/zoyYTW/nPsy0c7OgT
meFbIqaPkrSTr9HjQOHVTFfWoewXZuuXs/7DfDzeSLnzyAdmmJ5QBf5ueYFbf5s1mQIsMMg5EbMK
S8HbwhJdG2HbTqGkVG8cCmo+lEBB29eurT1Tfz6W9wzqiA94m7nJbt9gBsC6YiBhrV040Y47DS3P
Kpvpisl/4yM6pu8Y6gN2e3GF8ZC63GS0ELL9tz7rFaj3/Zn/2bZwiX+XtWdRazgvjHYD37SRlDBH
dXAS0+TVuk2iH9iQdGhUMlqQI6RY6KxY5u9awQZgimzfvZy4FRb5eZ+MgiIViMrDpjZeY2jYmtU3
dAZc6g4yG0MbMTOiUQvQiAGpqJANTe4oj6lJLHZLahbGSo4RGHGQE8OeSfJWjxs7YJLvnXkQwKMO
KtM/HKOt//QgSAUT81Ri6UPSMe/SNnNPrmt5yTKZt9H2uJV9mJQ0qrc3TVZt12Inym2YgfpDLP2W
V9VpnEiVrmmJaTPezBeXz6mQdoqU+f388Ul0XwlE1i0SE9n+cDnD4gVGFE90vFVsu9Yp2XISkTA6
OaDEWNk15gFczyBzN8mC+pjwSTzQ3tmwzb5Efc43HSPP8W8l7kkVEJxoiruA5qta9wYI+ERiBRlx
/y0F5C6DLnLqs6dSrDovfZzJACmlsaWvMfUvCAXB5eUIHY1Y/92rs63zeg/gmhwn8eHAkSmRaiJ+
GQDsvI/3RJIlm1kKu0zzSrOv1BT2coy0Q6D+Owl2+3x3Z9z3JosZPpcmVVUcXaHcaT3CbZ/TY/xJ
s3bXWSp9UuwnsNUSn1cqSDPIpHXQwWzXj76KUeCuYXB6nbU8nggcrIK5GSUvhYFShzXhpXiB7d0a
cd0oo60V0Jfvov+MZb8I+cH53k9gWZ6l0qoNqnZC0qabJrVf+spMeWpVZpmCWs/AkOjJIMJCI0IY
FFz2pruViOHMO3hL7wc8e3bo9qaTqsSnxn+7WkEgKjSGgzgG3hiXZQaOV/eB0Gg/hqZMjhxZuMGv
+X3g9f0LzQU8m1hD7Yez0KiHUswZiaVGHBgoKKtQshHkyUplucrk+9eF75OOzcxaA9EPnBnUb+54
n8RzcLu4xm/3DwTE0ofIIPoCGW1Neywm18Jmjd4KJL2/66ieABe5K2rjECEnn89NtmGPRUM6s7Ve
rdAVqm3AuZD6prLzqvhbhiHVQkR9tMfjvX9Nrwa2yCC7V497KlnyNiofvzET4TEFdUrW3K/N2pjO
OzhbVZhNV55nrZ5Dylwgl/EryFAd54+5O+JGtKDBFDGqWhisFHErIISvZl19mRIV7a/C39b4JE29
iRtQteUQuV6LzRvIsCPZMAf1FmtpMD5+eHo5slZhwQVgu7tNCHZiZico5qTjATQAhFT6p3QpWQXO
pdm5LxlFTndXyyLnwVReJK2I705lqU/YnPn0014mZ09AzD2i3UmQ7O3qbVCLZxRkL5OPU7GI3FxB
MWf/0kxYsTRHQsVubo8GLXYQpKJdjwMUujk5aijNqybZXZcRT9U418VUQyRyiaeNKV60DTrFtzrU
nJ8fBUEvwFPJt8n5J1XgERX4XGv4WlcMu82YLCr4az4Yk6zEU3iIgfXJadopYluNrDg1tlQrlbVY
mfxtf2R1UeDRNf853FgKzXfcL3io2/5sIT5LtTyJFQkIdpwl/g/LyjCBDArxeUWWsx2V5lB7xtUl
74sMJ18Up9ATJ4WBrWTwznXo0IJvQAhvH1Fs4DMBaUU5uiL7XkEN4tZ+c9+hH3hQKBvVQbSiePMi
jssW/OjmwbbT34BiL4pGQzK5rwSRUwTjtghCaiu7hPHChrD3gLDie9kD6O6mGudzYFCday/Mslpl
A+aQ5ZFZumrTMUos8E9aNiqepaBh0NYzQXY6bhd0IAJLxCMJSOGQGpPMQV/iwc4S+R3DxZDiR2RM
FNBy4MaZScK1uURVd7iwXer/VGbg0uBo1LdcOLZo6CpB8C2xWZek6BWBlS7f7Td6+hlJTfEh5F1v
EeNuOLH/50KhnkjX9OyicQWC2HwQ7O+EB+63UYj2FZP9EB0Rjf2PDLv31hnAk6B46VUXWBK0puLH
eDZJtkCxfIjX3mND6FZdzDfAZ2GiQz73G6QtqEm1WuGht2KSzqpxGYfB2Ve0bql9dWSHy/lD04z7
ioxNKy/twWF7PrSnEP3DEi2/5fYutVsBpKcKugcdB64K8wsCXDm8xDqsLgWEOG5R1Bcg6YoDyu47
4cS6Lv48qixqSb8Yg6wsNVH6PkxaqCGaMKPOPbR6/w/3IjXdxKPhO0M7l5ivh5jdNlGmco8zplvp
h5xGA8pIBr1j+e/w5zIQ7ZATp7dk9QyU+3gZyavVngX2ZRv8tGYIscpKuT/AVfrUYccGM3j9NXL2
JzSaE8GOHI8Gho0UwsIGfWHHuZi7IoBDe0pCAFjLg2hp3RSIJ8ciqTk0++d+qn182hV+RSU8DZfK
i6cKPhDKj9t/vMA1aBAYDriZKogQHIqDBZB6hyuq61PmzNuHjSwmHk0fmvDyhzu2+6boyfGcjVnX
qtAHUKlrTJXDMXvg9z56lLJSY8XOwsXPLqvLPH5Zs4NFeqa8c12mLsQGB24h72yOAfQp8XiqN6sK
LUzRnf6w1cZ/109fJcP8o1Eqf6Mb7r9S01wCwL1dmzXofFbBG3ilyDG4HGnIoR+XjnsOBF1rO9RQ
rdYfJyn3rE/h5mYwUcMm/8LMqCW9mvXMKFUNmHFcLdvD9ySo9oEk+wnLrpvQDIBbVqZ0yo2nv4Ho
vwl5cRZl4qpOtLEn+7v/cwhh8uVLsn2S51lWpSd/moYthLcF8prb5UCZr2QuU++wQX8ZccAyy1ue
o/dqyi36/OGkZRRRNmCUbCBuYpZfod7ne+9pZ4oMaILEX5gMqtmkicnrfR63DvB5oFIj4ulSWx2V
N0snDltcccC7CNKg71h5l7ofbVcw+sb+bY2TUFWuI4eQCkNYCtV0n0pdQ9ikVNY5du1Qk4kj9Z0K
Uzdyr2pD4nZyoPJ6KzqcBngbYQ1/kdeeVObjz5tw9BNh0KzIEmYgI8aibXP4E8b1kiyaxv1HFx1I
6SXYmtn5wPoUDH7EAyOgoXnZYoNbLu6toNvY9HNcuHBfFoHA8wZ6ccUML4IaelxT6HF+e9GX8IkZ
H6iZIxjKt6fadOCMwqEL+JgTaOVyFw2+oXoJaep1P0PH6QAL3FC9jgWYWn6JIQeMza/QrwPBGNso
dsaictyfGKmsfO0GLqnq0WyzROgq5xjJ51bD00w+8lsKQLY+6Dd7v4TfVS5bxklG4znVRnEVBaMf
MIYtxssG8ytQGoW74AMqr799ShpYrVi/KlTwGvrbn4EYfZej4BSji8a19rv/t2cvhi2a3EZBv8M8
dppBh7Nnq+taH+Ak5N3StkXuyfh1aarzrzQce8VWlrFlPc0DYB6tIEoyJliU0QP9Ba3sLTMmwV25
FL+wasslwujo4QL7AR94o/5lytz+OSu4YRCKqHVannL0Ngfq8jkGT2X5WzT6+jTiV+WU7wg7tPqN
VHdHRrbq/216yw/D0KzrhQ9MaNN0YC13xV2l+A9lrp5v7vchoc8icA+oqY+9XARbHyOsCQb79wTB
uXgO3UEZv7CXkvOBMqN5JHh7pJoN7Y0K8pTNqAws/Tm3eJSrgpDUZtmJw+ic9Iokd1engu3fTuXj
im5ssfKD+2dySyLLLTi05O70Z0zYFJsSdiD/erSWnmnXjngQTjhB2KwvUqdUmvRmVV7CagX5QOlB
MVwm/kn+2EzKoVhliNCVVzuPKeB1vk/tHku7ilEDj941ic1GU1jJDOh6C+uL5TbsLnlD5bRhBWWc
dGJAGZoCbBdIoT2J+201iakW4xB3szRHlSy5+oGstIy9l7c9YdK2TNZNj2gMiTIo0mG/Xb0BXHet
Za6yy0ldp843gW1cjd3o5MMYAvdrIZ/4Uf6DybH2lPkFxIz5mMLk20PViXGF0hZwwiBMXgEaV1Uw
qVGipdCTeWNgiO7d51R58c1KYq9kz21UMr+Qd0WpLjVOel7Ek9RtEau67sHGZfi85ushFfJxlRiB
DldkoS1S7hp52mbgKgWcfLTWhb/sVKG0vEOY17pDXuUrciTs9FfINp6sZLJ69AW1stPMP9yASZX+
+QCDJ57xGQuXPNLXuFlyLkyFgoPmRTC2sBAItUR0wl56fyd2PxSogeElm/dkLLfLxj9EI/8/OyoZ
qkOyx0mD80MZJTFhkAQ+P6clMM4XEy2J6Cv7qOuUxYOa8V2yOTtS0Xs5oBukzJCQjzezY3D8uLjj
3Cft8jDyn6gjn4Em2GpnnsArVR6l579ovFS5Z19I0DgNG2Z9iyrhxhvMzL0lejN9ikyptPA//v9f
4DEYOWUsiLCIocBrX1jZQqUyK/jUa5fP3I9+NePiS7Wnv/C7hYK1WlE7GaEsGN79NvoON8MNfiCC
flqs+xojtdIyMbW2dh/ULge1guNfMxbd2zTkIlYY16Q8UcOgAGhGw41QM2LoBPN8Ui0JT3BbWTOj
SCcWfDT2V+vuA66U3dPToGC1R8uAf2Z2Q31IY2AZt1OO8xDI9GCgSLNQuyEyc56bnHilwIXyKTkP
85MMcYhfLhZrCSyR1MF5ewRyJg2kJ2td/2De3rBMdfrKj6c1SadTZ/9KAztLmKRBIW4RlsMEEnTn
yQpTeiR2MAhAdc8Hgd0adbZbvPMujqlx7Njl2D1PeEynSbhOKUcOrQFv0Ur4ts0MWrq871L2cVEI
EzhlYCGc/KgYO8t5Zh9MuawPa+8CeytLM0LI4uPiKAcZk83A+1w/aDDMCPhNlAgOTO6eQKolnI3/
DLR0bcTvgprbZmE/vC0v/xsIkZ462+ADw9Qs2ZIW5N72KGFZbDs16JCs42w4teDqw3W5NRmaUh9v
uwxOKm3yorkuVF1z1G1FBhW8ZuTViJrHDyggmzRY1VQ8GsHVMz/H3hrx41/dL+IZaLFBsmhTdnwM
v8ULmuAytCqckXCrtgR3/bO4dOda6o6Sqz2HfsbSBHws5DZ8gZ19mVxfrPlD4VSVDEEzCO1s4Vqp
8TlXVx2TeQmDjYLwt0GXYSkSsdG1NLzT0LCb+odZmsP9KIb3UoUUmJ4tePV2DbXvmKKGkMMqEqby
1FOHFEFU7u5rUCRqHBBGMTW/JJ+tOXCW9EDrtj/oqYTpnTlxnWBhI017pEVzDX1zBm94YFsMFd+d
mfj3hNJgar0Py6TB+RebyNvw0ict0lTOBO8tM5fkGOGPv2ulKQJJE0ftOsgsIQPiv5dKR7cSoA6g
tyxHlIKGMboyFb4br8xJaOFvMHrzAW3L5JJV2hIg03K39d700esu25Aq4zFyyLPPqTK2HYNHDNXf
E2PoMu4j9/aF0kWKN1phYHmrMg673GUg2LuJrJFbn2NfV6LoQIavocHOqrkovyfsXy+yT/SkXsNE
X4Va1Vpa2JThoenNNJDtaXD8N1wP344aLYOeyo2DTQfbW5yHLCrMzs/4gKnV23z6FJH5MtcVZG8i
L5upXNqBU0QIgbjH+QNWiSfB4kN7Huv6L33bom+70vnDkEyl3IRclYms7DFwwX+Ac05rvaLj9WjI
/WJZIlBaJNrZ1ULjoTMl7NlOhgaOEGa8amZn9k5J5sU1HMfw7PSFGoZ9fle6ltcpwR3CKgwKoX8h
i7kobtM91ZgtdPrtb5QBkx/ABGd2ddiaXHRPrXJ/b08c4JrDU/Na3dzLEH1qqVm0w+BnRVwbF5hX
SeOAU9v5HnyHgH/uG88pR1RfKlFePl5/+QoCM+euQqiS3PoDjqdaLv2StepdbCalEjDziu71rGGK
CQK8XoVt000pUP7uZRoEF78sYknfDqYGPqw/s3URcTHVt/QSts8O2RFCNnB/c7Akq4xsB8P+7MAw
wGC9MT7zfNrFkCErr098J7IvkHWF5JbErv8Wb72QW58d1kIXFyMxNcrUtaiCLq5xnMxk537kX7+M
azYLXqIonDYAu5ChoU/nZvyC7niHfnsVJCWIP5PDBKwNKogw+R+ZUp6ZnEKTdVUqauC6LcZMnsij
Tiz2cPstkkczeMKWTODVsz0AS2CWnJHQkC2hFMjWsEy2yBzC1csjrAMBkIsxs10vfe0dJ1CMzZ3R
j/ycMa3fS2tzfU6Oe7WbdkigloVJflaT5uXBCT1wuVpVT3efAdQeZWT0DOBcXXcZL9iLQcxj5Y9/
ViwzJ1CopYb6mEKroac7/wXHmK0m2rgq+lbCIDTr7/F6R2B75dO+HM0kkBCQt7Ptynu5DL/ItA8D
kD6XCs7npzYLmhh4ew9966p65mpYopvgexnPflubzmyxsfJ9r4KKT8EOXQUqlK4qbowqbnIKnjgx
CKNqGXZR7Y5CWkVgKhqLYQhgn5bC1YMu+6NORb2UZZ79aBGTCFmYMEomZ1wp27ymXgt5PQDYbGxN
3JpHPqY5KWJ2QgtdR1qG+9MjXtiA6sdfALeqMhPZ7RJGGRi/fGw4/Ti8f9A6Zo+7X4ts8DoHp6aZ
o53WH/xCUS1m1EuPpnCdCg/KngVC5Hwo3oKBICRAMCIBo2IgQ0Glwys1T7QG6NH9qL5d1wAGZ4kU
leO8XHm29gwL/f480f3NWiiam40V57aLXkl/F4VOReR/Pdm2Jtx7F7TuQcF1eoxGSheqzoOsV9gg
xNBvBQwFTqbppY0jYR6PDDi7DB8hBfRmnK8uyeg5TkgN8t+A6EZVqryLYt0LqBE175cwTEHmyFoB
Kb70HVi1xEMfTbfuJugjB1s3NypUJ044Mr0VKh7AwHEA4bdWoekE3Kn/11mJbaTpGyxNzKIPc8Us
IVkhDzyccnUNOdRoVOzLViMjtHJdNVdHnRv2ghJiMUtD/aLAuIDrVu2xdr2y3a6r0T4WMEHS8ZKl
kZQQ1+sg9F5uZ5Jy7/0gXMSw48FUvjta38jUXeaTGTd3lCUDJNK0lkEUcu3jqi+H8x7DuL+IEaQS
en/HxAnRMNDzDEaCD29b5ciQANdIqMThJu+7ejlOhuPEL5EufA43rrpsOlM0GaxGcAV4NsWYA4o3
x7RYOovh27G2PgbL4Nsyq2KXVuu8firNjvKWqIiPIEC627ctY6nVJGw9v9JpBpI/bEoUMgg6v7zy
+em+2X7v3AjI8MPD061pNb6ZDoq4xAzAxAZX5nVAWcDFQF2jenJzFCBhRmLX60rjG6PgOveq2xal
mz6Zryh6/IJZWFmm6ZPH+5eNjZ6WkyVLTg3bcZ5GwDdKpogdwsH6iPiyyIKTseoEJPsSVXZpjcAg
7lOakz8KhHDuSS5EjWZNBJblbyimQy194Ri2Yi6Rc7Kgzqu4R8BggPnfE3ylfHQMGGqlYcMvdQCN
ngkW9pIjBodE0+UVBR3kNf0YrcglBb5DVMNdrLZI7Bf96eyPLzkOFBCjTwzelwYRfGTvYM/YpRqe
OUhoo+1Vo2Z7wJ+ZUDzLIar1I9PDoL0Zpx6tj9RO2jb/FD6WXbecv4x6m8eBhacgB+CSa6AN0MSb
ZLpZ1UOSWXd5RK80j4aHvvXol0ffnW/3VYKAi6tLgqyMiOL13Bewn4bnCnZuKStlUAeqAUm7NWuF
iFIxjiM97TmwbE7opqQr9Nvx/3E4zQk3rgISJpVo513mCZCJgmdCSwxDBYn7klJnu3iP7TgLY63t
BmgdwdmS61AS7ZZtQklKJeaTcRI1UMOQBiCrT/OkeUzF1vyHG+jyxC423j7mj/4mvj3zkUu0SQL4
MzGa1tV1jmNPHgwRd5r14FuAjhvBHfdvv65f54L1mtE1BY3j4blX9go27Lw4J5vR/KP7ndC45qwo
bxHJzFRti5UUKl/Rbfbj2REDph5oQm6qqhYRHOOxUTEC5fl960B0luov91CmcaqbAa/0iHDCI4CA
2gEXTR6UYvMufEZ4pEitYnC/Z2LRd+/0u1NJ9vrbWW8eLGMCd64Sh7vyIRfgd3UFGoAzv4i43Va3
G0afZP30rrJjb2SnknhRh9TSX1d8wcIf9kMOYRWlQrFMgtGxFRUsotYPtvEGLGHPX76CqtaPojIO
OjkpRv2W8pd47sNza3KRmYWiWeeCPy9J/AVkac1ZCihXUA5l5DLoEATxTKBzfYLoxjfdmFM7wXpj
vvg1oIDMeZuk8EheHaMs6ahzcWu6UIhdMWYtPY+v1TmUNwobtH8KLy5w4JQdGNqMPFsRYw+gpEAB
7bJAblCLcC0wi/mDZX5v48nSOZEai2YVB/yfDUPgIcIsyiRTzfuu9lTSJ4J63C8XG6endTGwr2T4
bQ8zTTxZn2tbsCmYp+xB/pge4qLUVEhVRlnoXWDBaQFO95zyNzG4Wa/ZGNiGE8rM9hVPWsg4Azhr
uOFn8k/R61fUMPB7Tu3vqD9PtNXE+9LUyWgS9ZOoMtyJ7IMkK9aG8XM7dscBHOJ/IalHGC4cwMom
jrrSp2gdTgdmw/1T7fNnvUojuoglk4RO2OEkBH6Q+TYSXw4mz3fhFDrJeL/ZrBURGCbsoqrxNE/i
orP6jxBms4gcpLm5m97tMlH7s0NTNvUXtUM6iTfvUm/aGHQSCS3uOV7AvOAjLABZeHBPOfsOqAoD
h4RlPmoO2iF5+7CwRiYL3JdS3flAxtVLiV7GQjni3pKB4IHt//90BT3RDyYMvNo4xEBjHw4uKHMD
X4OFUxgRHlNJF1Tkg5qkfMWkjeakE8WDInMcVx86xKwx+9uQl8bhQYngMlLI+aaASVAjig/mH4gl
8t6pS4+sEhzoPubmU5eqiVVUWwSaUQT7ZkjkcIr51bzvV7cPXtxOrpypLCrkq2xFBF8CJWudcVeM
qq240U50Nz5KZZ/ei1Qw1IytsSz4nWINVYI0X6L3MNslTeRjjSaJYOjP9IN509KOEcpDbzc6KCzU
5J10DjOZxTU+1zP9QNoStdOhiiykFDsKOGiyIMSFrbgrFzQkhDtJTxWc/6Evi+RtVs9T4tHvy08i
4wyo3UcnRYJ0veaoD0zDkDUDYNM4jelQUJewIgMhpgTJX58um/CCjlkY0b4dRPt18rz3LQkzwrg8
H4eM+/LTh8GHn9WQ3oDqo+cT6nMlu3MKLzrmrrQAGtaPu5xteKMABfGTFllZKpL2MBpiVNk6CBgT
+lb74X6H6ZvByTFrNDrulzvu0v+7Z1iQgCAdfmjv7rrmK1BoFCxzq7v6OjWBhIiTvIbn9vr2to7d
9Yf2KLIM5X198KZ4WO74iRJBekZvSkGKQYZI/tyxq0y7iHt+Q/yFdRARecUhl9JuQBFb7oMXXMGS
0MxlLjnplhYPi8ukM39rBJM+icKduzyYiYUe3lOKzKbKRnQ0IeJnWZE43vqE2pTswMM4mpKPmCZf
uUjxz8OhkKdYvv2xsFmloloG6ssRuvq/FwvVeWDWtmuAgt9rmFAm4pjaVGccuLn2uMoYzsOUzIyz
p7gf8sX3SaDaqKke8jbj8wypQrjx6FmsnXAvbc1DRTGHlRYpknGJOZN5QJdpLwU0SW9g7xBJZ5p4
poGZ1/dhDz7IdzitRxllvbB11IFSfM4isus6DTlwp3Q20r03YLndEvAj7GLH37m47l2imKt1wGLG
/8wyI1twqthhC8aTKERtLXEKYgj/ul1UhHHg7NOnfcDKKNu+HB7kSs5VaCqlK+BDz6WshQmXDQI4
RqNuxzXO7SyYP3gc+40HlF+JWL9khGT4V6cc7l2Mxv4DjFG+a6xM3KiLsnZ42qMd/+WgywPiJn7Y
FskE7dgib0yw6eI1+CAXLKI38TVqB9YMbQTeQyRk/l1I2TmKsNr4pboUQv0H4Mjwd8EKbmwbAaCt
SOcc/7Wt32YkX4JIgjXK/PUp9CXGO+M7RWNTDQ7t72eDhXL8aCeuaOd0b+1FcUmbEl1bL6jq6UNo
Kdy4XEK37aIR9bFDeunlrYLX3upHLVE35TL+gSNznyE7NZ2YKZGjKEqL8gTRK7CI8VtHkOaZkfwg
5V7iDiwYWCV5/OwNM65XCQ7roL9iH+DtKlPvHIjTxI6yBS19mR0qmkq030YJkcCof8xkVtv5f6rx
0vtJ0t7und+FzMKWPtrsAOjHzcgLyUXnHZyosgZ6BqS5QrFztBK1L5ivBh0/HjfjnVOm4iQ4KLWm
2MpW8OLQgvNyPZzg+UnNDbVh4QmGJT6mqNyGrTlE9F6p6k69rOienZjucrOpwQBU9tU/I/Qs35+O
QevbWpTbKTipC0YZRGT6hmRAI7FhveWWCgKxMxanvKZmPIVioPI7mgFAtkOpPmpmIKUVe92Aj7x/
ZiCEijEEGywbe674Uc6PKvarVEjn7EjXMR5c6PH57GyqTkuA3tF8v0V1fsRMDZZc9s3nuctFCAhd
wHzce6ad+06T5+EIOqzHbRmLv2WvFLuTTnaNce12cOHVKzhm/Y+/xRWWZjKOCmXEefX/FaZu0DCu
yDVvvp9gOm5cWFaTr24F8WqgPGS/BeEpr0U1ZfqaE9966ZfVWv2EvVa3ak9ovDIB3XpBvwpkVjta
zxgsWUIQOH5/tDJOqF8V3p4QJsnrfLSv2XU57WNSGCMOcXjKTos4S2YSjk0an57Rb5zq8uFgzbXJ
tVy7sfglX+amgvseYwqKEY9eOtUpOblZ9aleXdzKaPdKW8Y9aVsKRnAa06gzHhOzvcAwOr5BTLdR
iJHiuk7PO30kQnkUl9ySO6ZnUaU6Fi5vEjZKwNJQDdA/VfGGdmXN4cFKMhE+Ia0U7vFnQ5+WGkJ/
c1AcLp/yUbs+uPyaeO/wAiFG8W1SkUujddpYFUlVC6MQx9XABTDWkqgcKQQbFzP+zh1v6UZP8udY
HvEYWltKnSWuuYTo/ETlFvgRLJaj7XSBbYCR/DWqfXt8tvrf5KCKGSS4z5kHyPCuQEajpfxYJMRz
K7NruQWMofvqtMoqtjhjDbbCQKTVucHqg4OsVR6Xhr01iJEO4k3DUSwpzRv9ZW1irSkXJReSAkIr
yl7NL65QEoQCznuiY/ENTj0M5n9ZnHFvG1rkD6A66YHCe/mmKW4fcEbKsqkGz6Hfympmeap9fQtH
WtlaYpI5YOicqwyvMTYH0Jf6hibjmaZR68+Mr+C4geuE4faOexjN8TmgapD3o2vxhbQGG64QSvk7
jOFdkjdyPJBHvcu46dbg29HGn7zWkwRUyR9y8VmDovw20wnsiurcuQC5YsFFwDLCSjOOAwnPOVNJ
pmqHAuIkO0nISkeAViCRVLrcwcQDYoRfYG6dzKZoW2iyiPijBOMsdpN6c9MlsdEFZkCoPxR0pi1Z
n2LcNFjySK/zY8dCmz69Da+D2qK9xeCRG27o+TrHvbhU+XGVhLwbAah7HGrEnDzSxkGW37riyFLk
HgBspVsv6d9whxVVUU2T4ZHDjResDtIPTeAuMYwedPXf12EkStZP9jHP78GccntUosJtXoFAsc+4
DdmE85pGo7+CeFHoAm24c17n3jjDrFI+u4EFsiOA3nn9aI09RzFMvZXS59TkD19/QW96sUOjH5Mn
boWJb7Sc5nzNyFMH9qwHy/dgDCNtlxoZ8Q65YuldIocrWzSqqhtKnLZ3ovtrTtdqvgwzaO7f+1lS
u91i4L4B8wHZpXq5F58hcX+B1UsCilPrhvzS4Ei6MRRE30PvZtH/JErCjyjJt/QO9SG49vfRY6yJ
5Z9BMyx+KAYV8rWuKO6z2rpHLWjGMro0NDXmTKGldAbyizER72LRm/S51LskoRa2bOdPeNOAIBRS
OyG/p+xhNI9mussO4mfKzWB9ZaLGD97ckp+E9fbvWlZtM3hCfuZxozvUOcUGCyFRABbh0nqFJtxR
P/mb6vweapaZgYFbmbX8Mxt/0DvX32L+Yamhkn4mLKHRPulB3qKvXXOoLit80asmYnMfYW4vnNwp
wnR9kmoLvoy3hfHfh/Z2Mi/ADBBc4NgyomeUPou3zdbeNGDTEflFu8Lqk7YvpkpO4VaBnQnTeLUE
MRj+jMZdqpb3pVddMTC2ZP1qHtyBXEeZIUHaEg+CfzV/aNxwSqgMZASNi8tsnXyUa0cMMoWnkaW1
GkAjKCMoxCeQ9Sdxke1bMKZExbCUrrwdCh6w51DiQEHszV0laWdLumKBtMSBs4ze8lN590Z2//73
sSX4wHbE/uxAmWkeBJtHrqJ1Wnh3kxyrT9O16KVhY5KpqSLSMYT6hrDC3rzwOvoLffXG3UV2VRTX
/2H8M4JqLMuK/Eplg1YddeAjSO24BA/JXWzkNVVf2pCW1id8weDWl+5FzPhREmpY9ypABofXevuy
+OQtiUr3sTE+EABFvd4/sR7GpAA/vZ4fvsEWum+MHatPKUTTfl/yKOyHROcjZ6KhfhZjzG25y/xT
E13353VeQB+Zz3sfGEoGAHTrIeoe0t4tpEI0i/FjJkv9SVTlBps9eUpYPFwLNb/Uhf3JxAsdiyAi
RoqWT9bVgbFuaL03z9vmoJdYqU4QEOJr2odI8v3imkA4qYEbo7RIi/4wbzu9+Ngfg4Ky3XXypHV7
TyeqI1ummrldCQhS4FfzF2LA0lVXhDQXtjms61qgjXj0np41jtn9TPvtIVghjvmCU5xHpXAwcAbM
LKpWFq6xP8z7/R2yD3mg3s7zcMYq9StZyoUgymhD7+W3jPXf+tX8rhfOe6xdh597fhbJBOPc6F6D
3dunqV2wiHUhfTR14Rp8np8c3BYTtuXF/FHqVTA6zLh59ohT/tLWmht3wcwX/zMHIWDBDDeE+niO
EPKosHydRk9xoB2u8iAe4I5exhqcNXOXTRkx8uFDleEwgzCvoKHkXlvMvqPTWri5uN/1lMom5hSC
/9bsxCkiY11W621JvXipBQQ4LdwJ16JYsy4wqNuDT0B0+QqdggaCI1L4sBxzuXvrR7MiPTQYhKsj
LBwEGS8AdUZj/keT7DyOysiIO7oM0jeTTYVxz0OhNyp05jiRgbwlELXvP6Xtq0r0NIZsRzJfvtS4
96qe12p1Rx4NCuWSx0LIyYFbqIhYDmPRBhRlXz+qBF9DtFGQK9V8cwCtdiJoMsthfZhFgOwefMbc
RDsYb8gL7b9312Or9aT8uzSpmpcnVcWgaO0VBJOJXr0uqfFL2DGD2WIbiAosu9ms+dup3QHGiKy/
dtbe31fludclVPkQgVQxmNHTe2nC+r+DP12BaGnaaCBqK5v4LTw5JSSiZRedbMagjU0qP3ZDhMTF
WyLFyRmiiCbwykpaHxDUD0WMDdJPMymQ5BUZSbLLM6CQjHAbn0rKeXQUemEAqViky9Zp0FKsGV+h
FbE5gSL3qGXmWUM6q1oLufGhxOz56oA2ibmFhaYsSwSsjIzDglqnvpXR0fxRUK+yZyCl35WI0RcT
GTFo7bbVBllk+DNgLk1owP8qtyfnLBrtuK4aFjCHB+ITKehhpTBLeIyZF8GMxB/KSr86NSdB0sw1
vTvPg+12pSD8+iZY6/pftjbrsEI1FJ/dK+86k70rmbBSGiCvYhjIQvbxcwStEeDRMoGkroJ1DD+7
jquY8uOesI7KzP6LwUECQKL/KJuoc78l6/y7ke7eKyb9U3ZdEBrTICgq1sOeK2ONlZkH0mSOnnTd
tt1r9XO9D5iktjq5i81uT0evZ48fS6nK+cIW7h4BPqe8LfvGbs0oumlD8D8RCHtuGI98NBsQB9md
UDOD1L+jXU5L84Sh2P2UC21mVLTxaNv6sgGiHwEurcfTHUAv0JzwscH5WUZTpUOj23Cz2eJeV1+p
ClENSbY5bnFI9zJoelE0cWjqECsJUQwpaZ7al4quDjxfc9RzwyDafdov4ST/AiYPM596SPjUuSCF
UdZlg2a1euR/nzBQIJo1aEB221xZ74/gwHYP8a7dxfkHJ/aw6RJdb5yJIAvfZjQpQFTnEvnATbow
BpArxuhT5oN8w9DQIP2Hmyn3GOEFXNXzytcbPi2O8NTLfhXrTyAw7gynSRckcTmZ29IESrjNGgaS
SbQ22PQGQROA7FbZwPL0dDSdiEbAv9mdWPH7AqVNL2SXFaoD8gMIbM19JS+yrFxY8odOrLNv/Mg0
a9HV8wHHwaMvlX2VUY+uUzDVjMuFYIe1nRbF0w0h3atlzZtO2bYc36phZqs59k0SjAqbNcJLNukB
Reavv9BT7VvzSrH/6qRERpeHmjJxpKVhCB4iHgWLM2PWD6h+IV71bDZnY1btNHqyz7T4TjWvuRWS
ksT2YUSE1aA3ZocYleQJljP8DnWLF6XkGArVjD70VRmKAyvKU+tAYoY4oNZXw5ChtwZve594tgUQ
nOvv76hQCwfmTKOdFCuning/VMGutz28TvoeIssU6/dkvMhNDe2qmKuBZJm87vY6G2PvVVtdBcKm
7N4X0VbelAvE66zWP8FPGP+KvxP6rdyaj7vYWKoUpkCwJ6GtddcYQYNO8UxYNmf3yEEROMA7xtU5
vSMqV3ouCOkraF7WsBkyLrMs+R+++zQTe3cC8p9AKVgQKlqXKQYO0sGcQG6ghHCjdgIf5OYLO9u2
VSh2cbpRd+VGFpDyXZAy/gx3SqlqWpu/+hxWl4FfNwxwL5N3O4kjiOKM5ufC4hV0ZsN1G+3M7wmx
AMQiWV8lc0uMGP9NN9fqQfkKMj/wZMbqsN0JryuASHsk6abq0/n54uMwgJ+HfefWwt2ce30co5dP
NS+4W0GU7Cv0Y31W0lMsyzMF2wH3z2jGAMLjo6SNPiukw8p8peQMNLBKKRc85Kvv8/w0SFAGMEhs
S1N6phrFfQp/E87cELLYW7f3zTTx/woDqf5e3gsabsPqBN40LqaRDTAqElyYhRhVt98S9Vp0lZwu
+G9zQMdckSl2uznT5cnHckKap8yB8UgF5tH2MFbHwRZGLsaMg1G6m2rL6aY5Kk41xx1EAPIHsON1
Q0EKI2n9oLhvNBjzHhz7LAP+vHKrVD+12epB4q49ytVSBffJPeUsnXvTHtbL0FK3KURzp46jTXTi
EjpzTucsbG39wztJoSohs3oZG9a69uH5Z9i2S7BHev8H0J+0mgC1ovZKO01+A21vDCJKZitJqj+s
+gO/ctSFQbTZzitahjLAK6YFfW7zIpqaQbEeFr/2ELAhYJDLN/B+RjHh4kiO918lIjirCjAcizPX
E7PcQWF/84+5HYVmQPvVYPN+Djo04XaYvV/XKlQcwwewaam0ileFJxJpoA/O+sN+3ruyVi3sTpFM
Rws8XT39iZAezhf7ejAVaSo9C9XsxFcmAqPAl/iN3kq/KMou0RIulH2A3OL0Jsy8zkYVx1vzA4i5
cr+XuZm7JQslOyop2pG5mSF80nKjmlAUtvKX52kJO4woxhoamuQAnUDqPZTEkET/NOFQwgbUWKcg
d/+s1kTw0t6mA4lIjuedKuBOm3zBuLS8VwdN51FDaOnbFmw/ERV6UjpEQWAfDwJ3Fd1JgZzhHE93
RPs7lRdBKed05DaHuYbydvDMM334atauWWFxLupULKctCwRNPeMr8PjbfVKLn1cLjB302BvX375u
FGbS9ciQtSAXWdtGArCc53f1IdjDV3gjBIpkmObRBsJwfHrBlzHFJWYp9+d/ZAOm0O8M6H3JNa9d
lQNG3SaiLJGuB9ZQ5hBSxhj4SLBDBwKug2WaskqsS3+ScMVfAgXvE+5MSQIEc5+xkCf4i9kB6J2s
JsTZuzRFsYdi4FDbOuABcRihgFagdmi2loVrMdGHrzMpBBCfmSUikmirJlnJTyCxsT2BhoJxCxux
y+GljwN9+ryEpjW5fnuOcHgrSIf3BmUDJiTXrj3tCGti+FnTG7hEyHhkdk43AuZDiUnUORKFrws6
JDwcot27oTjrLo3Sva+V/TvKLAJAUPfAMswwR/sigRBN9xomt+adNAoNKT8ImEva+IEItXKMbEqk
iXURaLOgr5MCDd1XfhTssxJ+0PjWuCTJdMzRR5KS6xF8aZlBJ+47GuPZcXYY+Ap7SBiRnIAPkbLx
sJCb9xz0BJNbeWXszK6jUSytLkPZ6rMibD1NGxdo3OGNuUEhclK2WixgeIT+uwOaYvMKJw65GpTd
k1Jdt6CknyvoijR1SzgbB5Jnz/upscyAcX3QwBGuKnQWGpXQ4H55evas8+qKRhM4nsAn+5+uDcm6
6LzYGoDpcT1xMM4/M2ZXY7fD6nx+6XIrDUfFdJSDEu4B4VJPK0SocFq0qA+c+8GNmN3DGu7XwDcc
xflpJihupr7bUlk67Clz+s2BCafsDu3zk4FB29cU1KDL8aMgSOuUYaRWYkQHs5vBhl8IoQoZLNPw
wXPpxLddOOHhwnYo2gEfWH4rLs60m22mvWeGhj8JX7+AnsrRCsM6HjA3A7ohJh3JLtzNsUa//T68
uxRReQ2ZGMkyJ4E6coXOtcmA2Yxv701LGugk1MqEiwEUX1EpI/64jgLnXMQ0w6OtT1gpCFjINVaY
qmGKw1xFr/MqpsqvYJuTNIqEGYttGLUNU3TrHv8DOPfBrUAQ1C240Q2QlGmaJNZvRcpJRilJWnNs
WHR3Z2nSMP6cBLkXGJpkvBB7RlZGHOGA1BPRim2MsvFseQ9bnaiCMtDlBm48+2X5OSZR/u8xB1tt
rHhp5kperKN/9sTK9r7VlelPGAECqN/noSIPxVk4PH/Dy7hF/l5CCuwDLT64VIdmjjm7vhPHHZen
XcEbT/JVkl3GML+x1BGg9bjjVUM44CS1xWaECeCHAiwddaNp5RuSNBiVKgy1QOtBzOXB20Am2MIV
bJy/R5vQEvFEHvjT8vd814QM+VDEIFP4JBCtdG9d52jQ466oek49x3u6X9hfj12YUe3+TUvMX76d
pJLDA90Y2dQXfLPDQFoiQmVA1WjzrNKCSTWMxTZXTesR6M8bS6nHKy1bNKerAINdN4seNk4Z2N7C
5zh7/rL2CcUDvviUL+XxX2J8fvxIATLN5oQYAYXwfqacr+4tgV7Y+8VymXdfIvlOnt90Xbq9LHpS
LQcZ6gGpAvT/GZ1+c9JC1TmHTDW09xWdVnvwpJhTmba5xRa8uZ7HgcyoESqs/TzM1dCVT+wCznMV
jULfjaQBZQzoa6X1BGByXmkFh7OkWFL6O6/2mjbglr7DXdrWFjId5wn5LFpsxfz+YIO5c3frpjDJ
0ekSCxDucvKpFsY/VwyfJRBKrPmgIi3oq+3PzA3bTn+b2IOaRwRT+YTylaD3bg9Y49Y4MnMBBVtA
b0j5+49gk2b5hhJJlE62ZD5sT+yDpq4fug81NTz2wvx0nii8OtY3CBFmz1Pm3+cHR6+zK8xHveZI
DcZ2Af8a1yISHIiOjre+lCoHXv2G7gpxXWXT97WzF8Wk/vrKbO4rgO202kQQjgREf+9LTZ67xQgz
jWU4Mp9BmwtGI/B7OopFKq89Fulo4V35U68paJGiC7+0iPVWNmcQ1prhJ1zajb8x7iXO2EbYCq1u
M7eUpS8Sm1VIPfTpmtWYXLTIy6ll/itlWmF65PEGFycckqW6zGkLsvYmh3jdUTWZAHMFg4ZK/+VO
NeJDz0yXKRwcF/smozzeBY3OBX/qSjrew7qeBug5fuHJeWz7hugtE12mf3ErPGh39DzQ1MEZeYnQ
bxnRsrEPOhhsFqvhqKL2rA5Ip9R/DWAHh71XG8K6AK8YzX5B8/5lgK8kW1y+vjTCRLEv/aNMXe8f
RgEMhDMdqaikcgQp5TG2WwfvFRjxNU96gy+L+92cNuqRK58ZzbNuhgfR4e00mzGtV4ZOhIj474JC
LO+uR6fibWx0/WrCnixdeBuqXaJlkFU4DbiroqZRmdW5IHP1LGtUzqB7U9mvuCGnaP5qKVIPCBLA
56Kg6Zo3/4AO+evUx/Oy04j+meryVlEAiiR4R9Rv57TanwfowEEbhDANZXKqVgoEJIwIWCDsSDgg
Ke/RZ9iEUan+ZgNP2Z2KF/1vfIZDKFrIn8Fmn7Nu/ktojs5kJG3jSsFrAgo9l3KgfZRVcJAOfZ7p
q6tBxumAnhjzJ0Nes0JbvrEo58vYsuzloNbqaODTTDgOO5vANve3golo9OTpPwhLLL2ZZ3fdIoe0
rjklsGoS1CLEZrMor1+qJNdtLAd6ijT7pkwKTy/S5NtuDVb92CDlKk7vFU2y9MjchvnGDqPMeAZ4
UMGE0QgQbSBlIU6vMk6y8+8hUcBIESC6pcfIM6gA1wKFTtcY/JFgMjRPwI9y4lgqMwQ4G2nsflXx
/0xx1Pr3TLH/BwYgYjngFPNjDqsLyvOlOVF0wUQNLPkdWpZ12gdc1ukI+tTRe3o9AYEqJ6Dy14Pb
ohWNDP2l1jaSGEKYvq0ZvlCprprfx3Sob0GWmPW590Hpjueh8XskHc69l1VGpKnbj+tHI+V47wzo
ttxWR+rLg+Pe7a4ovXr56a52sDhg8xC1MOmQpYw0T8IlNQZ4PmZEakJxUZQiZjI5d4qGL31/5hhU
r7RgMIcsvBhjlznvV+W3tDsZO0/lYHMFrXCabd5QtUi7TNIQ+jv3L5Xr5IZcAjCx/ezYNhIgEhyl
JgLB1tGOQ7vzjpt8izARFyI5Mj9TzdnvQHFLC1107TPNqgL/SBubFB9+2pRaxsvbsoOpF1IhDPYe
l7yCFIWwWQ54XQhbz9fctMw6NV97FCtLvCjUU5eCL6AD2OW9xqLBqzUhwY61Rtb2HvgVAyL+Gi+D
djbpaf9z1PIkPRzZNvPxmwK9XRss/igYHmHIrXj+Axwb2Pm9Ud5yUZSJ3BMd8L9oIT0+S8JkI4Vf
VV2AbhFGrNK2M/YrHvcAdtjHHXp9HX5vaHzr3cwdW0+8Ef5hTKYN/t19gS4H37M7I9mqQfKsRzsW
Lp+/qcoLE23M1ZdAa0XdDb7vBLIPMvsuaYEdTNk+XQ/5kLmvg3GNLMGe6YjU/lJF4MyK4dMFmQsY
520E8mygMblE0TQrMN+Mi8gb84zIh52M5ZOL+9TcOUAWScmj18poRQid42/qMCZwA61LUnhwOUci
84TJbLFMmMcCa0fG2q+bXzmRkyNXAy/xqkGegDNjCZkOgP699k1kzwsC5XgiQcOJrP8eJx9NQ14N
8SUwY1PAghkLuA2BDJJYL6Z9pcW9Fq5jq5VvjCfvSubjc0FiRhDrgRvQinc6es3KGIpei7nbP3qm
DuH2+Sa7EfgBpiHQlG/99UDMNnUP4D/UTrrY0aq16YPzcyF5AL6GMIaliy7i+323TcNsy6R3Cchm
NqnovqE/l1ZAXnDJT969ov/Jl22Bip+vXlqK/Xbb6CcPJMOAERIQuEyI8ax256j6q48Z2HX4Z12A
7M0ghDIgScFb68Ex2MUX/QpFIpFvJU+SQvSBFK0VIjhzxKE+ZBcJA8SNJ2DVjvoXIkDlUu8dn1io
85vZ1+DSKLZUO1jmVUocUmeHdl+yd65lTsCQILVcBWM28KRrXcAMSlO/gd4wnEYucx1DVPbk1nsY
+/T1gUCIMzMbwmHWm7i2gMtAKaSm6mk6jBaK85b5nysGNHJa6jnGti2vKf1y/wxmhtFNA2BPwYN5
CCirKMUAqfQKEjDxO/HcQ/asgd9KNf07GWi3hc0WWlBRUzepIu5POMlrpj+UwKqrI5LncfbO7zvu
NcLjyPKtD7t0v+2AHgiABDfGfOW+t7Lp0ITquCo2lJSWec7+Wucv1llt6Ulxuyj9k3nDu5lARUZx
dqXeJAxslIJhteY20thxW7NEJZexVAcEM/Yp3PMaAGFx70Hx7mLfhOwsVFf4vkQ4GTori3BGAtGH
/LfgwF7t+EzNu2IzN5cGY8W8xnWpXiaQ63Sd4nZ/5IWxVexIBV5Lb3780ZM6NIwer53FJKleNDz+
+7Da3U17MOlA8UKepG/lxtZ5Z3IcZJtsFsgaTf93TR9SXv+b+bQA7CKwzYACzeM68qYvE3f5nVkd
RskF5kgBfWs5hoTTgqI8oPsHRROhErS05fzXpnh+UfiMtRXA0dmzAltIJVCsctrzNNofYDbbVeuY
KfdlTQ0hWoT7GgQiu0UY8CBw4A9AIAQmCZ/QyOKrujQWke4h8kWDvnWtnlLGH/7ni5jbZReBL5/S
PJ8Nh4zF7h1r3BAkSmNlMc5O2cEW1G1oGDktWVUJou8fEMxdxMgG1eg6+WRf773pNnQ19xSkDgEV
V+stIcY54jW2jDF3SCs66RErXflrs4ai1yILqIemgNZDblRdoQXPBspWP+lLwausQIcqjBjIGChZ
dKBQ5LKHfoc4V+mkPsCz1VDuHRm7ITrP81dXBlG9nDA8ahav2zr1h1WjSFYFsbauq0wLWFXVPOeG
29kV8pYVWKpIExqF6ZEN5xKnCBqvkmt27h9ZlEM1sWuejzPDufb2/FzLpjm0hZm7+EuDa/vhq09A
c0IQ6VX3TFQJ/NpR23GgFJbwzQK+wOtcJGb7rDcUAvB380lLcVOiD97wYJdsh6OsAHQzuxtGN14y
gSoR4ke3K8cxuwmbnnP108h+KHVYrlrKBQHTJG0SYRINQRVsVdVPXcVt+ANGXHYu1pQoD3PcBnBO
cYDMtemm9V30XZtY4Nk/4EvfWjUrTee5kbsXvzFOtCeyU+Bj1zms/kcwio98E7J6t6gXoZvAuehB
FXtWzVui7k7f8elKkuRu1FflN65VKOusR5KtBX7uCGrJwDmo0dtyr75cr819s7sM98p1kyjqDdvP
UV+J2BW0ivkXh4D01wUExz4NyRTh06pS3s3u4koNiE/sbuAyIgX1/jW8EbmlQQAIQSCjBWcSJAUJ
cO9IbRJmrMPDdXM1F3EK0Ld1qcIX4XiHAGlIONFmMNDe7JVbstkP5f2kzWJ8JbHSihlwuFf3kEuu
EFJLNoxKu9IlP2lG9mP5ho6r/c/S8MwIkzdxt4SNhzkBXAGtyRl/C2PBROioueLv2IZ7ud/rKqpe
Y9gjwLurFjR9loYcyYo3cdCWhgxi+Sh1l3v0SEo0GU3AJrTHuX22dTVotb6pe7vtXgW/dbS2M6Fy
ivUVo+LKEu1RNXuTb3uwLxHuPyn/XFnMypxQOBq+bYzl+EipPp2Ir1NPfftS13n8Sy4hy9QQWvxR
6GNW1cd6Ace4OFuhEy8Oe9FvYbZ37gh5O6T33bs9eu/ULRRBoNPi54aJ8vcod+jhsiSGgQ2NwQrK
OnKFE/Zb8tWRp4MDFvGjeBJrp+22Tf/kPVm+7BYO1n08RF31atjiyObEXRiP3o+v904F5KaJAms2
WJ8TXjnImzRTTqRFzV1ev2Q1cqv/XFqauPXzPDdwgXgWZpLlkrENjATqIMZTntzo1GAIQQ5vYfOf
zNmsUA+lXt+fZOjgF9YlO5e9Jld/0K5BCH0LYh6XIOasQqhdquWy2oUdeGrcijtg99Qc2zvLUhzM
1U8X3bTzhB9ExEluDT0h4gfO5NpMwRUIQyTLdGaVZoQ2+VatjvmntssC/lXaCk8i8cVFUnh0Fgwl
kruPD/x8bhRiMfDY5CnCcsYOxG8dogl8eLiba73QXHFQm1sWPKpn8+mqRf4dDSSCANas0l+UJgF/
H3dj0P4D9ZaRlNz0rorqxf1OuEfAQ8w8bdFep17bgG4hUfJKPsbqWzmX1SiUXAknXwoi1OYslS9P
nQXRsjSSML1IZV2e5aqVpkfVuS7B4ZZJK/C50GYDEOkZHpQ6ABc6clY3a0nr8PzJqVlqwOj8dmT6
QOX6tgvayallLlVmFcCjlOhcVWa4aHeuBvezJRW8tvPiRk3CouOFE6oH4fw0twNJROhPZtQlo4LL
XHk4vmoXdnQ5LIPFCjbQGVzYqExKieu6Hlz7D1pO+n+nWgTk5Aaqh8A4nNd9b1cuutUWrjVKT5jD
V5HWeKM7qyuEv7ugd0Shr5WwSvRI1EBfGRG8pkylZaGybeSQ5N2KkW739JubHrIy2I4cF6bic7oE
n33zpJarcpZnHyLFfCuUOrgdB1I1ft7kSpnzGAxqJ8MZ9IufABsROvOpezQUw+48aEWyWLVbki4b
aaN95xK87U7k9BLrVsMMTKLmbgMALwO0xw2pai4pEB+Ixs28PBGEYAchz8qcqMT1RsaXP18OmMu1
Zfn702uiVFEJWNDbzlUVUnJnYIPa3t7V+lccwZv/Eje6164H9YdUat1u7WezR/jU2VOpV9GxsaBJ
MawfWOlyFeEFM9E9OHPtG2EansR7at/1vLkh4GG+cqkC8a4wTLp07/aUC9wdvj8BdumMl2LBEJ50
nYpgjWW7LR2/vfZL9/bbxM9Mi0JfP8EuqbIu2jaoMgTrr5ezsiP+uNJhS7jbWJJPGpdNpwkAVFlZ
gr9wD1UEwHu3hrjuUBNSmSDmuPTbOPgZ7F+P9CTcGzvbrAXchj73YsITmHQK3YbZzJJ4wSE/ySDI
kFKtXhEmZaMorHYdsUkM6zY3uhXQPgaMyn1UadNxsyUIpLKnNZyDgz1Cs5y9AglgxV9CCBjqMuED
mpQ5LS0G3ql0KhfL2RvlvKqSeiBYz2gquMDHfoiYiFjgEfPIHy1ZO1k5/NE4jXo9vtFCWddIJuFO
74wYHKeG0JUWWnYJXS8TuEBmS/U0se1S4gW6T7uHJOTAWf7cEIEZAw7jSkMRHjDhl7H0GH8yTSl6
ATwc5/hn9wa3giAZpns1W8G3zNHUVHqxfw+e393xedHghZD8NII6P2gxgyvARQcFuP+k2kIJd5ki
VqqnpJ7JB9sDLsJb+ezl8OMvMS/vQumPUST+2z+cMzimxShN9b5/X+4GP13vdEObVoMJ8wxu7+hx
8XfHvtgFUky/5t/HOtZw5hizmEkGAOrhkIJWYY4t4HkxCd6Z7XVskrSBXE9IIPZc3SxDI5BbILKP
CwnegQOGWYbdsxsayKGwbKuKiU9BRt06XoDYRutO4ozJuGgR5jENLKumohcIg9cKFBMjFaOsw3To
ER+EJ/owCKAvWq78gFBN3gznKf0WTRuiYrzZBnvXpW9MEVBVwOsI6W7JYo8ExCTmh3/IIU2jn5kf
jo1hYFPLh79uz0t+7db0J9tUD9tsSJz4Is7dTZtaru5RwF+I4R/oP4lZ2R0HfLbwxdR/gXErRKcd
5xV7D6e/QX8zp8psMjT4aIwkId6WfTOySN4O6jf0SNvTlxg9yuRve7rPY9PacuXBQHQN4SMZPrBM
h6tgHLOPD5MtMbmcCOC4Y0P5wqY0Gl5ouwagjgkeiPfeWdytY92jXsHjuj/6Z23F+bbLpqnF+gnc
sSbPmUe7xcsaRtGb2B8ddCEj1bWs8ksvHmPbzZzJW7Mxgm8SA5ZGPFn/NMK0ywHC58SfAP5uvk6Z
z54o2gifxpmW4gDb6EEfkssvOmV8rFHKCQMc9PhedaWa+mAP0AeLSJymmnOKHkD+Jb6Xe4TOESG8
tAmEBpIJpjtpE188YdIzj9B0I9pdybqf2peLaoF4rVBBtoEO8N8UEly7u5zzfNvQIqmILx35tuAN
p5Pk2PkdUm4ZGlv+uFTYUzxUPNWZLPsdx6tyN7BQB9pT+t4SETp3lQre4Ce82IhyR3lBRYwSUwyR
S/4Og13JlxA4A5HEBQI8T30aOmQWyd19ObsdAzG4qSZvomHVcMcfu3GyUoX8wGtFFfe7s7uwTEzc
L2Qp0cugBPtytkjtyoXQ/Gpmbl6zQi6vZncaotonPPB/AShDDv/gR20W0plbkCDJyUEIL88zC9qt
uHuMOfUOCgdlCp4skbi3e+akL1cV3Vo9lB6IaQxoUsQspQerUJdsE/xmJ+kOh4q9/JQCHd56DD8R
aQL1o1Y5mjMe42v5L72YKSXOevDUCtzglI2at3RNhO86ENrRaDRWN7ZAhVu4Hbf5o15Uj6PI5Rcz
eB/LFAeozT5S4PE2rW3avOo/VppYvsCpc0wfhNvRVBFpn7bNc1pX+ySqCmOfssk8gVOV0GG1D4yO
afp7AuNyaW29y0+bt/gIlC72nuwLEiYePps7Q6ezIIPaIoye8Yiz5lxFiIpbU7OaOoJ+gF9oOzXm
1R2Mm9qoRjd3kQlIPw/q27LS7sy2WM/DKocxxvjEAcIbf6F21BZ9HjFSrdWZo1ItNJksyLk6e2aY
vsYnT7ZLQX5rONrQt5Iw1aKWBw5JT0MB3bzwA81kW804R9ei3Gna2L6C52kg54jT2wxloQ18B7Ij
UFfdrRY7uzTBETGkV1SWP7kcQVi5lEsNqGd3ptRrjIBpyuMi5MJRPt/tOCEAT4kqwOCLZiFS8Ous
E1b1wziH9grB41mCJ16NjqDp62+U2shwMmRPrTwQHVWRuhcSgGDhAiKlh/uycSceDR9cpgNkYOOn
jZAzOTT4U3LwCynoPVShyd+YbMtoeivCbtK5FPIzMgShxOGrZQvzSEkw9ILdi8104oa/vMntmQd1
9Lr9I4SV/Pgngxio6Rtqp1bjdUPkzPl0O6TIMFs6CtGxDfPUxIrgnlp+tYeP9NsRG3GPpZnu0NFS
qpvP62S2UGssaMqzKbuuLn8ABzR8VLALGDsTBdBltlBI5Czr6CchiNMj4n9NGU5/jbeV59NMzmHu
9TKybXvDhspK+fuuv5Lske7uCeT98Ff2Z4fpfhiutqekwnor5lfYiVCzkuTee1LypnthmSU4Fxxn
av+IcVU9fydw/DauzvY/5PE/sKMt1aeHFzhpNOphsrjhcUuqOSRqRqz1DjeTZv5mkXwQ0fxre1Jr
hiuxlPOEYzNFC7Sv/zvWk9aPwkhn0aDC0UwgzOh2TSwiEGLOQvk7JzTbqzW32IqLWBj87j5JyhP1
HtdfQMqFI35BBj4+U/FCJQxyj+NJej+t7lqAln4jpmNzQmoL4iKUmDn8+3A6bGESW20R0QU7ByNF
wp1Fuk9Co/paWEHaZkeWuQiSYFhgeXX93Ums8+2CIYURCvkOgiXpg5Uk0P4QS5m4dirym9ZtKdXZ
VJf1s/tUdz+0yU1Bo8aB5KdebDaZhA/6sY4ohi5OSf+YcTbBXRjPGaAG92up5fpHOzwyYvoWxVO5
Sj94BDV+axzaQjxNBF03a9b6JMWEc1lvRiY7ncANdh/m3v9vp4mijUGZ1r8trJgS4/7pIZWsSyfV
XLOWi+u+9WrUFMZ4b7OP/Rk7W5bpaK0sqsgDbinVghG85hzaEbsh6O6XXpDZgE3xCtl/grG0rAKN
yZOQS4g05q1O9JxwKX1WXenarGfws8BmH432ZKErtzYSJHoy1To4cGq6WwIKoB3XRh49JDyE4qLj
nKN06ifPHjTxxiwTFdRWY/OJMjV4UeXTvMBAh8Q2Yq5SEzqpkFKfsBtFdU9HHqJfd5UkI0KCnLmO
VHtELa7G0DOFpRMRLIdXEVpFPm4gGGjk/NYODGHXZskSaL0kxoc1fessq+2ugxFGxbm0ctc/R+23
AKPmKkhmFtCw2yiBY6HYaJoDvHuXMNpBAEoOKm9/tMW7Z9qYklCCHmCpEqSifRnJzLi85B+gjwfF
1gRhJGap8LxzHLvHVIBchGXU+DXsOCrRDVNcNwzgfW+JcUd4fgP6GMTKM6qjRNb7WjxAOF7JSgc5
c/bppvNtP2z7MXMXEq2nxkOTLR9ydSNGmXM82dxAMJMET4gkMrwWSiIPWCCaaIGmuvj8KTbjELhS
ew0jfzAf7l+eZNwgK/2We8EaUAhRkwa3nVc1qys0pvS9LAgZkANVYVxAxA4AA6qM2i0KjcWUGZLv
zJ8ub38W4Bl2TFYrF5uD1DSVDVEwfTYN1OJIF+iLurCSAsS/gAHRQHxC+VwWbeZZkAZ0wEDnf+vu
CBlIIEiU65oVVvqqcNQJ7LTP2+Qj70E7ooCnzYuosqvZyVvNnkDbbWL5zSJe3PIpS8ZHglWmyLqk
BZ+H6OEBww7Q1HnJ7qJ04oe/IDZA4NzFU2I3U3WLnM2WhprgTsICV9HdtwnRqy3pjMwOQRBY4SW7
7W+Q94Ws97axrjobPW574vefSpms1YSj/ID//TYOnT7XxOD5TMcyv10JQsl792qQPEhr/yrHUIpD
ZLB/TampSzun6HsHyEHPAuXYM1gURSp/mlGYvVhTEsYOTDIAY0aXxYiBnV3Qzp5yfXVEVPZTZFTb
HRDGjJWVruxK5OJY0WXA97P9OeYEHTp2iHZgnHyhYQ9nL42n9bghMkufx57xK2mN19BayKnfuynC
mbDIu6la+2USKqoxk0tr4mNjxGRyH56fsCs0znQ4Es+uQ2WbathuebLK10oe3kON9z+fLmqySpgU
07xuONgxGMzrZnMFYR6yO3VJXuEIgahjftqWAcnsAq1+v768krw5RPNWDeq0tQjxW0W+w6S/Nv/M
nMOJjgoz6NdVKLOhYb5R6E0hdvOLK7cVrcM+MVDhB48t4rL5I814ELM6Y1zB2y8Z7klkhG+EGkbt
IEIThMSINgx8lST4ePdGmy6a70/NPDwXcr8lN5jaGWZ/Z1Hri1Y9u+rMUaSOpaDr2TrBxfEXutAp
xjwzb5oXkYyQxQYU5Rix+/+crjtrwhUhryfiLfGYubegFjdAmwU5hzA1t1GkZ6Fi+xlKk3VUZ+yZ
oYIpkfdu0j0KwOmeEeYmk2HGlk5RNV3rQeVyfB0Tfqew2QnYPKm+BBjWDbPBIimCcjl6yb2ZUUsk
CTsl/zCrX4TYIA4fHxeokRw0ZtnPUL1BG2T9gSA9t19RrhPWa3c5BGBfLOVmMmKUj/65Rl82alCc
ydSMQMWr4UB0waCfqfdO37CRjFeDc+aq/DodwwEyjWEKYnotwTx7l5HcyKas1tn2tb+XXT3bR0dw
MYt3nX7jF+Ujok1vd4o7+id1PPw00YzIOsTANZA873qY7vvKe3+lASuzRFLyMPjPu+/MPsB/G+O2
kLrqF5r+cg6KdQi5Arx4oCvLuB3VQO0BE8fg5aQMQAEf015E7Tpgd6V4rNk5K9zYZtiQ0zk6tByH
oGnqetKy5ZeEdlpxkaH4T2xggCdZNwR5KFEdNZ1qeq9IBmNEPapXR9vA4oBhO/+OjfIk88/0IOg+
skLL8VzMq9dAjXjkbU6edlvRgkpbDEoofjDEeSgxjI3Im/BOi1BvhfAp/cUgCRIA22qEwbF2i50X
1es69VBT4YJni1lx+2CKS5UNyZ1vdVV+xlvL2/QGXTco5jHWtm+u+54fruvNCUY6ouvZJfadwqEW
6UkRwHOv57zYwl65oQcwwFbYc2BnWoJ+KhuKP0yyjCLWhc2XCvbJWGVpx1GGa+vf0rSQy+nUv/Eg
WfEwrUQlgl814PdzQqf9XDU3iC4/klT8Grr8ARv5QAcWUi4rhbU3/ByPRjbQLelTD8aV2iZwMxTP
BLFSVpToTT7bSa+OuXxxmlSdgtjKhHNNmrrn3PVbYLX75bV8Ro8EAdzIML2x+3+hHfV8HtKzlcTP
bevyaveRlEtvf2l3ev4k0E61lZGmypAel6qlhXzDoaRYCdzAY8EPaRtYF9Ox4oyoes9vgZ85iRKR
/bK/rrMGD821wusTF46cPHj7tjF+0d+VJKWbK18GPHGLojGm/AUbGlDN+YEAwQ/P4rSggGvJYNeW
DgdxK8lmpIcB2HrEIEbqgHdPYnLuMaRdmwPxTaOjogbS6UMERp/R7kWYergw5JlENit7n/NvTcNJ
Y8etebM0R/qESyEGBNCAdeppB2BU1Op82RBKU+RaIqF6vlXfYjxBJItX9w33DM5hzluYq/qO0u1q
jpLboR6PsZkkZMWWFLKLsarepYS55fKwKa5IqSUFec1KVna+662d4CrZi9Zlz3Zsl7SyGUh+aG6u
7MluLTsYX2WrGhJWaH3Yx+gp1SPq3FF+kSHml7DTYLk6A5rTFtyumDWYEkP1KoeWFQp64pu0pET9
j7mUn5fnjokzM+7Diu+I0CgaP+X9vTD5M+QHRIauz8V8AMeQvc4l6XYJN068dhf5w/QA/+tzqI0t
Y7/yvLhhtqAgLwZ8X0vU6D2mtw7I6IvbwNBMxftPymupNEX48VPmzoG4Ho00GLdc9mpcqoJ28cVQ
j76VQjvmGwcdT9jcSe4iqunWmWzFEHgksROu/Qwwr5PE+lzSb2XiZ+Ge76mOg0E1fvhfaAhw0QwX
oPu0GjsJsO5Jmx/glS52QyB09wSZZNclHOAOjJj+6YwgBc1yXF3C2YF6DMGMMMCKi8TL27ZOdp9L
H0nT4pzBkLr1uOdtBi/Gg9n/sv744yDSq+UrIqDS5bKvoxk6r0so91iSvRFkd8Kx/wggFmP0FANx
sWt5Z9JT8X8UPx+cMSaj0LoyHE0EF1HH1RaiICl+8Hn9SKD4XpDkZc41LcwTEJvXT70H9eFG2Vrs
ex993T7w0tY9RGj5qYzWCaXfspjX8mE4iWOr5a9LjV9QRs7Mo6LVqt+xmPssniNAnqJz3U05lAeF
h5WAdjrZKeyrPA6X9Exnk0x+fGDNpIXfncp4z+uz/5Fd8aU5+cDZMVLv8jRjIxWK8XQba9TXQQyW
zkmQedhKjR2QcDyH/Lgc93XaWDVacVkBMmWFOihWNGk9APmhxfygivQ6FQLGEqZqOlfI5H4R1zun
6+oyvQtSmdHY/h5HXehsmNtIoKmopWD+y6QpXlFvdEWLZ34pmRsswaWFZEefYsV0G1ni7iBxszNa
J0GDxTq5zhzrjNv6Jd+gyeOcnae0ule/JTpKpqC/8+YErWqv/jv9JeKm2pGg4/LWR4i8VMNRjGaU
gURm1gykCe7A53/aa0/vIiCi4edlSDo1fpC7HAmcnrRfYG7mccr54mdOkf7rAdxMOD0AEm6bidlI
7gNF1duNwMDjEdN8/rqCsCh0ZIhAwr1serMVypYEHnx1XESRer3sSNDmaR1HygxYTyKVjCgcFBPg
21TlAujqdEwSByeZW+pwa2ArKnd3pE0innpRIeHAJU5U7dD3XJ/GfUoUOFbLQIVF5VXg4bznc0DD
y47UJMFw0GHImzhXkFG2FOh3Xnq0IBGWFqv2SohaB2i5hjlZgnzq7Cs41516h9wS5rmdjjTdORU/
CcMcW8AIGZ01A49pB0BFj8gCEpErl2VG7/vyW0JPmA/bm/nJrgQr921HcZEFaKG2esC7ey6YxH1k
rq8bKRoIorisSucd7voorqTKzqctov+KoDIZtCxeh4b+NdmHyVoRyoesQMO2aXNWNw9qOd8cgrDw
atn8mJsyYwtSVmbALBrF159QXLBcYagInyuTn6hKzpMfp7vV7RzZwK3qxH6wZ0Pn8THJ4iJh5DqQ
+EuKhlm+l9zib/6zCoS6tS5M0GdIpJqMsgws/EtdwnAApaLWNfbV6o0lDHBifRbVLHzAAoMWVHY4
hnIEzAK8agP09/Cfsc0mvp/TPpfB+eZCFuopowYx0JgJNDpNaaf4rnYGXLlSG8nH/kQtAvfA4/qR
bmYFxm5DeZ/ArMvJZh952GTJSUxkn0gZ41pGaq4WnWcg1frv1kDztlmzT4sJWLRLu0TMsZ6ricGY
iKtnIOK4C/wJhviHX/FQixcFmC4DNt9ZKHdtFCu0jbC+tSUyJSTDwHYPAznZEEAPESCfJ3pyDyPI
e1Riicvuxc4FHaHEhCw5x10RrnKEZYSHfarNLOd4m8io4Lan4pUntLhluE3v2kKsXZRoXcXVUMfv
K5z+GhHdH40gsRGqfB23gRNVWSiMz53ldcaqeiz2ctVrrCAMXtKqYMPMEPEZamG6jZF0Pdh6qrCf
yYlYgYnSzFyN+wh5rBUu+3woYfVsbY6UsJtrps02T/4dIo4tDVcYe638iINsK4k7eWehlUrD24v+
zZsN7TbxU9c12cMMcC5qK/wFSGDCi+Y5eaCQXZtF17yJfqM/9+RJnNPFsc/EYDuhtvq+jixESbTw
ofA0YgTUl9jc9PulJDc3CMTQkVIwwPtI+AZlM9eWvEdyjz43zTSJwKS2djEBeKl0PX5BBBqjAme3
JurvJeundn6WAJchX4wEEWV4PL0+ok1V80nkfpUEMJJfr8mc8ea7fMQ9Bus+Hdn4fzx1Y5xyyax1
ym1TvdkTC6A0ajFfW7LuQze2eiqlsEen9Y1UdV1+LNORgv8heae1xo0QbwixDNqwkS6wcKrr489X
o5L99ZaIVpzDgxfDolX/Z9QPW1RgqlG3IMEWJt8r8GA+oi7gyV8IWJ+9N+Ubx8XRGjRtYys10oXc
r88NZG/NDhSmI9suH7JMqIMNih82MWIzAtO9OlXQUzJio9pBYFsD1olv2PNoZ9w0VbflcJf1ZtC8
bnj8brAuuoDwjCfl8w4JZhaa6xhxIq1Ah4ItbHM9b19CismoiVaFXf9rtC+DRZ3HGuDu6uv3wsju
EkTYeOGwvc16j2Achptw7fLkamhP6VTaF/Vad2tqbLknRewwDdgVGgjLxz6S3r5Wa+ypBdBJS+p/
DnNU7xeS87yno8VnnebiQAj3PQzO4C0hsDo4NCFhJ+eBKMK75bUJwp+FSuZx8hwmsTL6I8PGiCtU
mcNFAf3bBcvBK2nfCVAigsOMg5LxGiEosXH91KjsecvNocn/buSdcBW7ZJJAg3ffAZ9Xb74la1Us
PT5UAuZwghBmpSch5L0R2LNWNn2C7LJMbkQv3xHcOFrUCqu8E294fmzdC8avpP/cBiT8l7aq3Rdx
9eWyYrx8lOfY8FXZcO2HF80hCP+mARX1yUFaoqRrJF9qufhB1qxJyZNQ3I2PQB/JR2zWj17H05YG
hUM6hGwAEPDOds74Wjhj0L8A6UDHc3nyYgRs6IFC8dLGI/u1JPSImbKfMzNWMNpaanU7DZDeVH32
bOwcseUQMBqbb0uo6hlJ/5EguvcH2UZAL8/0BOE9gBM+RfD320q6aQH49tyjWD8TsxfnGMso8THH
zK+7FGdUTWHC9HLzpcAYpl4IwA4e9MYYm4HFJU13wlcNGqv4Y0NPpVqNySeq9hPljx2IB8bvz74I
3Qxt/oZ0/DD0UpnuZ+YibNdkVwfpyFa/Qag/9gLSDZacMlX5t7YReOWIX1dj4rs5PaRDPfJoocOw
fQRYTaeC1n28EwbEA0TyCJkpj6v8b/ZDMngT3M7bZO+WL43yr7zimX+3krS8U6kWh9v6cgIKKfAH
x8qo4j4ahHwZH3WWEhcriP78YjkHNNwqaWFb5Kjl8sokRxGSsHKyECEOGrzgLkY37geXQlnU8xOy
HAvAE0d1HkqQYiWt7UB9PrsMuSCfQra73apUeguMMgJ4fNVhAB1TZ0We9wHOeQxS3xLp5dSqC7dM
UNh6zlqW9N+vy9hgs6kKlVR4uL1e5Od3oL9C4Z0fIp8seC0tkyPZTYDmZ00Q7xflXGK1TaRNMJh7
HFJAppIQgUUiVGrvpVBlZzZCpDNdOBLqHG7GXVqr7ShCT0tOVY+KuSKpzVzP27KMOS5Al61x0h81
4ssdkp4FwxdasXijtUhjMbSVp/mAp3R+8clXlIvPbNeE5ERlSj+Tzy0yPBeajRTbvsVt13/2Pi84
s+Emq2T5qEeW+kvGWcjSN822HSnmgKAiSNkqSBi67W2wLiCzrxqEXN1bms7Nw7MsKzyZ3q0uBP1F
83fWkD72Mtzo2PXiDWnUMZPCHkGYzZh7t9DBg49G+cUThQUPGnozuXCWLqPzDqyozC9ZJOD/GCfx
BdB2CJvcQKXQ9nfpaQHq63FTVH7XiNdC4ai2TsNluBxYgX/aRU8k+HDt38VfwwLjIXKHQnHenjum
spfakgzu4ulocVi0cmBZk7BktiAG3w7E8Gb7deASyq2tI0kG3SXnh3qVVd3CP+ETy8g8/2+3Dzg/
+sLcPc3A6qESNKJ4aPs9MePip4MGW2qBLHI12bnXPG1T2sdkrHrtFm/sPNP6QO5TTi4Rc++1VQyw
SjhRQItEGq6iX5ysLSutWKl8A/kiyNcvtfsWceXwWU7PaGRSuKmpBbcxQU+i/f40byEMBLqkkcFn
8aCvFMK1YKznePmNEG/ts438ZZmYjmtUvhzUAKaFuqyVDfz+/bpDEmRzWnEpTJIMkYPmCDGnXNCY
ovbXMFfdc58cSiMIxzOB6RBQOFnLNcbHCv05tUAGo/n86TagVdYpihqfGLDD61/NOoZ4Isq3Ax0R
8zDLahGMzMtxtbps9z5bxzrGa3GYXiDN2lOCISRpqDsxsPkoiJNeNDoLk1wrnKrYS1Pt4vyzZ0LF
S/3O2OmuBPBfXtnOhtETCrTc3OLnfdlcqot5/V6kq34j3WiKIUuBc6KZWQNOiJHZ8ZEmRsE/7n2a
j7IoXsik3ZAjK2zBzL5yOZw+jxmJNzYFIe50u+X1NyEduF8YcbbL9N9JL4XzbOYYEioYRojS3HJg
f2sRdWhZ2O5A8MWj0JONLEDGYfvzBnZ21soKG9AzMZ9sM6usyZ4rz72oLVC75m3qe3pYjO7mFZCg
4FV8xfBYOsHT+YxfFOHSmGkIYIPtqwesgAnFzMJ3gpKoI9Dp/8xvGEuPdM/sQ/yiife5NA6F3kZp
Z6hwz+q4O0gtsmvFuM8NJ1YeluDSWBhfSnhv2sebw2I4fe6SfRLCswROgWiGdjzWwFbCq/Xn3EHM
6Z4FzBsYcA2/hMH/QJOCBOCWoljTzviTm2uzD3ib7EpzlmsR5u19S/Fn7EYDVEa+VeIfIov6ek3H
ranT+WMYtzWlJooKumYH5o0PBNcKdF4npHeG55hV6Qph2SN/WplUxEdAUA2zbPOz+cCRkAg3nUkr
Gi+054l3L2nPH97iLxXRiXaushunKV2vUKxVr+U6fHLnR6Nx0Eg6mOaE2016Vijtor2UTpKO/15G
OmsPxev5+4XxL4lsuzy5vra828jsN/h25WbDaayZode5RQhbzXlo7LPwAF4LIUDDQ9dl0SLkwkDp
csWhomIh8aFwUsQGzdXeoAlj5Nts1uWm0YJlbCJEhEBCIa7YEgrqN6iLNDxejw8+rWvMQRJkQDqb
dO4BIjWxuzK/tlb/TUmgJB5tccsdK1uepbONi2zCr3MT9Jo65QXrGMpJ/mMeUBiZ+tmOjK4P8oqz
6hPA6NKSaE2jMm7rxgYDA0R8WB+xFJrh3KvL5ye+FXBFDj/Ek1/qaFerlzEvvEAXruIaiOFO5hMZ
L1UkfBAgAXKkh29B/JB0+KdOCGlDz8hf2ipZSZFy3WomapjWkF12ZgQHyWPR7/LO3Kp/x+evn3vg
eY9nrA63N23Hc6d7u7pq+/OQxLKw17x+fXiqh96xnFVVq84BZy3aA+wisTVC6/m9L8F0Gu5msYjt
CW0eatGCXQQP1TU15uAHwYTwcI9E/4UTMbOX+qzheqnRDpMHIcjnJ2ui8ipLv8a+gB4lkHFKpdO7
aRX4rzttHTVyiDOy/A5C7MxvWv4r59ZLTziYDETlOstpQB7FQdy+rN7XQHZQ7dmzKOxS0H13VeoA
YsKrzGs3IJDiKfy6En+qwqVMVXFcgckCorcXRbTxACfD9BSZWAmaNTj0TYH07v+jOzdcLfK8LbyZ
q/diBSqa3gzTTHLOUoSEcmlBqCRRlcuJE0a282puG98GixTrrPsHpQ4JyUCHZOPz1UoRsB6lbKFZ
q0zSG5Ro23Bb0dItAcfSaWZ/qf0i+Qk4l7+NEU9feTV2VtctOEfyj+JExeMjhcy3H/8hO21PGkz2
JXHvnn3SJdt9RWgXzeZVY2jY1w9B538JRfznWisXr7PGRw5TMbZ2hPh2GKZxczKSFxH3E37Ge2aY
9fKyGNU9AndEfXc0twgyCFpJNcXm1nwBNxgPv1UBsrrkXVEE8Y4jMhK/bkG6Q3on1fF5G38BdKxC
3Ui4BIZhpf91w43jQWMw0MsNaILHtwj+DqE2qn87stb0RixymHDI7fj/G9zd4981FmW0IdENVP7K
tx/6MFPUg2uMdelRCuyZ7VoPDnld+b4w3VObw1qPBDIMwm7cv7FvlhBG41Qy3Xi8s0gCWqTqrshD
eUWm/jy+1eVqFbmlkT5x20U2XaWibsFnzskq1iv9Z6YizQ+799iLqJxQ4zCW2q3/mTRKvbQyUCGZ
cOjECihLOzgRQH0XojKfBqrMBnS0wEgfBNUqMSpfUDoaKrUQr18LiYYLmeoTD/kNLIxcpvtdRPt5
XR/eiQHGpCpzXmcpc1o61lAdDa+lvQPjiMSSG6SMP1YRccuOXEGdeEabxiP6Jsrhh9G5bmzFJizJ
3JW9kr7xYJGp4K9Q3FhqNOvmGkXAPzP+7UjnfrUivMOaMg+5NUhFJziXVdkMAKslOdFSbN/7SKxG
jCPnD+fTgBZzHoauFE7A2F7xXnE1/59YfVVEuzI+x3jOXqPuEgpP4TPpjk/v0bdv+S3O++oAwd+0
LyGqTxyx8qbnZLgKZfDB/1q9nZq1hof71m9XB1dnxfrBRqHfZsBkFhQ4vkFj96rzWKICPoAn3SXT
he66o9UfgPeJ+xif6FMVny0ktfnRrNSOunQffB2zn2umDX/mJatJ5OXpQN3yw21IwufYdO1jXimt
vvAOUWpaWLbv3VWUD82HkZkgx32FT9IWqJ3olBl8ifOMejT14odIvbV7mZvOo+PIjEoxQjmyB04r
duUCbViU8JB2UjI0u56JrcAIBiPsj40IfiM9U9XnghFsnNzaUbnpKsaPMvW3cObDhX06K0FctWlj
ViUCxAJWteNzLfqFcX6eWHM/jQazP6TNSr/MHHf4sGgKJ4TPP/EUuvXZdQXr7Kkz+GvgHOVUG/o+
BpOvtGA/JJAiSY1AtUdiJ9BQ1HNNmI2yCmgHl1B61qsvOKsx5J4ZOaXhztu0gsbfz33/cs9bg67N
yc9tl5yt0X3TGXbtRrPumwZ4WxTEfcs1KL7VA4dg1YedqUBJH2/fD+xpg0L4TcWK1q0PE81QcAQ1
rW0OwAuUnh+wsP6KYSbmInTf03jJg9vfvxNPLFFY20RogZXR97I/vZIJ/8FeA9VO55sLw3rje2qG
TgjhvHCRjaybTm+9w1ISF+MRLE3RGId5k6wg3y+Pu3WDa7w4p9Vq7YZFVvnRZ3DgpgeBoyGMUPCe
RlA6v2aA5Gscb9amIKm8hb75pZ7vUZTzRqsFb4iZotziz9vAHDDIdyWRP7ou/1QH/mX5zfINwB4D
Pdj1mOH1qEKwYF+V6iHmOkpgslMBZfi87DrmHKUQJ+eZtbAZiJUft9O7GisROzX7kgZQbUtiIjAt
BmlQpa+GQ3sIH8hhxaB5DTezTp9XBml92fBtRaml2P9HaX7lQsaX3vDuiGvuauug2yxEo63rvekf
9Rc5zHaXSzqLBByTwlGndMdMEx+f5njqTpIPKhy5Bxd9hqvov+MgvizhLdxml8h19tbDmfc9Aj5w
mnZuPQq17SJZuEtlwzGDpGz6RwG4eTp3plRg3F0OUWcOonwZtMYi8y/vlnWP9zNJ0b83WMJuqIuy
RNK0fHGGFlZtGqnxlbdePDYgbXcLvi7QVPwUXSAAb3IgwMjWcFojHhBAytaOvYF9/XDs32cf0QlN
bNewQx4pQbFC3ROJy0AYo2sAjbrGUIcCTOeZ+xawjeiUh/f95tdRcSMUn3c+ptryFrzg7htqc9t1
Phg3RnvcTki2bLLbzhaQ9M0pBSf3E3Bg/5gADhCAS8sGjefA7jOgSAQIu9BDQMmW5ubaNrPQHVDb
3f2XupcqHCEqH5wKPySFmUp/NuX6/XkhICjBPSsj5LJh11Cmc1Uv3w7sZUBX+BMHNxdofRH1yOPl
QovABW+VTFWxgPg84wZSvkj96WJ56TjdcenkxQbBpWzGiu/OTDnwbZxkOwVp1dMgF7U73FrXAp8b
3Ecl8pcO770OUV8NTAouAvXJcKzd3m/b4jKZr/y/llR8B9mjNLE2v743wiHo8olDQ3NwMVocQzBm
2AnjogHsmIcb0mQ362vMnqMWOh2fc662R7/w6CL9RJUr/37FstomVfVp70I738sqeNy+GsEC2Efx
A2YqLu+DUqYLOPgO2jcMtWsQ0tICAA45CMOFwhwPmSKPTppS3vHnl5hX0qJlVPV1b/YaJlVFAwwm
B+H64DHKeZsxSaiMwgO5ptxLUhN5ddtkv835l6YG/h7cGSLdYZRVEFGwfamXHTqnJNMUdPlKL3ju
7EX/yq+MPLok8297AqU7xlb3siEsAVLSyuSMOL+p6q82tuH0DvbklChbstgSbSU94D9WbpblSVrF
X+3Uz8sEKxO6x3GvWqrTz/R0m3RYhngcolP9BmFWIZ1hLudrEmc15WeU2d6STZiC+NikawCJJnnt
lWf4NrzhWZB0JzEubOpMBxXaPTBnzI6Q4L0ArP9wicHESXssXw7rdJlX39rBYpCPtm82e6ZPOis8
PENaAU42+IFduN7d5mdFBZBJBdfueoryHGgEUNOWlYTe68NXQfchCKwNk1YTJCKisxryyDuQws/A
gunECm8LM9dueLKTXXHo7BXEM40oWieThkmtWQWu2jMJnVx1xUJY1j8ddiZuMoQZw5TsiENrSa6f
AdBOUHjCzgwnEg81HYd77mgO3h3v1tczUH1Po3uVpBYvGyTvmJRGe92ak8vWNqdFI+7CurSh69QH
BBNnRQh59d2QyDhLoWclIc4akgutbwaxPtEWV37f3jwjAWI/T+QZt5nhhogO43N4+8VIBt5F2ELm
YzgAmlQczQsmUiAeIDAB7V2wObKc7m+pG4E4dzJ1YENYszaAi8F30YeoXCIva4Tb2PSXRtnuuztA
A2VugeLi9eN3xlikMmvpptgTZw3dlSNtIc310EzLIVi3Z2dXsDrYgLzq300Zgn1KO5jqB0/a3+N7
3qYMYkNh0xywjvkW0cL1WQpSuwYNYBCid/fOHyI+gXxsOHyHTmxXRS/CWqJwoZfmbwZFIY5PU2pg
ii3yIy93uO3bgAAKBNmZEPuJuPagKMPdnh/06+eiGonrJmyPNZLdOwQ5pN9X2FlUYuQ+xwmL80Bz
T3O8KJicNDkXDXxKm0Nyj59q9lWBjftiJujyvnExx4uGenkGCvR7BMNTbvLWtwGNfGSwXXQpdYSZ
sK/oRhK/tXoQh6ZBpl/gD7WrWXG9p6IjmKN6DdBKZRar93nQhO0yxUlClyCZZ/qwj4jmxN9UoBEW
ozbh2MtTlVbkk54oF70afcb2C5Li6cpB4/YrO22ctpIsiPZhN8zeCu8b1X84DYqFJSQgbFoqjS3a
vkkpo8e7KT9wdUKzUMT9SWWXzQ8v6PwiXk6cdgW7W1fKjx+Ym4+dtp08pf92HW6remIC6y1cK1j4
GFR8/GmvM74mMtX0DiqEoace+f6nNtA0+aE5O1H1WgiiVTQl5/5DXuUNKpuxBjp/KSVTptGI1kbh
KrePPaffXS66hcv5wPieHo9695lCc657hqGZEY/l0Vc54NodHL3M0UErKEerpHME6SSRXhRkr//U
4Ij0eE7zrZ3Tu1RysW7Wla1qYU7Bnm2eEIOMdJsckZOiabIj6/6aAB+mVU6cA9F4dtnvqYNJOFq5
kMGAWdNy2zPVqria6WSA7G6AAjaw4ZmJFa94EEX8sRAuO7Wmcx6vfa30oVnu77QN2VaEeiDMlqVL
r6u5HCA0FuZcgUscyXKV1Vo3/DEyYsWKtpgO4TiJxxjDrJhL272ruPOsoDRmZyyMDzh7xixQq3XS
10r5ZcN4QQ6p0XAc6BhAjpo49vPzOMaC5+0uDRttZTBcURH3BE0rEVOggETzy8o5Z0kEzReR2xtk
m+qZCxav4AXOweKCaPwNWKH2/z8GDJzSENcKcNYa/rM5MH/x3bCoU3swOb55FAgRu28R4SPnBHUZ
SxZ3ZY7J+13Dr/KZBkQrTR32ZFMWtmus1GF5M8PGRIU5eni95Dztp+DxpO8GYDGVaSO2c6ry5u4W
fsyN0bUjefCyajghr0aMgbzE/sUzRoHxRx31yY6AWI9wi3pNWg2FI2NVuu+uPwceZA96BuEJZ7g1
oqxKwNHbDclzvD6Ylobtrxw430Bui36XKt2t9ruCEkSeVlrmk8rdnAr7aZy6wmYwN1HJMOOXZXkq
8jyPhwQnhL8qA0YBOr83VN8Q/l0fjVa8EcB8z17MiYpx91OTWP6YVPQN0Gy/DEUFC+wTy+Ttmyhj
sr8ABV8A9Ll16xbDWAufY/MzccAnhCO0fM3LibFV8fPx5x6wFI39O0lVVxXKv9cjWewZQkE8I/kg
zuy8a4Q5i75727750oiYTPNNdJtIzRTJCz+ON1g1Z7ccK52saWCEgWmE3koJItV3U6oS/amV+qaS
5Upr8u4UZ2jKxtUhPjJKsq28hCnIjIwaoehlWEOFk8GZInG11xHYHvS+VrpVA0IZgIM+v1T1VyXC
QkEuS02wzTn+FUbABJ9qjBlHCajEP7GJGpehwCkxqzWpxOZwohTP/IEqKCTwnYqHBkH1PxMFob4o
ijt5C/27jqxzrrTw407BoQUxic55ZFBkNbcirg1RMaerFy8mKc/dn5yDr4cRiyMM3zv7zH7VyZm2
u/emNVtiLovd0sfJGfGavBD2J86/Occb0eSSQtCwgE5oubuz5BvE9xy+tfYrmZJu/aMIzNV0+Isy
BoS02IfdKd5Quz6Oev5mDhYjjSCw0ybBDdh53EvvfAnxy/VFJ7XHf8cUM6AdU14/L5R8SiPBMD7s
s3jQJemjz0yspJBeHlH5Mk2JZGu22gtU0ZnDiDY4EopMChEcTRgzk8/304ChpV4twZkbxp39klLH
8g6ZET9xo+TtMZReHOlkUubi0WbaVHqAjh54eQIgbEIzK276IaWVae9OiYdHkV0OgfC56sEVLaYd
xPKDB32rWyqk03lVpeG8Mvvnq9oct0mI83ouzidKH+IFz7wc9/9YsduE9uJ3ajyv6N2JHonJY5/c
cVLyzciGIncEY/9pIAJgIzMTaGf/u9nkz7EaPqUg0kluJFdL6LOInkYuqqu4LwIXOSNQiR+XsKCa
fSB+5F/YmTCgV1z+gg68j/zanIahFykT5apyIdI27HAROtXEFc4GQpTDfILmrl9h4Fr8ADj75Ba/
cdFLZKiGh7PtZu4YaBkudsMHDo33EV0Dj64+aS73RqKVToJonBeLqJw69AFWPp19YvBZvmT1rHQ0
8S76rcwkhksAX3gcHvHYekh1tR7UZF5aB9jwUBLGtxH6o6O8XACOWDUhXTWASxUT9TU7leQ0YP/f
mMHf4156TZSGbx8JIUaaIGb9T1NqQB2B4SzfO+RdtYjIr3w3CIvcEa35qyC5ilUmqYWKftdWT71S
iAdEn7+QrrVuAmPFYMUi1hVMoKg0597toc6qATkVD+Wc6toEGTiMUB4NWYEvbAeFE+R4n119Umrz
A3HSEFBm6no/aqODYyisJz4dKjfO7z0ncP09EhzjGTozPxWiVhUttIxBDAcCwVFKnCodhgHO+QMC
2SM/fNHqOh68HZu5lV/xY++22RWKhmY5eRGf8Qbj4lVdBVY7e4seswKZrlG5bGDGSVeOuhLKoEs9
5BKq8n4E0o2S1NU6cIBCOaRaOwGtuKgiZfF4d9Fc0CiwnOmiimEKVpNzYs5ftmpKce8O5kgpt0d6
gKczLk3XIddH72QL3YXjIkNIVdatDkqAWzO/05tV6z2eQCmmbJybM7+tzgmXEQdNzqKuVA7D0424
hMRJoRdcIhn3JwKvukwsBoRRBtMAt9lGDsivO12Fgt/yLX4KSYgwDvbpA8QQIVL7/AJ4Cc+v5MDm
ccwKY8Tw75YHZ3Fzb+rx91798QJFwklvtTPfgbgSobyb3DKi2Ts4q6wz637bmjIZlSIcqUL2Nypj
0HgKzCYJI76DgLo7bpxhUjo81wqEjX2OI8pxxfU+N4m//FgHpmnmBFJOJv4zS3xFkgGomk3MAmAe
9fst93cenkWtnCrQ54J/QanbG9H6EMFrZJoYmPC2crJvd72qsFOLGORQVz4Dk4rfVtXnBUOALD9P
FOSpXssu1DYUzInJeUe/KwHAdGg60o5ftlbfwodx7fbcxnFxVSv919vi0u690oGdyEiS9bUSUtS/
6sgD3XjXWrBdc3Uobbl2pkud4VVdTt1CFfABewYIpP7c8ft7lL30E9yyZmKnR6mcmQrOKDxfDreN
jyeB+buDZZmyYkBMU+bRTVY8GmwFZgCn9weEv5w15WzdD8qDEYoncXxmyC9xhLzTwRSXU5OXVlXB
H7xpVpWTUc0YKcXjgycMEtBKv1ppVUEZzFzjLeH7fLsDYC7iXXYaV6BmhuY+S/V4zcfh4T5NWagf
SCw69bhIZrM3J6GxHyL+rs0cZit4TTnvRfhb8RpFJZVKCxJVu2OmWxdIw1NP4ewmpTZLMjrIzShc
PUfESTtoqUw0jXATmMNyJ9R+u4LtVRnK4yJZQIj91ZgCUltFedS/+svub4p2GtwIj3kq4u5ZyG9m
uxdjLJ01649b3hmqssGX2N+8mWc9Ok9SKGQ9YWk1daCE/Tl5ap/f42QL9H35kPMpQKWYYP5yo1it
g+tNda5wurijPSrlsuNscEryPLdG/GfTdF+CixHZeBfWEt9BALseG6mdrFO87ML1LvPscNkfWjyc
jKJ7Q/VM0RIEmhbULlN7dSUSqyivbElHXrjQS3BTWT9Zpx6CPohx9NNe06ltbfUzWKMT3vIXBc8T
v/RSIZrsP5BYmFznkVLrqH6GgfLZPSYseSW45cfMDtYwRnuaxHO4jXHm/bvuZsxmIydGa8tYO+Zq
zGIbZnZTzbJFZsbQtMcCHLinomyEOMiQdvZ7BERWHzwFDucJrn7SWjDcXvad/QcX/o3liQSBUbM3
zeZ6IbQ6Z5LpFaRBrwT76uxj4NiwGhmeeP9SH9+gVDwdw/GR5/CuvrCFqpdvza+nSTCgRq3JFB/+
qHh9TX3PCQdH/bmo3RqJ4fjMQsr2GlTLSdJKpnG38bAHAQe6iM2sNwp4v43qWi/m0nEDJa641/NE
F95/wNkPfFXOPTQbbG8qV3tSdDrrgZHxQUrEmVoIWimTikx54QYwlhIMmJKccUWOya3IRNzlfSc/
P1t/QLLR3zyol+I4rT1xLjjEEx6R4WTRUTHpy+qALPMS6UEKb5mt7IckHIgCYxcT2oU4AcYDKsIF
Ed9DWSMlIx85hrwfA94Oar8f7/u+baxmN/5Y2K2N3s/xYBFJwmb8ASelDQ3v+C084rbwX2hjAQb0
ml0F0rrksKyBkPcdvBFxOl9/FM1uEiaGsjKfToDyWb0MtmoqbKaSdjitamrrvajskzLFon91teuH
U4T8C6rqBNfofU5Wpv/TiqXZp4m8SwkaB7XPALUFZtFN3ZyRUr501Wg2ilEMMS7u/1Qb1ipAW/6q
ie6HiBJidsWjZ+UtI1a09UHbzf6c1Idasgn7WRcqAZETMiij4QFnfKl0HkozQOCLI3D2T1iFv4uY
cZP3rSmivaOC49qtuW9Gl5OHZg5AuaSyendzZovgA2XNCewM7Q2l5DiyndwCc4QLtPnMn58KZwzj
Mc2J2+KO1PsRtSHV1ChWDpdi4z6+EYLgj3qK4Z6uel/60yBkeEhSiNmyeKtYgXe7nRQKeWDIFpFV
/2rwIl4dJAqSj9E3dfxm8hGRkVIJCwFOXQVcKk6YnOP+UPwefdDnczDasAgcgXIOyAq1avDROH83
fonJXpidiFO1z60FDq5iN/wMCmAOO0Bajmo+adcICJyTf08Z7/MKu5ZlH5/DPaTdgthbLo1shYxu
bw6g2ysLzJtzplEQ9wtTjmFxnKa3i6q5FmqqzfRcqrcxc2uyE+uvU6Wh+Z6r9WzLtIlCYevBNFy9
0vMteY+K0liCMdNAtKkbkR3h7KTo7CoLTZsPkOIZlQTRxgvaiq74asl8hXFYwxTeKyeUXPkMfH6x
Uupf6mSTGdUuF/fC6TpRnDzMhg35m4++Rv5u1Un4ylbvMQbcG6jsPr8Irds3k+CMa74kY90nKFID
7r9wo8/JqWbxsGEvzwqsO1QSMZQrg2yh6m8bq1g6eqzt7hB7CRxOmX/3sFsQmuUYU0/p0lhorxul
GGhpE/WqmW15fE+nfi1+dwJtvpOXuIZkHau5sZn/BEG+5SA2b8WgJnv39JFqOXASyHUFQPJ5sNdL
EvWLi1nHiuMX/Vv1fsUgtJC4grLmni8FbzCQaeZWUoBmEW9iRiYrdBEMuXHs8iXKHq888MR2PPns
qEkzlkXYHqaWvkdEqu1ml/4pYTO2TR1xgv2PAMeOYjYt5QbpAT2tozZeYOE7uwf3YkeBHOHy03Sk
2X2pG28avik3EfYmJu9BZNP672y7BZ0M4yABZbHEhLeg5y8fhfUaoGTMU/XT1sLQoEoapXP0LFPf
8qz+XN0KK4zbaWApVM0MZhkHLlhfCjhWBO3Fb6aG9DiBkvMCYB39F1+wf8tt0o11XCcHpB/uGtV6
6plU8r3+csVoZwSMtuMvZXFetV5q0bg4CDRhuuFktDNKLuH3yEIV1+zPngqU9BqDxByFz0W/bFVY
iZ+/s4bBkTZJ+FZ9VmrUBJAWw0P60KVNIRSeApkdjFtlucCxMMtHPs0DlqBLRQIEqhzYlhHOtEDk
pk9Iv1OictfmZlfHCECYV8V0B3z0KNl8nRGf0Ty21Tp800raJ9N5VZSRYPUZtUqv12Gzef0k9FaW
OKHnd5EBfBLpMg08jH87fsoc79m8M2HIIHM2Q3Xg0s1HyrDKWs4fK6+dwq8q6b8l6a9+Sxy8le3y
90V95piwbNhCBhK0YyhA+h6NblWf292BLY7ZAvWvg6BorhL8ipNyXyFS1Tx2HFy4lVxVOc5BkJWs
xGW5sAny9k1JCpn4vr+rnKoUfse9pBIUKSQZyZC1m5Wimj9TfUsKLL49quNAixziM3H/EYwz+OBw
hNH4PaTeKAPzvZw1aYIkdFK5ZV5+1qbs3QgAF/FgbmkB4M/a3iFCGJmfd4RHH9fGqvQazPH4+yQD
03ED4WsdBCjwQinPEfDqJC61/QV3mmDrS7du+lWJr5vJuQEbAoD7JFXTFqREsSBrT78gK1Sx8zxM
2fuCAbEcKm6UaRe/rpXETcIz6s84HU1fTlxryGh7Jxs4UCDn/glUMgByJQ6ZZ/KVQ8IN4OLDzPpa
5Epm323WMtN5tvUOc1bw9ASfGI0PUfCi94riMjznKYEHRzZ+dZQ2j71mHGl3EYQ6pNcY30mE90SB
1R3skLX1lNhXOivO12y4o7+Vmcd8gWlM7iioa8TwBFdY98ZXJEnDWe8InsIT4HFu4egbE73M+Rl5
9wwmnf4d+3f70WoGZLl3CNtgK+w0jO4DMkeLbRyMRzLkUWU7/Jr0ojWga44LND2wdnGAZ/n1iRKH
qpoBFDZjw35M05runs+34DcJvm7TbxU5Z7BNMWlY0efmttMjTcQsTa8cF+Opq6wC/zRWLAdTW9gK
8rFbPYMnye1mZOCQGPIbiSrlwufEka1A2IFK7Yhu8+0hZuL/6mM0WBMDqFxMMKUIQyKK+ytBH3fy
j71QEGoV4pPh2ZbCSpftNvwRuSkwZ4viVHv+iMHudWglqBjAeBPGh3N7MqG09f4AwVo0J8nSm5lu
5Xoekiy+aP/XbI2qaYdx8odCJDL4stNYzE0/UOHRKec1dKmjOCS4V+kIDPLqX5boIsOg9ewuV/VP
DVDrfooqYL1euXZFqjzgAMDobb+slXP/0vmNci1wcN5Ke/fAdqgUyVkd0LHkUgu/OUXHf60BBxj3
GP/2bXD8o7lTSY+kwrG+8qWE16hXeKcRj3Of2KpRGwXbAW4rMW7ACVWq+1r0zd7gcHxIBDj29cij
tfA0n/quIBJ0ZG20EnoaHdWVh9OxTsTpHJ6c1kp2VzflqP3il99GUUxWKlqKsGD+7XShG11RNJn6
2ND5KA7JAuZYZpdPxLITUiLCajkZl2MHVvO8OGKmCEDHWRw8ONsoOrV8ABi0ykYpnEb02956HVRU
OOcl06MThgp1dsu/eJNlGJoAp+bXCQXvCs5lpLsTPWjdfK+rBJATte6L11aOWBCcZtSG8luRGeKu
4Zn4TjTWfZ0f5XoLv5+q1TRyXMks8AgRlVdpYFDW7l4/7WMpAjjSR7RHgHj+AEp6lflHezY/sdxv
OMv5XCw6+PoOCQbUxUNElPothHog009mACLSQ4wl998IbNYPFVOWTlg7JH+d2KeZ5pw0KBftoD9c
QORwMwttJcYy+8pcsDW7K84mk+IO4MzwNiBLS2KLKiB+SZirHb18V5EDzlxEK8KNvIUBibN+L5G5
5GOr+Gy5YNBS9zsDlcUMuzennybRSS4SSGDgJp7H/t3MctqOC7Er1aQj1zhV/dbzqFIuo/oplPlk
qKHLgJdKlbo4zf5crjhanHlJCdqDa1O5P0lwSu6D5qHV51FU9HtPaN5b4UjhNvzmArwS+GlKGabR
rKXiVl93n6afPmRSfDwQlp/jI3oJ2YB3jYZ1vcrG5f/nZgV6F065KEHn3Ti/BSuj6Bi+U3hrW+je
hHMuQq0KpLADlYT+3SK0Vel8SoDLzU4kqoiyKk6sO2BW+UG50uf4teW8tTS5xvB8ZHjaUhV9pbjz
m0QiTM9IwoY8fyEGHXxu5f3/SvrjDtjv0id5oDddPkFbizkxPaSBZXUHnDZ58fz69YuZSb2zEXQG
CY5GUySjtFQyshBNZudle2RjX8Xkzif1saFg0LfkfSDeadFn1+x/xKy/cWZ06UmtfL6zxEQYX/9Z
BQy15/L9oJamGYzW/hsbSUhjOV68IuOsdd23hYKT3aqgaJDyU4OqXS7ldYXHMGmUCTqJ7GJL8yq5
PGwYDXlb+e40Imhhw8wnZ+E3VzREfKGEQ1Ln2CM8SMVbTTBQyGJgKb+qsJUyrGMp7sQBjnrYvZN5
/SH+IOeqO0vkVh+/EKgqww5a6Min7h318B0n8IuWhlOT1V8mj+Agj5uvP4i/eNkIEIlQulbIHFTw
Zxrl7NgoQuxM1PfV5QPqkMPq+bbTsBgKzeYiubMlcEocVRJfo/Lu4rAvNUP1DuC2+XUYG5H7REiw
/lqUfuZeEoQwwT8530/pSKMTjqoRyN5OlDmLt5AN8bARXJOunJCw6dCAzydjnbu+ZgrZ/N3sKbmE
f7i+W3XNQhOYQXHjoEpBpgZB2F1fDxRT2E5gkRMWYYQEMauYkCYAa+2ABaceRIAriDNpwlNlZ5au
+vbZ+EWmD5wSW2ogpJVa5KJjXE4iQdHnuBoYY3KB1KS/9n+U7U/KaXYVhBy1ABvhCyTgDfL7Oo6B
b92tg5VgWMvur4JCBrUrKlJNLsAOZtdtF2zBxqHMsBGDd/xAqV2VqPJeJ+LLbkT42bnBB+gqw56l
L8E2LiFf/wzSeBpDCMAx/SixibhlmLzzGpZGdMG50OseI90Tf8ZnZi796iPa+xFXLxj+hydkl1GV
dGS1LqQNe35op2rhW4+iKcxbf8tTymsRBKIocwe4+ZmroDfpjiJyKv9hkCn6rbSo9b2QUO/SUpVC
0CYpnH0BY6qorif8qIue03E9zSDggSBNyqztxD38nlE5SA07XZ02+HAECT4LBpRy80S47kcvG+rE
Nbed7Uc+4xzHVsfUfnm2fYNFQkq790vcKGyOHGvfhlJ63midViVqzKmebM/GoT07+H+ZgGcib70+
FUtLg5wWqH8CQeJuxfyBQEnEXu8GsBfv3GC+eKYi1TjtCyPRREmVqwpGgUuMuB/IVEcMEMqxcmcQ
HiY6I7lxXFDk65urrzWN9NpOmomM9NTEzZO+DIx3VIcdlehx+sh8wtnkYCvfapM8tHelfzER3YD8
b+xWGrWFxMbbtb3Zqffa8Md/nwvT3jDMKgFEqBuFepc6x8skDbtbtduPe6MMDp4Gy2SeYs6LISd5
LO5EGyIRudpRG7mD92+788d0gZ7+XdLFBXV121wlSCKYQ6qsPHZJagZraLSc+BwkRcEE5OjujV5h
wpyxfTp0dLX8xdSu8t3laQeXrfT/xkzsXEYJPGev4eSNJ8WciE/3FPMA+YuYeICS3un2VXdIEm2a
zb6XYUJDu32VMFM85evU9bG7yPvCgQtMMce9xJbHI9AhpOIqNxa/roLZiCZPtx4i86SH7K6k+x3t
O5iOF+l0KPYDQjbox1Q+ffevkczmpjwka7dVvT7QXUuTlW3LF/mS9CTu5iT8g3hcw6WHm3z7YeGd
CSLqfHrci0AqvPqZQLHuRMM7TmlxZLrfUReR157CDGTvcBHWJHt/CMSxTsTllulkIFDhds/YHZND
1N7vrg2mYbkdW1DI4PGLrBREuccx/QnT9wtAFbyLBvXnJzkdyEeSaiiNXEYSqa1wT7ZluD3MhiB1
b0cvpsaC0K35jwYdtd7Nhu+4R+wG26vQK8OGYJ25l1nJaqPH1EB9yEqK6ZbuOPW51BawdE0LaExr
B28PyDZqkfG27XQCmF+DG5oEUeZHkQdlTXtd6sxf+FhtbyfY/dRaAEZVpnblXW+a72MwSUE512Fo
AjeYQiuUWpmSEiMk4omsUMH1mieJw77wYl+jz0DD2TIvmY86kXLUIpoi0kcJpdxZ87C+qid+be3Z
dd+AG8xk3Z0nvC/B0ts+4NZU9A1yUQt8Rl2C96CAkXhl9LeVvUl0qPF0iUdNFCoyuqTzpdsYDoL6
5OS8T/ACnWFtT7C16gHc33L9J5b6mEBE29gJRRARoU7E77GLpVrkalGe0/8zI4qO+beNHlcT7ghQ
RCuLyd2qzKiWkdLOHfdvE2Go67x8ekqDYMptRj4L7b95hvcx+Vy8ziooBxgV88CYp6YFGbfnUslq
pL5wUw3z8bugy2WOkgGl4+Chg0MYAFp7IQpdO/2hTyeBCaavLRxAXWyd3P3mGmkZLP/xtDVEiGL7
yyT6SjDg9nvI/2geSgPlefoDm+5g8laX++lkSBImcfulKFqk8Tnk4uwpxoHue21fb+hvPiFfxvod
WUVj1k03zV5uq/so15iu4lTVzI36+ui4pyVyFdz+SIHOyuDALZ0PbuWaN1hp4y6uKGQrYd+S+GVS
T/VNZroBsjXlFc3XLrvevTDDk+cfPi4NaKD5O92dg8yqyAr4W5NB13lG822iiPHxz13R7mPpZ75a
3J8wZbAT5ru2Mra4A6Y9ZoCKWw8WRaHgmASHoNSq3C6AevszJEub4/ky7MwlU5y8PxIEu6Z1FB8T
RAyXNHclCvpbHOC0cjZ/6rOjwoACSxaMCJmA5mx+pkOCVls5SGc0/8pWYP28y/VaMglnR+TbbCl1
6a5NUyTxsL78QH/TLcllTbjzz5TT1mecqUK5JSRItUXw9gWCwZBSDONJfsuwX0PDKVKKO/KtBGyz
oVDZRAq7My0M7A17si+B83ooAjxBvQ6k6mo8p/wQVrlM49KJRAFJGwX5xuQUTAQcWXI7PGp8Khqt
7ODvalICB/mNd4jUyyGyL6cqYVUCFw+LQ5K9InkJAmDiM2lXIuPrl3Y/yoDaiqspzCSdnMAntUAr
0VdKdxYp+Uim/XtZIbIw0hODaR0ihY2FB8gkGoUI0KKBESXTX1gVfw91d0VdDHsb+wZsDdaJ4OyS
T5C2Bgy3TYVWJ6nLCIv85/McBWnavWxTTOT/wu/nbh8MevI7y6ZMNjBk3+1N2p8GbKEKqQR+AV39
j6h89dySn4ZhqqZp/yAqEgax0FUYPrwnOMN2TlSTSHU6oJdMbSVOVHl2aWHg3wbGAyxxLe21pv8L
o9htfE8+VBFFTh0AAdE1KOVE2stiPrCMHsU/p6Fto7DxmKi2Z8DSt/173v1npD7PQyLN2OHEbz18
s78EGouM8HjuMNsoyEYzs8yqLnwvEOmqv+mkT7xd2SgPEowaZ3mZ61X/BLOYxfTxDQ+FkPr4+FhS
2rU/lXLOMduF4p/MJvgf+Fl8NJIzQ2jzusxRX7k+1O3ygdb6oO7xbXWN0S2jqNMHcI0ekNOcyNu+
QaZHnrI2DNDPwY4Pun0jl5QPcTV7uAj5Og1yEh4wnJLivXOYm2IZQyvdHkYuDAjJ3xUBaAaqfwUd
353Espnuj+i3hWETT4I9L8iXe2pLw16Si29aL2KddLg9fWk8s2z6cLacBVz4ahmj9P7bReaqO2S6
i7SRlBsD7DV4IlZMhAopAsmMcgFd47Zo8WX5QK8rqnebyqk8dphhe44W7i2/RXU0//cIjmf/kcqS
436kFIquhum91U/vm6nYICLpR1yd4X/FBd44IsHqm+Tmq3CpXLqprm1M2sxUkGGH7PuXdAmoXsVv
d1cWCJYfyyt6JChBL8oKGfD6hKuAf7GiDrYvP8snXAw3CPAEmOsVVLJEcokuL6oRtiIsSvebqVE8
1WJKrwDJeLlI227qAPFZx+U1OfOWrYNRccAFJHiN6jjJvKEwYKLKsWcrK5RALXmJUWe0s1mxNngJ
MONZD8D0lGSgaSjsIWvwTBpZPy7ejiPqs//TsWFXr3fElP4+pHkpi1vhqFhVb9VMOouZ3afX7kBJ
0fdoYWCnK/vJZy3srJC834pLV0xvUQxWeaC1JqEhajwOTNwCy7PtE+eqWz+fCoia3xXMVksO9kER
Z3F5bJ+RciX1whKBu0T6B/XZ5YgrVqmm22tjjw9oA5rKqyrtWlTtR1F477yVrJ1uHwCN7iL4ds7p
j1BJb3q7nNSZTxn69A36+9/F325bUtf68xXS84u4o/CkexS5XXDgsFsaL73ABxmDVJxbEvDA4WxC
XSTL8EM9BgmpPmJ/+tCX0ARdhEVzHzzfNbJKopDfMXSPTY2Qs/kl0ca8gTXYbQ8HT7aesBDTvu8c
7qHdk6M2ig6uWRc0AwSJQkl2wWqhenfmk6P/z5z/Zh83uwcrD3Bx95NhVYCEPn9FdVELIoeMmfsi
i25HZduyvkgPBCwX70CSc0CNrCPWZN1Ci8Wg7pR65/pN6iKxaEV0hNXISjfAaSN1k0OAQA9FQRHe
aOaKEP9zLo9d6eCJUzVLbi0Zqjoz0oA7Q143iv7dZUES2HPDP9bNo1BfsTi7vmdN+2jx8kikJ7v+
EBD6D9vwfrMoSseci91kbnTBka4gqd4OonbYzAhJI23ZPPJ1vO+XCe9QDTy3mHeC/fEA7RDpr0dQ
dU5Z//8wjFYTaU9yB3azBUBIwxsQKCfsbrPkyzIF9i1sjsWgbYCVV3r5N+1cMSU/XIbZRVluPws+
AwvZI02RfEKLVoOGcKPIcQPbqeKnmVg3tZvl8f2YvDxUs3u0XoOhur66LU/i0e8eqV/AVuQrPK9q
xOQs0CBVuGARancnjFmVKjuy8TzvoPCzV6dcEgSWE4Fr/OFaBJO5umx1NJkGHdIhTAhXjRZOhhTl
3zdJ3LnKe2B2JwF4n4hrMrKPlX2FYb1m84wUSxz/KNLNx5gktoNW5oRt67ZIWBy+aCHLGKZw13IE
HfXgqCoCaUtgrVChq1MgukYhx0o7a6Ti9l3TuLKRRSKhcrzG2MgNvpRO4r6R7JL+DbxGlY7OE4Fr
UVwjH4qBhXuBCNBUnw0Vd5M8Ek+CYyqf9Mkfuz/VnvOu+3FPag63kMxKIpBBVdIl8eG0GKUPB2oa
e17Wi+d5m5fy3ELXTmoEb/VUcjsV126xefHd+spm6ZTPaynH2hql6i+tcjIjv8eZwVo99drZam0l
x8IfdBM+7Up4WRSDJ9kOP8FMyrmAH+ieKsEjYU5CI89v/xHQiafNRkM7bLTetn5ybEC9AffAeBrz
HhqoxAGlg/rzGV1rr3vBfMyQsL8H5KQK6EeJuS5e8v6ZBtbtBE7QDoqY3cqJeB/UrEJWtw5MI1iS
Lro6nGfO5YWo9uqNPTOZGKfoE5ywa7EzG5zt1w6eEdL+KlhAIdA3jNdHI9eO2S23anh9QHReZnPX
QtIWX5tCIqAXpr3xC2DuCylMOjVhBEyOUc2BEoSzT4Bayk8tAa7Xn1F5vAYyBb1yd5UQmw3jBXPY
H7wzL3CRIKCza5Iq6l03cFPa6UsBnhR7a4u2Z/R5Elp69OQVi3OCL46UKwFPeVMEyKOjygiDnw8K
REw4sbZanGjDH809u85kjGbiEpF/b/pgdeHTXCRaXNLfprZ3IghxrodZ8F67lI4s4hBY6gt84ewz
SfL+aktAIKAHepw+xoD5Ec13OzxOMMP2WWgqp5ZZ9qFKnKAsRbkDQ274IDaxF3urwiQ6oTbB89s2
ne5V1WLvbRIiuiPONSTTE9nPVd4IVDfm2A0uACmVQFUnDxA3S34/EZWvK+ekd169hJEBhLX08QME
7+mjoOo+h2JcUvwuNVyWX/XMgpqE8iY+BsUaVigIJTN1NRN4BSrM6KOGbsy96peGvKh7/6T+K3lS
I5FwCwuhZo42pKpt/GquwC5hDX6yzoUzNK99/v/dAdVZkcGaK7AfK1Ozd2JvAoougW7MGaF4DkOt
uKBig8zymD/zO2pfKR713MGz7mZ+qSKOsKIFvdFkziuJZeb983kxhkoG48uodvGDN8goE06dEK72
/kx1rnGo000bxXcZ3jjT1CIwDLTN+j954PQ7ZL/DASYYIlH9tCswwWbflaEP778CWiBI5ILMGF/b
3qqXy96/XTQDEDwE3mKT3CFGBZ5cCvRTSuPCNuhq0DFnBMkmxjPEzvHXUtBgdgzs01ejJ6ReyKzt
jgzC789yICRyoqMQakmW1joC1pK+ZtgMpTZXnY1AKOSgUj9nKluwDFIzRsYE+adOISWgOouq5yAg
KLT/Q+Y+2cwSDHKC1pSXt3e0G2cjjcq3AFC/dN0Tcp+/wjAqHS8qXRgYWRDARK0itNnupc/PdUjH
A+EftBbK/SVIOfhLmkG8NXIuBEHNCANa1zADI+Jdhz1V6o8z15TA9ZH19bV89aAPBAYKphsCM3AM
gGQZyAqYOTnwX4vpiQgKIse126XnmwbSWcxjnEZ4InEv4R5JBOTJteCxOPlQZCYPSIn8LsVVJy/c
eRrCoqtS3tJaFmdVR3GhBSX432zBBenB4eTSg8DYE3W81whey+XRK4U4YMvF8WJGbr7darMWJF6x
cCmwhLPkjm1ijuAcv6wiZHN4+yoXKgOWK6Fylr89pbtlKNtHwJbptiokdo/EvgV3ChF+cBQYIMgS
Yivvqt9PgB1PPUvxiMikgL/WrFQhGVWTyjerhUs+DYEd4Gao9uekzmQnRQ9NjcuwihFwmnW9pun+
GrzMkON7/nHx4XeXAR4+tpbd+0VCoF17/5qbeLt3wTymHtE2cGm7FTmtbU07pnWFpAZet1Bp7uI3
ZrVLAtL4rcCoRAdcF9RbMfQsHBKfcjPuHDcV/e/s+pW0u5VA5RD5Nkpb/xcYFc2dezr3bxWsmiCS
5X3tMbwFbk24WwS3b3piCTh0uLvB4kQSfnO1mJiLj+I3RsLPwbzZLOau+aC1MasIN+CcxSEy+ZxY
q0GTDZbrGxPFKP9ZfzU0lRUL+PI7rhzBg6iTQnwPI+Ox7nj5+tI3S4QYWIyvWuPYmtcsmSQehpg8
SGpUGeeStIev6uaTJYJCLi8Cw9xlZQwu6qFft+kELIklkCoYR35vzFVrucNKT3tt8n7qOhwY3PCI
lv/4J5KEKaaUaK7+Gjz2h6obeXWvA4RD+oog99b8fHhdd99C1CHBaNfTtOLTzyJXflsqu0vRq2xv
vVtje9/S2cmF/kZstorNfNxxqe7Dy7Tfz9yM8ecsRZK3lsXNnRJZKuZK2EKCBAEUcRWuYDlWqnwV
095dqciMW8if9W5b0ZHcD+yP9Z+aOVlsQiqv9T5TQoUgC5qKomRyaYYotG0os23/AlPuRifLz7+y
/dEI+VC80l1l39qa7dpAm4F239ZXdbWbwVpPZvMVNd025+aySg4WwlOXu8NErSClqH1egM7uNNFg
xXJkEKzTmSgZ7B1SUHEJvRIwZ5FZZLVqB12sasO0G2pLhiJa4LpmiwJ11WbMxhXRWIO+VcL1OmxZ
UJL1ryzYQ5yQaxyPHQNSiJY0B11J/gv9tu7gs0bat10snYuEAhwn1hXN0boLgwxdK+wvYFTozfcu
FqHkU866gG05bC4X0F/JzzeajxTcg5q+cLCMBSjrXa4pzPlUy+PyxHqfSUPyTDel0XkcKpNk0OUF
kbkgPGiyYV47UNR4gOg7nd7GDE0IioFEpiQ+SCi1OIrvoPBOnLUEHqjUF0I6n4hKXa4rZDM9M3Cf
4Cd3U8plG98EfWIjaMM8sdYjFXmE0ZNZ7UgTLPkJx2yNzZHnwNZ55MZY78S/lAiVLif5PAupGKmZ
gPy5hv4EwAPyMz2s+mF7oMXxK19Eqwb78f8pcwFsdeslTTb8c/ZvujBMUQg5GAmRMpPRxMPoBl0G
c2ozhvP5D9V8o3eYtEYSvzU7BH5M8WvlI+PDfKZZWEl+Xzou9oKZagzcm03a8ULKemUGnhV80wVY
W9PoEmIVX/M5BzJtfGjYvF+AxPOsdsZzRVcDjF7NI+DB3853yHt4vjTNgldG/ZqkqgqOSGo3kUn4
M58Q7YWTP+LpFBQ/BRPHYZSZ/0mqR67AtYmDqnjs5U3Gllg0+NCfqghA5df8scG+sKYGCavfvoNe
5eSBpoHOsj9xfLPM7/DMVitf4j7Gj9Nnm7Ff78OzeiV43AvSoq/Jjvzb95b3mhXjSAkUYuYPTl5a
KTWBsg8d9h9kviWhtijFbyYqai7LzXJLDnAywH+PQr3a1jq/mSzfyzbhwMJmXVR2a0AkkG/9HNMM
DDX9fB1pwsnc4ajHD/cuDZFDYEi0yAA2gWsUCxcF4osZMS0ZujKThZEMhMaqk5xyx/l7fIvrOVpo
k9iJYVyzPQbGVvf6T2e0vRnz49xqMGwvIsDNjszEY9Wap+LD+sEj53iPjXSTvp2In9zu5i77AzJV
Uxof62sFpeCD6m4mncrsaK4xcZnJC8LNFMQXP5KekJkpfiXV+kUcQvlSv4HDurxVs2BYSLtOQkwk
OG2A7tyefAwympw5EFqQbaXlUq7g/7QbLyFpdgnhABIzj2rNjUqIuA5YSd52QA+SNY8RoJ8b6JdA
zWzvYg5LE7RVbOWUtsU+zq8Tz9zh1vH866jEaJDuK3ZuLOhQlqzdKfmSrISnbX9oU+I9VY7BI3Ti
U6rU7eeDD0ppaMj93kUWP/6Ax7tXxS7+pTnhst/GFTh7DYLoln8gvuhldYb79AMDF2RdecngxtCR
GyTvJEn+000pnePPZew9bnjmQhy+xAS6AZpdJm8EiwK7rI8UqaempX8ysr8QYqmZeB5Ky5m22V8X
DcB+20Q4s75g/DNI/r8vaesnh9Lp9KCOR9eaOxePcpiXX70lKnkRpMagPw+kpXRzfFxXf7LJtSVx
0vrTVP+PiV3h4twnD0kfc7XuekAaDCHNjX+Mo+DmrqQAf0qXegRlpWx5hZ/22JcWzOja2TupQqUD
dcGgTPz/gr3hOESVLLUlqFghCYVXW47GXd/RHULnmaWpoq5//SsLpeuFRd/LzBbPxtUjqYTNm3p2
gvueUpzQBQYOxbvUH+W3eH2FAMTkXv15l//dVg2Eyg/gMuEnOusMR+SmP1yjO+9e4SYDCrtiHqur
00F4WvqHaMCLCcb+k8pnj++g2N+0e7q2w75UJx3Af7CfSvY6OJI+eBNlVYe2h3lZe6LDWkMYloiz
MKKClJo3o97RD1nghEJKTJ+NiZHLezwZueKUp2eKl+HJ9Ge0OOwBsuFizF0pP3qQ/krzoDwNJsvy
ucPzNV7/F1K0/TOL1uueQhQEhap2c6ZkAx5n/rcE02psvkO/Qy6FC5n5bcg3pcvXn+Q2xLnDRVhZ
0qt8VJHSjVboXrsy7LZoO4MRrStXXgOPRYyNmnIpt3Ejl6Kbcv18FMlkCdaNZfYAvM3kymKd4Qj0
F1fk0x2VjhC+031uFDksTcayoEwGces106Tg8b0K7Zme9ZtieSNLLFfKxxNqw9NsjgixnPCiP2xZ
ljG70X4dcmomkL2TTW3gWxz3u2SZgXAfe4tncuYeTgyIwG7Vj7XiwJ+M4f+VDOl89L4ppD0YXBzf
buZt6VrCTmgMM5AEeCLvpXeh9AfmPArvyEOfMHOAF9dy0vLNB5HyLEwdpTb9tw2tIGwCOXX7NlUO
l3mfjlWqqmSouSGbYRH2iTU3QjRb+Lo1xOAk2VgzrNVH08GPG0mbRNVrShu+Jfrcp5xgIpB715WM
jg2uax2CqrQZ5hFa37yZxcQyjLkPKDxhsKYQsL7MM7xOgJgoMK8xDZKIgCU/Dhk7P8oHFP2JaRSw
MeGRhjbXJ9aBnQFJBoMZTnf111GaWJ3hSz3EyhHsTpnlIrXqjNCeY4r2jbqZeS862BV/2PuuoxK0
rR2crgrEyoXH1h4rfUu5DtZOXrxRzokfaQLM8edti/wo539WyysOZHfCz8HG6u/a/NJknq2Bot88
4crWtuyJ+EoBp+OeO03lOv5s+gzmp1nnyoBuZKZxzEotDMF8LKj51PHTURP2BEQFXudK0viYU9RA
39enx8P3iRXxj3CergfelDZO2glnt3lUi2I10TEuhllgbbvsXBB7o9WPu0N66Nri0g+6jVBt2TB/
lxWZft0YOIZs4+oB49CuGNJZL/Baax+5jO6XMKyFWWETqnVypXbPnRqGKxU3B4tRuzyT3Mn/3AdY
dgAcs6mwr+L/fvur9s15J8785cLVbHKdBjmLrhiZk/MdcurnaxVv0/Ily8QoFhZYm841gPcR92ul
DVN+XtT3xO50PYRd4up8avV4Ix1CEf+sHsTmaiotRvzUOhsKR1X79+NDxz/M0HwveFLXjeaOFD6J
uvnZsRtzH6nxaZUXiux7qKkt5KB/5oPXNKsLnHBCTGRf5P5SaOK0Y/s5mNbwpxjgN03J7OqEOCdO
2sn/e2Ffg9ZgsUi7Q/dmMlkcZGfv9VqrOSOOlqVSN4zx6GPUSNUh8NjJRHDkJsjUmShZ27DLHqpn
Dryn8A55ur+UPWDHpPfvF5l+u/9Bz3L0gwjbgp1mYES3aoUAHNQOXsEWg6a1vdU/gY9WaRaZJIpI
d2HV/3RerY1GhM1Z8xXCCMk2Ba2SGkResXdp8TF4Cf42/qQDXbRMtoxYA/OlAiyiPEW0ce4fbOJw
aZYzrgWZvNGHq3y3xFCt7lhRmCluRte8iKVoGDCJnUSUZascsO1dZ2CS/UnPmdcKwI+3jOM/uwqP
5KdR+2uJox+Y8DrNTFj3+pQ9XPb2KYlGgIhS2H3hHkMKQWImmrWkL/wMgSDmNQyz0Rajn9mVS+Nv
+DH19r79Gr3GgFoYaqoUbBoV5DZn4NLxrtVt+Qs74imvBKQkrkpl3Mkb2ADDLCykBenC4LQ39D7D
OZWIxT4fihd+kjPzKlYtdRNI+DJFGlaBoUJwdz4rpmB5X0zOAZCerGGbC21TL/YgMHvG0KcbQke1
fHqHGSgSPyo8Bc96Tb79jZDuOxASQlymfcbhqcQyj5ud2eueDS565D0odC0raUXGu67LDOXiqn7P
XKmHS4slx/9KsABdvIXNngOM2hN+v/U13FwiSCR5X7fl2bgC/1gUElEZe3gVThlCy5qEeEslnBsU
aR12VPla9NIIS7DHs6VgyqkszPTXX7Zs1iBG87ZdL2P2PLrxD+fTICzGrioxD0dq4uHyvnGjXTCy
1dfvXMq6WIIErL3mK6N8+M0FH/tudsq2eN3ydPch8iU7pLZfaLyqWlWc+ggo2s5eoRgDkp8zT/mO
AMZnJFogZq55L8v6RmOuHK90Buzwr24ZPBN/Pmd6aIa4DEIiyai9BvHDVFPlY08fgYqv+eC5KP35
g9UFEvalERoLG7aju6ALDcJ8Mpu/jZBqsaJE7aRsEnZTr9ewk6n/V0jIaiBNGNNOB7mkLF9vyrXH
y7crFLV+D6tPW4FfdnkXvZ/ReakIAiA8x+5YjS62cz1+mR3Ka7ccimuMuAMUvrjaUi7JWMEBsWHO
jqLqIZfhgmq5L7UwAs2fFQVN368Ij5N7EluFhi652eF/wRN6a2TSL5D9pMfiaUFYIbmhDe/de/hX
l4HEKGXVlDwNY2oxbzQt1TfRiajJJLz3rEQLIUwrwrYpP7VFRas5x2Tk73/DiJyqPeOBhLkKMlop
hiQM/iD/5kzUxTFBX3tjiKyGPGrzK6USIeWqIOWsRodGBOfU+iH538hmB0y4ENG021SyWNRmj6in
3wxwc841p6SecxBgmKRZtS4du9YiRGxKQRwJ9Er46sRabsZ9fhvi+bRSXJozO21M0x5OyShYn/5t
oq999xjNVftGXt9i0ugiILutLq0F2Nu7F11vOP7dZRof0gdb+lE4u+inU07wBujTmHOoSfy7eeFp
qGhUHSsZll+jji+47gviOZ+rKh9VQeNRjWFnBKXk3jwCusQ+qCoHg2QCmslM6HSas9icfwAVLzRf
bfF8106LCH7XOTytUtezuFCXQU2SsdV/x+xGDzPxFPHseaoScMm1G3/Rr90jbvpuUv3GuQkbbwJ1
Q0ma1b3Ewq5kY63gWlgxw2pgmKxoE3mztJE6Z8ymrTdJSRma7VRv0ITYXkMO3ucs62pjMjjRCCqx
lE6OWMi5ytwq8jNJ3qxH+jrNtc8ltKWvflGXS/MuubrmvHZVZmAJX3DYnmIG93h1TM27XmVtZasL
e+1v3pX2DiwidAiEhDZZQcXJkGjt/2CEC5AiriYdR4cclIF/iArVVe8W9jIXy9dNHb7odrkcpS2N
+zz7mZJB779LRBaFwS6CzaOVicfPUQeGghpTp9IiJxFo+u/CmxeDLrOc9M5fcbhbqNhAZ0NsJ8xg
S1CJ0bDdQMVo6tU5ysMFsqas0fGMqZEQ1c70BO41FbVlzXoNxdq8rUem9DyHKIhVhe+9jNECK+QY
USNDF/VeKczXz3v5hzQNBLlXirB273Pm6fOp40EYVnRNst0QeX9LcYAPamgdqIftN6epFDiXgsEV
XwDk2HR6HDBzSrt94Dl/lI28pQ15Q3ywNBFjdDpzCQndQpShSBbyjok/zKMxG/JeYMsTmNdRhf4w
RVLRRGGTTV9SIVZQ8GpDamHck1UAXE1NPXR7WJ+Qbpej5os5wGUnO7tlWL0xpnpKEs2rMjordAXY
QeR+LXBfM+1w1AbwGfauutuegNmcuBkEIi7lAxVTM+i5rv9ATlTrOFr4OxsIJSQz3lpcWERpYSBH
A5aO0bVjnNY4GCV9c+TeDQEOWM6XvEqa4fiLHPVX1Tn/FD670JGCfKQ3pNpIeEVqZo/AD5YDruWt
y+2JSmROWHOSTPOn9DLNzqMJYEa6zqIthFCesgA93A4pfMA6F4KFmYTl3bxdsAho3lFWDv/VliF9
gs/5VvEKT6brNuilu3KT8pKQAU+C+AlM5Q1TI52ZcbbyQopFwXIxfwVdfu1PuFp22gKFDfwxX4oB
yQImRy2nC2aN5QXmJO9j0Zb4Nr9bh0WcrzrRSucXWkL9sFD4hC0GPuB8NH2hagnh47x/Ifcae3SW
14+jdbFypUW1xNHcgWJ1sjlNTQiE6JxWdJP7ORKW20L0F6b2IGHCGRxw5BnE/9AkPTeVCUC8QKUX
dBTZxp8eqxn38JaUnIBiIbV1k37+AxirTMoDWuSDDKLvX3fnhiGmpHVS8dJcFlClLQCgipHgcDlD
cC4wH04AoYprIIhTO3r6nFUi/JuckP6j5zSeGQloy+Byk5/T9czdJ1YevG44uD7hjnrtrGINJtV+
Dj+LYgrR1sjIta+4K7Hp28ndWjJ1+BTzQpc+bgEFXOg3ZXpanMjOMWHpLmCphduKsMS/jeSP5P3Y
uEGgefHHewj3Srrmi40X1mnuSsxvmJlzz2H7rUS5OIaY+RKuVVIMqkfDq0l2N5yEl5wvLjICLKwm
LPwWZjUWtqJZbp3N1ser4s5zFYX4nLZqCusuXD7k/PcWBoWR4ZRm/wYmXdb7Gy1VepkHKgVkXMM3
KsnY9YQNWJYclm42DyJ/xLkTSpowOUWWv6/WyeDeB/8ZnuCFugjdL16qzCc2WhznrwPtl9eGEM6c
ztQw8YfP0LajnWDg+HQNQH2IaEEXbpYBdWT3xZnXkc5SGTtoUiSf6ke1kk27xsn5EPVMmhmcpztE
bc8oXVozhjWgXXM0DvRrUzuMsZ10tZmEB9zOLppZdADRTOw9+OPDVAaHae1QwNLC3Zy2ZOKcny9M
WRz7VlcLDvUzV6+yYwSdX8+Iq5hS/iTfK/aATBRNJsR6+BeQNJ2WtVxItZfAoAxE88G+T+URShl1
gG8VSEsEGm7XhNJwO+JBMwcYCS7Yd6oxpo2HQCtNOIsXlRhqpG1KRGD6JDehJ155IGJL61SNiK5j
EF2BV5rQHBeWs2FuoGTZ9DvAzwhgBLXHVIxaIhBAnG0O/0dqXy7o3zX1AXJezhtAMPTz+ouHyfIP
KuNFOixdVm8hf9zU0v0eFD7LbFDauXRBx+cdTj+BG7PwYw4jctCdgAxslVwASYuLmCTqb3eflFce
KokGTldzhETJcniGsXq3tGPjRRUxBcuDldrhjJq5enX8ISsf8zAa28IGmO6ADijThURslSzWZHeh
4T64sAeIPG+HmowvAAiUOzymLlzsko62WqWmg/OkUOlTp/4dDc+e4LFNkKhawNaIfd4Fj4D3GevT
qJxnk9D4y9Ydi484aYOYDZn9bl5mGoRNR7oLw9fXMZOwvgYJejomEc//f24UDBqlqvmrV0iBrFjX
TyHUKEDyJF+XK5ixHcV8tSMTjtLQpRiL7Lm8edIXqP9D+XStwMK0UOQaW4YVyChVDJP4Innq3JBT
erFkZqZve/egGOT9hWQg5e2tDwcQ9ex82DrWLU2ciQOtyfAFaBqNEaYESHc7AiOPz5WTZcIrFeAg
0sAukAn/Lns96QAZU7urxCDTWQFatlIs5t/SFr0bIz3dB87MR9+AheDlcf04T4ux6xWubIG3fY0A
9eEK+ksSVW6W4YXgOv/EqKTAokvdqFgp3iYYwLl3zg6jaXTW5Hc3+njf38OitTq6vb6uTBUiaPFK
vBcvJHpJxN3B+ROOgSaRAllIskcDddqZx2xwMH5Nvk3x9Py+Abph+t7p0ozE3jL6xsH4m3rxW0Eu
dIYlAes5EYELnlbJM7+EFZRk8zZ+uLVfY0yPxaBjVTTpPN8sn3TLh9IHUemuaL+uVvb/JJneRSl3
9HL8LVuTOAUu+8wmusIJicndu/g3Rh9tv9fyShtSyJQWXGvfffqrjX3SzM3prpTqw3w9G5+CRehP
LEaq733eTwIZbIu4lLiqtefdYakWwwgAlEfESPRsDbIqZ4/OwKVjiIHoS7VdVG8UPZ6GeJFwTjG2
39OFDNWP2kaPjMTHD+oEF0qaUlqEHmOeYfAgLaJBOlASJ3EoXy/YOJLbkga47RBavQ8EoSDdtSQ1
bNUfcDe0GziR3+aaFEb4/tXB/+1NeoKUah4ICI5Gc31WSTV2leroLu3iT3HAgbhJC6k3iN93v2le
r5ruOZxRLtdvmiFGIoN8CMLSuKvR7G4+HtdzmuXfvvh38bky71ghiMHqPkExBAQ6OHPoBOmygQeu
o5t6attqo27HsIemqRYBy8GdXkAXeNHdscLRv8l9A9zOpGJ4eGeQaG160xJ4TgZVko4byH37QFb7
mqrkcIzo2va/jXcgZGBKHcu/1xCp530bBnG+3/FChr7EYSORSIzPheVwvNQTiVof/5qPUpvDH0Vu
OnAK4/ZGORKiCw9ns+gyrH8HE55J3Nl0rCB35LtML/9zuUYn/dpd1zDLnWyCRQ4dImaWWAMsuyJF
sGnCLZK9iH9MWCUP5fh2YUsCjyMkXOBZG5MF6pHoOlPbigfHRB6sZjoMMsQGbwV49+HEcNncSEA7
EW/4Z/VL/hBXbobbWJ1MfaUEft+NP4cvBQPGmADUG4pUCpjCcVuruwrQ316NVth2UvkZ9ata3Jva
4PsVeUNHDB3lEiEvACasEzGsyV/pwKQXV50Nz0FBCeHLjXxpuPLWqIgPVFFKEuCryjR4DsxtyHzc
de00iszQ3R495PqJh2tdhetWwN5L9PbnjfvZ/3hgCYwJG6pCob6mL6zPFqMKvmMWn/HpExi67NUx
I3+Bg2yitejN0YryOVXqzDGj3935lSRPNNNYHQ76Yvo0BgtRwODeTCM7j61LR+n4GQNSHMykXt9Z
MAe28GxX/MZFCuWzpLhirTbmNxs6RhHjqkF3qXmldEOEENw2AjmkX3jxk/D63zC8KI+mTzcaB+zB
r5lhOkqHwcNHD22jzIyHfCfHCIY9wb+MWlUB0l8yTivpL5O37Xwx+u4KMms8xh7ap4lQSlWLapYN
YprvBX5aopaq1sqg016qnTO5t/sY7dJqIKzGibBbc3ERANt5GIF7tEEoQ0U+y1UGzjZobZQgNJEy
X4lAqjoneXCkGzoNk4bM1jKlogbIpSn5+IoJAM3Q/2CNo45R4iJVjODuE7bACBqrIoCSzxNhk2xH
KQTv03KLKDehWWpnZgVoVEwlWkhA8+tNA24Wff5mvCku8GFysdeJnoyMO7lpiHeYfpxawrjCZaV6
toIvsEJ+ttllMfKRi+xBpv993Innv1Ol2YL1PqnrQ0ReflcGHLX3N2uVDZwJ6xdTjftBDlnwCwBn
g5aLiqY0gpj+8Ga3pkoP2NKtB0YMId0A4dYrTtvnPLV9gx2k24yaP9Fo0aN21UbI645xvjqPjuIJ
VIa5KI22GQHtZ2Hj1zL5FQjQxKicSKFeNvxhx8sVomXeV3ZWmGTwxtrOGVZK6PqxZ1bBL7RBZgKk
GSXVybjWFkbaMo/n+WVpGgq424Cy9Ajyw/EPIXQQdZvKs5mq4kbs2Mkm4Bw5I3n3IU1tjD+hyvMy
He15Wh6owMoySvRYkYBRMjVfJYboxColUZGS2yokEdXAg+hInKelMOA5KQseyXMfRrcifLXyP8vj
k5DEg/hucfyRYb82oaabkCJ6PLBg2ut46+OeksTf9rjMOQf1bTM0gA9hDtjwiiKJ3uVG1stcOrmM
gGxWj9pkDyL2ixTQ9PpCgX3tRHUyNbcap8t4KauFHL0B/2aIx56XcAF35r7q+KVoendicldzGYPk
PedAaMIFyiowGGx5qi/9AlrfYBquZZXxTTljOH6UKKlKQJV3YR92S4J8zHO6+bYiw2sT5+ytiivY
le7kazPxOcbrcTiEDFvTtmwX0yWbzZi8UyLhrYTUjYB9/ibVgmRcNsFbaHUs2iVuu+09saBHLIzV
9yHRIpmqAQuuiYaWqplZC3pYCCj+NW7pVSAfEKCSGcxJAq5ZUyRXz3R5txzZmulqDBx+s331L1Ii
JRh9aujOXYdSQzFsPbZQVxCr/atKKS5ikDMdxBeP9eU7msLmzHUsWZfi64Ui+XDUZ8RQR7CHoytq
fUC55LHDcBB9zVe1DBeyFKF4fJfMYzbdwz3Wvg68iy4mQTEg0ubWYru+IEDt9aJumb6YZwbAZy9x
gO8O3BqnOM0A01n4Yd+RyyNaDvx8z1i+EdB0RDn/rQjIUYwg+KPoGHjoo9uSTqUfhRDAWRwEiogo
23RgQ96qenR1tM0hryKMSULFkCbRDMghil5LIqT4sZm5eWmjfvHkXomeRI3I14QbT4254eYJGYUV
sAx2Z/QcpBW0MFBll1/bEnaN9vonFZcVtCUytfR0zADXDxBJ6abWx/g9vEpk1BtcxxK3iDBsbeVA
HqeRLAsCLc8xdi680gYDXbpxvbb2kz3yGpVNPsnb7RQL5awcLJkaAdcNEPASAPfo328sl2P34xIM
+GdKckzZsl2yNpOO4i8Qvgz4J5IU/hYVXAUTB85ZXbKjOv+Ld8VH9/6SVpbbSMSDvMu1eCqo2aE7
Z5hP5QXnvjy5ptDYU0nMIGLTlU+wQfA3lnSTucDhwV6VhU/ggf/xBR9YE7pUaS85Q0oRVshum4Lb
LR1OXyO7hZ1tqPQMd2gXFh2P/0VLlKRapoaYdYm/7vdnggDID8kddG2+49iVVMCjNUiS+LeSWHdm
wQ3VI7LzQn+bq/s2r2xTqu5rsuCzCtQPZQA6atMEKVTZd5KW+oXmnijaJepcIs1qyRteRymcSFB7
ypatfc1emjiUL3CBVhlWagACVm7OHZKpt+rE5l6+x1hGUkzRoct04fnd5rLL0VYe/miutpNDZocq
Wu6xxWsBhoIKL318eGBKxJMh7NMJR3OV9FfIh5GGYOHUUx0iAtFPkQCq98SdJ6YvX+pS3teQgSOf
RAMnEuAvKuHAvUWS62vIKGMy0ZPShHV8TK8jxQ+twvcIEP1Wejhp6Jft4H+yPL7N2X2g/Twuw0jm
T+tXXF1HjwaZIJWjPetMCRyO0UkQHS2JVoPJQFwqiN/7zadlvKvU5EZcRCgF6cFMh4VeNmse9vSD
EY6N1HoITCufwo5vXDKmZhu1w6xNnlyEuFgUifMdv601aVwB4IEsf9TynBC63Ibm8EJC6+X2dgg/
uMTY/mFPsS2wcq+06rC5D4VhPKGTe1mJ5RdBw3Zjnim62DoOK+++kWBM+9era78n92cwf23zeRB0
WONenhvZ2HNfOhHfwsFXxgf4gcx78TFLp/KBzsQAc9altQL2g3WbZZV6E4r4MIhTkARl3yVcwMLr
u2inWgx7VbplinINJKlqprTAXNcG6N5HG3H+k2rk7/eBRdQeza6wWL67PrwsBH5xTVtUNpbhXgCS
TzLjFn05RLu9hMndrWT4aG6y0WFBQPIMzLDJeEjh+nAP4T6A4zdGPRC9U3Hi1w0aPpRi8oVkvDgG
NnGNELb9cklNVDYxhKWGwXnkx0rQcdunu5SY1xtz27tSb1uNszflWQ6c040xcSeTZC7Pn7Tri7lG
z5ekcRs/8MNu7qxYtTPizpsVIkqEOJq/yT6TChyOe3QdpRZHLrXzqCEZvu8hFYP0eqzwlbRv9kkc
fcTcmA8wTeJ5G4QeHEueWtxzvAwlMpl1HGFgP2fKuAvXiFLDYUQnEc+69AP92//uyAQokX1TO6Qj
uU91Dzb2ZqL0nh2+iKDPdhGYjIlcNs0HDRl4Kz0a6E6MrW6WMVmHVbpBujxm4hMhmVX9zOm5tITq
whY2SWyA7e0br5ALllENm/P9InW4yyv418msaU1osP9z4y5zTvNlUnj/qbvyxn4iRwrHo+CKZWnz
vw69XFjqfuoytKWnWoCUJt6Cjw2FPPoR7B7N7269ng9Mq04pkaXBzt4577Zkhek/q9wA9EKvGkW3
40TN8g8PEzmS7GuKHixdBZWz80r2AEYLk+faK89Ad7rIU+/t9cMyv7n1LQCBygegnkAbWNZW0ZUX
AowJaVCovAdaEysyINOOgBZHSYewkon8fI7G+YBiWPGj+JFOeoW9U+HKB+fc9zyw40qm5HdBAQRd
5eKZFndQMZ6XV154S/wZ7mvoey9cVkSWdGBTD+BlasxjR5re5uLTP7GUyU49mQOwyZ6HnMlnpgBW
jegE5l/62WvHIbKvfEmkXTuhJW9u/a7KXr6hvBR3W8B9oXSo7DFKPEo3OGEOvNM4fAE9gp1NyT75
SPu1O8HpKkV4mEKaI8zlJJA96BIadHxgD+Tsg5H+zmAGvyN0f2TJD/azFmlcyAJCrCAAOttcAXBs
jRa7/lGMFCxCYUtSoCoBd75eAKa7k8F3X4E+x5ZLphfmaiJnc9lsjyS+8KE0VuyI7p36ihMxAF8t
3DFYzHH+YsMBNo2eQaAV0IQLvaV4Afm17Zckj2ZuGRTr4gftusVIckugBBWGZk9/idwfwtiaCRlp
abD2KzSGBOUE/+IF54+uRWvkkgwZqSb2nPula/mPDLve8624VZ8Ee3oQbXFE95rwSVwEAQYbrJ4A
fTPTjiXVUVSu083KTp6jtpLlgShenaN4vtgRisdxLh8uQBCxOmFhGgrunPMJTpziKrNnaZhdq0uo
kcLQx3/bWMCkjHbQTJzz82BFNusOgPauDz0xaySdvxpoQ51+Kcq3E+EDQ2a++gvIICnPTSKKh+7k
Pv6R2FqFY8fq/73/y6LQJ3WMCfZtuNilDdVh24MSAqHP2v5xlqR4tfS0OkUcfVNHoXsJcKbsBQ90
1D7WYzKzujk7xhYOLDltRTeF3WsXm0+gXtXdS5nvB3UGKBbuSulIzPri/AkTGKRxp/pf4Uyo1bGE
7y3pH9UqXl+77rKt339qASmwIIxSF9+EcotafmPtZQgbjGrz0CuQa303jHwDgv84caXmvLIKoMOW
dLIuS/YFsARhEdQ6aFaZxgickfg61UvbL0n1RMVZj3hnw1cmLkQhvaAOMmuqyMwdUS+M9P4MUoVW
USyfHE4WHPmD+RNw5rydWYrf4JFNLVdoRXAPdEv0oSHn4GLiJGFvogjIZjktLl2AAqSk5tL9tvG1
HUsuCW1aMYwdpz4dkCJLXJMAbnfhbospQsXl4yKPm7RP6VAaHM+idplMGmqOkpNIGcNsTU9bINPM
EFstVPtheTS5i/FbRCimykwUTG3EG2buAzCE3Z9JesL/atlfhJToGbWiL+02438zDeRpFdt4LzOu
6IzD15GtrlMq6XrTW4/PKtlpYy6xZJzNb/lO80yb10+wrVOpC7E5lgoS/yFSZo0tnC23im9mUqyi
LQsJPutK7PldtEg783ZlawOI+sKNLZfKoMbg8366DkvQg5ox+rF+8yZK+ZWxY5fhnDnF3a1A7tvF
Mi4Tp4xKnj/j+wYBmBxdY+H8LVfIwY0muiFTsBNoqYrEFf86y6TqXvwGYDsGST0oXUS3kJICCxyW
AY+E2dWJpriQTr+YGjwehF6npn6IYp2bP4MWMi0N527B8G+LE8H4kcr2zmfaofKIJUxw2HZEnEEO
49hN4NRLXJt8P7Dcp3gMpp7u9Ko8ssqmuVyzMZAma+Ow7SYzKQpy5EpPeoJAMbnCPV7Ht+Uqt8ci
aa4RHpKewQyu4vnKgPFsLq9g0DSF01TFI2/kpMj0DoPxpv6ScsDVNXHuTVq6kreSIGNihXmEIlQw
MvaIQ0IeaPbfsQOR3cF64aCzOigNDOmJWXsHrt1gqFWvkBSh9vyuHIeNyrUaQ+G6Yw1D5VX+0VuG
43H8ZI6Mk3+Fo/U4ELIvVJeFL5OzzOsNIbKNTzNGDcgtuxhrHKrUVVdiavq/MwJY8f7FIMGcD2c3
r3zN6pUOLdZGh6LJ4FtvOKvKkRDWY+uxa/2Yh/C9i8xc2Ut6W2Hx+0AXqhczPDqn4bno2MN+nli/
HLVISsE3Hih5qtsFdgo0XRQtQNFUu6sfWY5ZSMK6CG7J3YGMbiNqI2AaxDNKsmwXOpg4gcN7A9NJ
YppB5afdInU+BCkbjCoygmX5dkGnN/VVCqaaTpE0eYI+ClSrYyUxZUXTTtRJhZtlKGwlxssDlBKY
tpypfw2ur4qfYHMLPXmI0PWc88JfyV7ac4sIIVpbdAsZB6en6obPc4jDzN3cFkLc3uqNLQWQ2u7q
2uyIqUt3LWuoCj66kZsylHjc0qA9ccijaJWu3RL1V3Ejwod6bQhv7ohtuyzQCf4OAnc44XXMBxIz
4wWuaPDLoNdrZgPaeJ/2njzd+H26nGiaTes+EBB9XZp3q5JkCJ6TO3lbB62kE207ZziD6CUxX/az
6uv0OaP0ZYjLmZgsxEm0woGq96yHYzVRy/Yud7vplrm7NpWjvQ2HBHAw0QtIGoc+cqCmQeUmuxoX
RulwbeKhbmkKKlSo9hD4x5sLHVKoa66770SwqYDBmJ166icdIPN+G7KZKlUNThiyrYlLRiZa5e9G
bFpLtlHlBV7tRZefiiK3PTkrMc6Ou1Y72fL3HGrBsZrG5TvMUrGi64Jd/t4Ij06QpOHBIGpFrgHe
x18Vf2HaDMBv5mD4lAc5IfZ6u+5rNGex7D5JUltoFD59f/vQ6IgxXx1Bm5q7AfKycZISQP36h26z
AnxNOcW1ZhJEHE7uSSUClFHdjxZHpG5cm6+BFPdZZYz2PsXLPRc32CvCQLuHyX6Zs2aSs00Yf0P1
/khksptOyQDn/IR7oyw1Du0hXOn4tEYkQL1NwW3Ffn6k3d+FzyBoLGrBA8GavH2jawVwmHPUCBrp
5wHB9OexGIUMT37n1Ho1EuuUasoTW2L3B1MlF2MSB+056MP15pST7KZJtVQJzbtqRYMr+KLnsx5t
axLfWy83wEzRCo+1LFzhnmhWgt/kyxpnsUE3daPR+f0dpkr9xrqyExhqttXvWZ8FyLwfn6RT0ZEY
uCt116Op5soHM0jnCVvQQXllTGOb1C/lRe+QLi38/fk9xbbueG55OOMbTOYiQObjqnmrVLdV2BnS
98jV+vi1r4pL3BBtaGntVgC6ujYIC48mCie+0ptOqir00vqvI2BuEV7r1mph5GMMnzloccNLW4gG
ZmxWXj8waMy16bx/uYigTk5gScSG95LE5g33q6nGLyx8H1q73rQBstfELbDsfelAbeD3ZU6Y0ZmU
XfiipmprJ4PIZiepG1lwBTfpNCzRl1EF0ECTKG49oS+5xaHID10S6Sij88qszpD0meHCW/HDr+RZ
CfxrvTg0F3LkRGALzLBYWEF0d/iri66QASqjTA54DuGwHwFP6LLUy5kv1YGDu8mRCSA/79JJ271a
u0PlAG+ar3s2YQhN8mkXzvi88YqlLxENxLejwR8kAGfPqvhD8Lt8741rn5hrXSBnSC/aak40L5ib
jwXTzRExEQ4GKZ2O3eY1ZKSLjMwET0JY7ibvCR5ZFfITaQAJlWeZ0GLjzNp9kgqFLsGF4JQ4BgCS
XABJAnbNTutg8o6D+jQfI3+W/rEWv5OM8uYwHILigitc/GCepPJwmXtlT/M8D6szKh01uLeNHCZl
KCHqTD84R5eMlWr8cD6K3yAZsFxV7L7WpSNY2Z2Z3F4yNxyt+kjll2HbuiRarX0RfkNWotfFvSud
js43kFB4cghBn516hM1SiZuEXoctYgjY81HfGAEqd/iEbZ2XzQXfXOjQnUhK5rsDhF1Zm4GN3HjC
hdEJ59LzOQfp8z5X9wBlEDNlogjRcozvRszi+FZ94jIPdYh6EvSSuWTuXIWISbbWr8QEyRTVc+mQ
1/mS6Wi7Jfw7+xudkwcLRx23dXH375h715F6MImix02RQSxX+cdy7yt65rq8uSF5pT7E2PELrGHT
uqk8P9ATLSM8HzJznzOvPPqHc+7ALwrnEoFX/MvJ8clvp1Z0eRK50AlE8QeT6bqZmbAxPLbF9vhF
zu25Xe32gxGw2hX/bwC+E1JonUyGbZ6gnwEgziLduF19XA77aWK1PDWjj0IysEsxDCSHYHZQLOlR
3iqqOaoEEk8s/hGcp+oQKkofJJ3uVMssmiTPR8M8QsDLb2kFs8QOYyRKmbWaa4Yc/QH90hMUXIzB
0J++Wv3PNoqn/3w2IybO2+T5jnzDLLLoCzEX2TcRIdfVV8D4F8K5CYeXgfvm1VxlGkF1yvgtH77B
kOdPlyTroxA8KkvAOm60Z0UuGROPhMxSh42vTE5JXR2TvCMLVdfOIsbLM3HHXkB/t9iYXAMfMIy7
veVTWt+a3O5evLCdVNLfHnfUZfODk3Y6vrfSumStb5qvDMmc9uEx0LisbhBfUADL1puJGL0bzIOU
9W0B3pS0n6YsL/A245XMz9BTDD5+1E8Ok9myVVQKdkBJh+icypHIjQeLQ+PR0UXtNfP6wb6VAl6+
5mqk5Jid2ZcIbTLii7keS03Dcy55XoW9XoQrq8AQJN3ge23mDv/4j1Kk2A5EPqvb+/aiqpctcesD
5YHqNqHlmz7ESq1OS1GxJeQwcSgHlABfvSRyYrgXC1BeBh67OJEgEXLWFDxlz3lKJv8wwnHlRMW3
wKhTh43FPLO+wnl9L2+YB6CD5L49tV5ZEI9B+pDyAK3hYMRtSwt6B/yKFzjGVoX0OVQ93YWpz3fv
q/FLxHLVgHU1Lo2554ubfuTgbL6x2gVQph8VRubkssxSA4wmsHO5a26Prg1cRMZ1baRCS/bYToEA
3QrhM2zd+CsXNCnUUtkDn3aafG4qSEPRs8+6FwpAQB3XigMLBtnW9kQQKZO2TDQ00Sx8qC+bPfj+
EEAA0NPl+YTVUHD0Jfq345pIZ4o2Ll1VM8kstkX+RPULl26movujfqoaHup8M6fUsQEa0KCtBVxx
bQbHr6lTLcN+z3JmA30CsDSqakg4IaylhYSzCzssHPMeJxtA2Ltlb9fxlRIpD3RpCRUfYQhawXBT
pQ3jSwzYT2nmwDNWSjloeORa8ZqmfryJNyiIkGJQ6PeGvAafaDnfEIg3KBWpEoO4P5bIKf2kluaC
Fa2aguSco/GG3OeoOaLDgXXgjbHI09IAW49Zw1PtjHrMHrZCYkZ02x3R9I+mYUoNixXM+8IxfMa7
C0A+1bPTUCILldNDGfIOAVxh0bv2iFlW0Qak+V9hLfnjtVJh7vzlhn7RCfkUobTDk6WtVzIcOyJV
3T1ZsoqmE6tUtlusXTQG3z6Zp8wosPzvkk9leJXqS+N/5XJtpuSCd4Iz7UqGAIaYJ0oaPmzRjXdD
+qa1mcHrYLN4Op9ClBGQqZDt93VwYu4q3AyiYYtn8j0UJw6sr0wk1aw/e4XUBWrQPrmdDwUlagum
Gs83wjDS5uEP7zf6J6BqIjm69QIbpvk4CldP/aEf6g0XwyPu/e4z//6/jCXu4OZbsFZTHxhixPXH
aoA1ap0MKmgcnbS9/SQzNOl75mZx59D073D790yUIogNqxyUN8LlfPzmUb+sAxStg96RAO5ogHl9
rrzPJabFr4P9LBjCteE1S0bXUeBtsk5aCWR1oHzdue46OvtuEs9QWPQ4L4PRdJYdCGixjqasZU9B
j1eZSqa5JruCjmVHBzSf99zS7fBVALsEC+S0GFAIf9nintXF2cLVxAU4WP6VFLKRJ0/Z8IEv30or
1Si3XW1vJl7FpMWZxF7W2eanf78QyeYazJVqAYc9w4fAQ5sUPE8nWmaHex2ujGlxIJXheF+Rts1+
DJpPIp3sgNxrVw83lbjzhu/xnVSfvMD5tmot7ATWoXjR2HYIVJOAu47Q5hJwnkaJ+3nWXjeZeIP5
vMui9iSlXPKFUDn5N1HfXLyEbpFONuQYgDViSDg9hk/tlg/IfU0jR5XJMoMA6BloHFKt0DWZ4GUG
Q/f6Phnu9eZRssBPbsBA3Z/wUf0ppvdTCQUJdeTuvFfNHLcdM4VILSctPQSs85H8DZ+mfCvs7eMv
H5jJSAb+RrGAggwPq3Qi/tNsxR2X0OTW/10GYZjQFS5LZeCBIseQn5/YmD5RIaWPtkyNlvAwHhXj
FURPmavVonA4cwW9evNOHzr2TqawVCSKP0vRo5teQMR8rZhvXB8TxMqn8yHPkyPfKE8KDBV5LoQM
ijyy3obdGeiN6ehS7gaSvOVnL6/f2mrSPcIdpsByihpqi/4IoQLgN5wj1HwRyJN0nCkkx2G0aLDa
7fobx29u0NjFZ6uenYKnUCH9VWmkGsndw+r4hY13j2AJegShtabUUKEXu9Z8HEdG3AAmSSYEdVHC
heIFh+3KXOuRMT6d0pauqo7/7/Y6eYhaTmdNNA0wKpWt8FeW0rmj2JQbXQwF9HmaN6F3hjalMChb
xOVlIOxEiypJwnlGaldpJQqMgOpeguAdjSCH3xrmWekMBLS6exn+eASSvR9ve6xvp/n7smDbJvRQ
ShNywIVfT50PTl1VM2kRlbpKJ5mHKT6cUAuclCeo9JnDibrNMJkeWtON9JDsiYpTcJ4bsb1D9a59
r7QyRexvm3P3+2P2xbqZSqpE8GgvVBdzOtItlxzsbRAKpkmo97u4RS59UTuIMX1njgW/KU4OQiXq
P67LJuSrAjsx5qSkqWtvHxG8bOTh9WjB3epC6d61PPGVMgU7H6cDNL0A87ZPjil8tMaecK8xAge1
DywiWepqPOWUeecqi+5W9SHi+qDfQqoYfb5Rm+MPuPWhZwGSD4bqbuD1sQWuOUoXgCtV42Q1IwGd
CP+ZSwE1UarX+jSoofInJHkdMCFnjmXDF+Fqay8tLul5idcFucM7/GpF3o87P/MUS8QM+q1zTru+
vjgHvQUaYkRJ2XFr8WYhibEYh+8sF25BZWcH9SP7jAshK/hlArdN9NpGPuvCDrDCoJeRM7DxyF5G
enm33lWBpSYhbFpG5HoXtVkz7xrRxwb0UbYUk/rZ/UXX0WSHm/sEBZVwPg1crp2LIPI7XYy30CCx
5Yf/Z6q+yJBbZe/h571IgM7CUdDvfcI9zCub7n/4auK78B8WdNy4qYsLD9Y5tuGU4+7yr70ufBOe
t9hgJ4BxK/EvCwr61135FI3v3P2i5SD9ImNrRRc7PYBT0CXOY8OA6sAdcIPNX6sq6HFns4P34PRa
MQjZeJzDYMw4EHyLfkTkg+HshzJzVnx1OuYT2zE/G2W1kVQPDc1c9i4bn4MUGyyBlAtkysBdy1a6
+Gs54r/RTZYr+1HuKTNbxGP2pm4Z8aYG1gy+HGg8O1N4r2YedxRadxsicnHfT4nFn99aaBvgr8af
4HrsIuU4eb3CRQxr0zJNMOAX5W1W/RyzJd5YKBILg5u3MrrrOf8F8vAftP5wKrMFfketqWbLfodM
g4JAcETRJpvRzQknZl60FiTLblvSKKt/PcVQMt6UT/lZOH3ckszBaQnCKDFZhvkt+o4WM2TaR/n4
eASmpEnwR4V8qAorM7TsJap2LL5ecSsmuczYvabGwSBmaQ0hurKb8CL6BrdQhZ8X9rVyFeuYK6/B
jZjfc5Ci2PKEswRiw2oj/MUFW66G1Su2ixemAfjyQAy6mY9NIrHYpWjjgCAlXSbuTqRCLj/WaIGH
LzVYC2qx9mrrxt9UG8yzMpHzk3DGOLYL4dW7NIXGAQu/kmb5m/uVHLrnsh7rogNtoeBqalSULMrP
5bWEgpFUg/7PkP8h4mQONBM4/nieTu53Owkst+jF/tGDgiVI78bgJY04Byq8gesx+23IPkROiKMI
1fBKxpffnzWYoJce5ZrtNUzw9fYjhvPpK2wwu6ulkNOQw1xKu7HdUz/W+MqqaE9Ucu6QFICGcqNQ
+W/BUlFsja/Y7KCQbqPUtlVD+LxNxf8AWX1E++wfuxgGRFI+QrZCInLPx4tb96o7t3nUjTEMclq/
qpEqzu6iBn++I0ezwU0wOOzRm27a4Dyu5PT90/eVGFCqRKsiS3lsRmalFHQeIULzV2EljfumyHDI
Hi9qdTZfAcarnxB3PHVRTOmq8llVw8IvmmOmsSUz9eh5cp3Fz7mWKMg/Eeuj615YeYi3RCwLu97C
asyVjK6AQ+l93w4+T0pYmS7QICqQQOGmmzQ487WQo00NDgjPcMJogM6cgmqlAu4YQ2NrUHOzeWPO
MP0NNgR5TmulUD+uTnJC8/IhFXveQlDg8Cd/Y8isbVJaIqjkD748ktC+z3PtKg25YHVnm9PRNKW9
X6Q/hwIxKUQBal0LP+JJu/1XHl0Xz5+R2xIY5GMXhnvNcUgnfcdTFwuUJVJDIkb0cAuvh1B7CISE
0yeMSLsxcPXjpzGSjWo/wnLt1KJoZpmx70UJuAz0gkXKsk4zMaNYmWnm+AO99R0E+XSRJ/hHiyZW
M9P1hqbmMEVmBV2YHW2nAV10yLGbJ9QAv4ldltNwTQtgjuSQS9uDTHAZgf7cMtnDm5x5Pz7bJW8s
LQuGqctnfF79LS1eUJIuJ0Dcj58qLQeCh7DCkBGd1q3Q4cmIgK8QlDQGIKFj1BSa7oE849HiCpSq
QCp/j/941c6UpvnAMQUnzfwkRkXJZUwB3yeryiKFBZlWypVRRQmj2MIzHAkWbdF4mFfxoro5T5ld
ZLB8c6Xhuth/K6mcT892xRAXH1fDFCm38LnBw9qcUnSTnHM9Y3xjbgJhMHM2Jmpn7IKGPU4rb1Ra
5n1pfeIHKY68pL3xCNQrFyvSAIdDQrGdO6Yk35h2Fah+fzXHNu+VsYVKTLmdHjLEcJU0JmuiJFU/
lsQuN91AJmSFTNBIXO1+rnd4Jh3c+tyW6f3PTcrFcV69TVdNi1Vr/dYfyDJpB/+HMVqOQyNMXCal
zRRgBFNU37U+emvfm+oKSZdqim04f00fZ8QKtfsxvmIhrphmR2XKW3mvck20IEBzkvXF27cb73nK
t/mesP4u3jD6pkG7U79ixE4cCwrAHXl84LrcNcLfNK75AhMDzIHD1Cnv0NPdI9ZnLKWigtWq8kz7
yz9Wn3spVxBTxmNZqzgBs0YcXMbQ22kCBQ6N0NxQLBsJBvatR1R2eUNlJznNsvnbH6UwPc8Pxyjy
9AZo/T3yWe+XqafbMmRvItssnTFSjKxTCRn/WjhhJwnEgATG3NNm42iNcmZBZHqLS3LMuLIs7p+a
S+qMCn0com//454Exqwr0zLFkrd9+Sp5gXSxE/vT+FUYjDvKUEbbwY7t6SVX6CedVSM+2DQqHG7Q
GqnqTn2/NBryRaewxxbxp7X24XGZ3oJsE2ff+XM37o1TdD4npyvduEORZ6BovY/0ifjKrkWn7uzT
sHBVL0cwbAOuuwRe5Go7iOruhQ803GjTgoWOJPt8xFGQ+L2QBvKg8yNE66teK1p2R4ZZmfaq1AB8
4vgh5B3t6IbnhEhrd1zjaw+09IlXvizYExDsNoNdhwzw7ByimC43MTsLF8uXF1WZeXse+Z6PGrxs
tBGP7TAEs2wsWk93ojisi1Tepu1W6JzoeFpONHrANZy3TUk1+PmBgrBIawBkkHXJt03tLAWMlJXt
0/bKARgxwzI3MJ5sx3PZRVz5bTJLisOHUFxACGj4W651eu+We31WwV/iYRC3syaRBnlquiL8myu/
FPDXiSNNAsFONg59DhXqZRrltee0pDTE3/imaYI+NyRDMGgaBjpkxF9W7hejf9hyN7rDSLGIIOJU
Xeb9vc2UuqhKALKpg/f1q9iWpHE8CoAUSTPr0egVqv6Xt/UK+1nT25/PX1AsYkXEiZUjZvTTjzKU
SeHyS5LoOobGnW9c2/Excg7wSxzyz1cxz6J2QjFy2D1u+qYoiYRa/i8lCF/4TECWbSfsfECvgnkv
OiBu1X04Gv+q/DMota5IVL63neTWUXz2ryvEqzzG8hthXd9w1dkdyDvfPpxw81Okbj3yHQfhMfoi
hZMWSlrb+F1CoURL3m1Olywvef+53tnfIunn/myp4XlfZxvVPkbtKEMMg3xWmqIcr/5PluOmuf72
rJ81OUTQ5wRepu02d4b5ewP2Iu0FJvdKWjz3WLI75liB5jk+0+s+wSKCKANvtYnvzBqgZqA88glP
R6nVw3ys0AlLSvXKD/EB+xjE6F1ATmhbVTYkInjkls2Xn8Ys0p5FNTzTETKxqNKMhWTDYynPPtOr
E5pJRXSZykBU0mDeftUH+0c2mtyZXdHATA0SBN0sqtvhwlZs884pykTXU/Uu53OE32OZYMep3hJW
lwZjgFAlXPilpWjuHT88YTKjSvgaOHNhTIXkeK6pD4tWtGgmNxAhBZ2Qdft4/TP+4z2hOGn5Noom
4Rn3kiU3fWzFAtdxxZZsnufUWYDNMNCONk5iQVEaV4H2N9DbQuSxa9hC2hNdA0VCHotzhA8IKHio
cmsUBbL69UdIPekVH8f/LzRJXNqRrb5I/ZvxWpxWl1sRjpkohAGI3VHpHUxlHnEvdxOGK17/Nt3U
L7+s4U0fT9VgBuqVuRCJzsKmnRWdK7ftWm1tMFmivRzhgsFiiwcT4byu015BA4uviMvw9j59Oe6I
jRv21TOXCthdNbKVOILRvis6x6FL7IEnHkBfN7HFlEo0OzYkPzC/Zkcq1PAQ8ZjFya2xze8Gn0r2
79Fhn+e+QeoCU7VRFZa4dk16Sp+DScyNuSRXnoT74CYdyz++LFe7ICB6jdZuRa1/Rbb2u9+MIltl
qRvinM5R4AN7RlwXZKfYiMbS2EbznBUe6DgHHWqcwTi4ny4JiJYyfq4V6USsBKHLABydXqw85li+
8EbyIK5sFvTiyWDd9Wjws1Di77x+787vBSs5FLTlh5M0HSHKwHyK
`protect end_protected
