`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oykMm7p6mF/nrTigfK6qh/L/DUU87oWavl/K2s5V1Lde30If3DK2fHQKA2BUYpq7mrL6Q1N2BG1IfDGwmw4hzw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z3Cd+zRCMRTkTX85B1uzeNljfY87HpOdX+r2hdNnr62+U5Rv50JAgkNLrp9ll+G90uUSkzbyC3EFMFjYDetqD/Xtz+PJ+pAmGpdO9VBrBi3D/D1bY8WSX1cb1kan9tD7cHdEbFWCUIY3JS3IKWr3E23f3ZlJ/DhLIxvy9WGjEtQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BiHOlOv0uFIkZRBUMtYvQysEU6GKVLS3jcGNRBHez00jf3LLMw3NdoDVxaYTaxmI/4jtW0T7CA64nOAfbp4OPrzTin4mreLUci9ztHe7VeUnRdbi98ndomp9XPm9ofGl5vwASPpMjplErnrB8zguufLq1hskXknmKZeZYH+i9k1gd0eV88cQBKl8hfEqQoKa8AkfejlRq/rHCVN+s0QqtpM2/LxuE7m8BRgFXK2mVmh6W6tJChbb8gi1+ESKDP5ZvxBGrsAm5uSCKEGEqfIfoDU1L5L1Z8MTXMQMmwxbSPzFiS+5SGfmWlrLdzzh0OCOPA4db409Zw1dXeNsR2KIEw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nsyx+4cnP2Drj51ItDP4QEyTOrD3ujzGU7AGhTrpaQHFkglykmXP6SOcLVWDaaJ+/A2pHezjUhO1+pFyAy5sgZW+GMpXXsEvOOrgmKw13Q9JFF4vycqttBMsS2/JXidoAnvpF0gAaOiUhUvKs9W17igt8IkXoUmujBo+3wIGPXY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
r2EYdB3BWE1CzpCSlxxSWGptGsBuLM8GeYHpoVQf0WCz8zzttGg9XEJs6MZCa6X5GbMs9iYhcSlfkun1oVhHJPtfIdc3e9c7zV0xCdXlLaoUhUY44AASk1jEBU5ODRtDrTdRv1cdaBf5WLvFBQ6Gfzc+iCgZELBqG+DRXw+zTr8tj1VZD5VVvXy4BDPwtC3pBjV41wkhYWmURsOutZoYP4B88nWyCUt05pT85mNk/ai63TVyXsjRyDkl4rF/mHSL1gYDtjS+RLUJJsLGwdvTD2WzkrTswr167PqETWvoTFCMG4LIQWocLJtT90W556Qm/npDgrbcCvx4C7kyMgjBrg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5437)
`protect data_block
/J2blDtdWotPdCUl91MqR9QT6VYbIK+s5Mm+wL0U8LB8im0r8gvJ9l4qize6CP5Od02wK4s+Xwga
/41T10QHKd8n0ApS6o5OdW7dec53jqnvUH5sLbhj0TRXqfzCcmLe2dI0qoqjfMWwVcWYHi0epRVW
AmaTTeOB7DgzAtF9cjRUKjhvy67f8i/HPT4xWJ1QrmJ9dW2lFvXtwbwK1yLitbXNqsj6QdtLy8os
H2wxNUPWujs2diTbs5RkB1hQFhJQtr1vJBIs+g7qgHZdLPRpcYWzjBF3u05/XYKo2RqX4Bzq5834
gm1IneF/DEoiwmpIZV/3Tq8xv1Mq+o8EXBHzcgE4soAiIqkz4VsaPKSb+nBOqhYFmEznyK3c5XwL
YbDUpI12CgYaD58ATy3uBgkBYyijIKoccSRquj4iwk0VkLdKsPeHFEmcHNbY8QOJ1XtidQSzTFaI
iw3AQUQ81tndcgu55nqwch/dSHicwiMaxCqAUy3PHm53OZZZojNyVPrdrQ9ACjWghzcQH2/041du
xqewHsXDAn7ty4ZHimYrU5Y2jjxpyCi/JCkvsb0BHRCkrHJTGxeLcRKKLeeh1c6419iRo+GQufG5
9aRNCq8sodz+EVS1EK2VNUzr0jcV+NAsaV2nheIrVFa/xkC15bjYLNkh7OoQu5ir38WA4fYS6XgS
ztENC5E59qwwTS8/DiYgBD2gK75Yq7eIqPGj917yGVz0k1b2GPRHUp7iBq02JUp2B2rhyGxWhjWs
UBUFjMGu+kFj3T4WlrqROy2RuqUpofguUU0HFvSuJrfi6b3gcZzMsZzzDPGlISxQ3PT5SRSkCX4q
qQGftv43dRRILHu7/6EIWi00AbRR4ssjT3QAONO99mi2VR5BP6LrEK+i7yFPx+idJshTMFzolQyL
FWJPlGFlBKHN/H89aVR5gTbh31Lw1Bbp7mGE121arz1Zv15bDApr2DC8dIgQivbOjEZkAkpbxuIA
DX/JJNiwwCUhTgbPmBdVBuWZRbvMWo4MiajVfn6A1N+p4Kqj+9O1qrXpwJ04exqpiHnIHZ/qDrIt
vA59ROYknkWkz5KYxxBooZwq4wWVdMD6U3Z2amcwjcUtwnPJIQcw6ykXfmk1BnjrtImeiGcUDun8
zgtJLgsmfkBRKbKp9C1Wmpuw+7zFREm0QCt0svsWD9E2tZQX7r+cmU3Fufs113HmkP7MnxDk2vHJ
4JC9PR1SIBY6VILFYqJtaF9XsmXTdZHt9U1eQfYXEy3r/eBRNFDTty2O6D0ckM3SXZgSJQ1mTlNo
QLeZIiF4nZJBG5j++xZ0qcbgEq/HNMwA7OE+05QKmXW6ELS3P72nlMuv2LIBLB+aC0XDPvPcLYee
stOY05FW+R2xTkIxUGbC0AfdWkbJkRmQNnOOV+07jtMB27YuYW3Y0TfC4aoJe3fT6eFDS9ICCeFT
xPjh73WKaD2RMAZtOg7tXPt1t5gXV7Kef7Xj3sA70eM7tA2DXlpo1fHpNiIcGFaz+PYtCx1DBWp9
KABk7CVdtokvlkmbjmR5vQtRXLSBGEJu5ETe3BMDD6IXxLwkt9jEffYi5ni5+iW21ynzo/idy8ar
bM183LWWhqVOO8DJN+ChNcSZIRwM90SMhgG6PvS0XLSzl1UWSHiLWU8YhmdYhpVBlZbZs/0XWFoa
99KW3Rh+AZx2fPoa3OU3RQ7naoT4cMYU0AEaDP6vymOsTJkLeRGe8z8pA2NmFrvy0tOF27HwwRhc
Rz14zb6cYQ0LMxSTm+QmStIylrP9xiDCc1H2c34Ug/DsU2FCJI8sXSSApOlR3KcGdutkErMUfmAA
z7S+ZBiu61UhD3440U6oBMsAaL5wfjfhbFFNBAEPSD8HWvy1TEmVnpk/mGg84YZZ+FKl7bkvOyVO
3NiIbGMraD4OJgeI+d4E0UU5K5LeM/BhIToC4BQ7WXwDu8wD3TRHLtm8ezfwgMEAQThzskDbU3F6
O89kxP7hDe5Eho5Y1G6/tq/8eQuRdJVwRVLWEK/eMuV5VD3CbjipybMReNEW1thcsYjh45B/NiVR
48Yp4a0RVvyc2iPoymdAP5s7EmAztwjcRaE1Pv+aTsV5ZceMck0+yksVQHJOI3T4w/sDeGBZTRQw
ZLRuTn94+cWkxpVytvL2stpgbNYJUq2nktco1naYEul85bvBE7QyqpfO0v3Egrit132A42DSVjxY
6y8KUloe3l94vaeDUhEWgGLfZwJnazEZIbquhJqq0T06kTgcqnBa4CnHII3PnECMdBSkMmMilUfb
2ycfYv9U5U9fDJ2ed47/8nRTYCJf1ZP9Ivw6nPpZrtvgbZx1hnVJ2FvnvTv6tPg3n2iHBeM/vMUn
MWaq+VJdTo56gm3aMQZ1qbPMeL5Lf3vMhk0o8agtR7yWdmr94eGLbbhStOVHG0UJLvieWPwmgHfK
VPwbt35oKeeR5B88F2noo/LK1U+dTDmUr27OLEQGlgQtuF4/EB1krOsWLqbQF+yZWdy2q7zydcoa
bL2KxWCXAAvkVXHK8tqs96th5Il3Og4Bg+wd2LxZrwjGtK3To3CELPo7rr35PiggLk/LStn1e+84
SGfMuBSDiE5YHrkJVFklbjw/Myj83ujzxAf2l2HZuIOY4tHvuu3FWIxYv9nAB8Trxhe5+O0da/kv
JXXq3zomZfyli3GJZQEwB/wHe5pZoyek5GLCbr9Dnc0i057zuR6834qAdNDBUGHV5RFlXKKgNQkS
xImwDaOVrNa6yjh6a+YE0yRQhthp7uSAqxmU0cnQGt7PpLDJLGF3e/AxwLoJu5m88KNioSG/h70t
kgc+NmMvjJH9lYpHlvY/SB8cjZa/hpsbfBiStqPp1Mcy/AIp/4Y7Sr1epq3rchJetA2WQQGIyqaf
kyogExBul/ULzFPjtuqpyb3JTel7tqv6D9SqO56N6Z1RdQkLqvJjVF2/L7aEQKrrk38ZG+a3kj8g
B4vH3fw0ebrCJKjVMX7H85azpcDbHGlvon4p6nRk1FoCKDwJPPaJgFv0AWSk7PSHJ2MJaWesLqQd
9HG9fCxeCiqYRpUhTNiHDZ9cNNOskmuQzQ07ZxvfN00qKUExQX92pdAfLK9mQZrRKngSrsPvqrJx
eN+gcdhdaax5KG4Qy9pFPCUnh4LnNkfS99MSNhY/jEgD+DaAa5HrzCUAiDVV1u2mR4gtqGCdObqB
jOU97BDr8a4PduhIFOa6uP2KV+S1Vq+7W75xNVy6MhdFNfSBj//EAnKPYgd9GzImA8Q+axsejJYj
NioVws5LuWgBWL6j8C58QxN5RDxBTqDW1WGFhKmD2dCIrFEfmXMw3PgAO1GfVIAHOpts1PEiX1pe
b6ex3l/xUzccMzRKo3k9ksmUUzC5WlxkT7UFXzbWQ+55jixH4LJjL4pv2bx9wRrq2/s8mnaXmhBW
ZZBBEafBqDEn/bH3F0+26LZPoLPqEIEso7i/JIm052KKf6NwVvnc/qBdvu5N/YydNRhnyC3yapRT
wsNWmwr47bz8TLtk3fcHakWvceOZgJT2JIM9PvQEZy+l9TNF2fVC5CtxfMEmbrsRXaGmsHdkHXeu
pRDf2d//uQvNQVpx4iMMCukMJD8E3TBiYHZ44bG4mKe4OwH2BlD0lWh8zHynk3uEnguMcRnsHkqS
kHKjFhgRopkjnBi65PT5PNvS+IoYxmlTN/f6k3QdIzPcft8f+ov9ezvv+VnkXbX8wIYw12A+I2/H
4M8Bq5FbglLXcySDPs9vrdSqFc1npEO8I7wIemxwxSckMM3UC0EJuMbyM1bS/82BWCk1t7xzTcVS
bUhjnC//Ip9PvqrsCzsnVqoXUmtmF09PEnv0uKKo63djxL8wDS7qBhLj5RGAwTwwYdji8n+DXm0Z
VqKGBkpPb0eZ8bjGNHvoF6QZKhBQuXLHdT2AlzCO3noRaibfUuc5Yd0GuCDghXEkKSMFbFSfjX+c
mcZD1Aj9NtPuq5eY+nLpQ5IhysvbbItumNA0lBqT/EG1An9rsv7rpcwmRAGxq4AF+QKiyHGWIKak
DeEtD4CMWSjMgtWSRxEVckczu5Ffob3AUVzJ+BAxtTYGW9BAjvek0j+jB3i5hzngVdTcHFcKgjWV
A0GvCQbIrhcvfGcGU7Hrg1O8lWuBW2w03uSO8bpgVVPHlN8h9auIBjQxxUNSfAPUVsABoYOwAzHy
idZd3UbltbnXZiO9O214f+zHzJy75tYI6UWifHnf2pHdkBuhTz9W0Qarsn4806upTFOHGEl2yO0o
sPtaAwt0Hopy67j2y2v+nt2htX3wl7SM7f7NLlAa2w7ZNHiRf/o0pRF83ioCaWj7U9hGXILb6m16
Zi9a38UynWLIPbTiTJ8Pw+zvthGJ7xlwzUomCTm+/WlRmOTX+ryNETsFUXqGMyKIiKmU0kV0HUNV
IlgHU/gOMfuPj4x0js0+z99M83l42kAzjuRymVlQVcqenurav+153DUVzxVNUd3ErCqUiv68Y5JK
IldWW7LIR5Ox0sj6iBK7GrdVXcaMRDsc+QXTxAWdDTycElnzhz2AmYc1CNHocMw5Iq8/XVmFSOQ/
8binUlEP5iXVJMeo0EXTRXozEwaDnoGKIeLqyn1XHt4NWpDfeSpwqCS39q2RzTA4msAf6cV+XE6O
rGGGsxcD7fHkrSmDzMU7+j8ocYBgTloeNNusuYLOxh5itqOLfYUjE+Zym6/s1eH7c6nYpRJTUFip
bvlZQTt0WCmLSxpnxN0vCczeKIrvvg1F1yI7KDiAjuQ31vXil+aQr+EJ5Z7og/U/T4z0zMlc5o/a
VJMiHUPSKHnRV6CPN7NSVSTkly3v6TJuLbzyfw9zePu5tnrQrXXl6VQrx1fUYGi5ROjAgNiTN0en
ARrmd5r5B0Rzagi6DNJKqLDqVTrtyiCnlJ4ZilhxdqKCfkEiDub60H32IUopH7HkNiF7aYip5PMy
WtYKObuoU7niURXYQyARsIDNAWjuC2zBiOihtWxzHxDDHjXGfxMjhL2qzKHupxqdBsU0GM7EXrht
JgtPbux/1sKZWnmAOm1Y/xBYbrj+p6LIga7Q/Ra52bYnV7WUNJ9usXn6AkcsedhoUFccr8k0ur3y
nGcoi+4275GAIVqgO59jJQQo0UyOjVhk7IeIbVTrl78aN+zfeWIVLfdS3efubFKhlFpWTl/x21k/
FUrMgTlGozsA5pB4JDZbFwe7Xy4MeCe5wRXyWjBbcBQf40wARTD4c/nJR2+rD/zxJIU9Tsl1MiXm
182OLLWKcSkkTmCY7gM5zurbWCgnuSBqOi7A97lXiAOyZjej/Rb8KZYFSfAa2PhUU4TSaFLfZHtu
IqEdzrLsOjBd5aaGd1hWGDuJsJJotDXK8OfFLLlSuvYOk192CRXkW9oTsL3g8GdgZlVt5Jq/AEza
AZxz2oxl2kM/tAr3KHHkOwEB28VqAXhHgl2DC2RHYXSrg2m60FVzofzY0qTDSxYUkSA41t6urIaC
W2x7ZNF/4wDaQo+GX2AMa8oyfqRGN4+kSXJR+NkHhIHdh+IIVdg3aOObvvQm4h3s33c7Zg7Xr+Nl
gEPFFR4ELONglIdi3yEX2WhhJ664F8JJBWkKBPSDapyrtMzVVCTRTmcAFLDflkF1qd/b1hPEBnAy
NxgDfRnKxsFGijbIeFCM89S5YGTjVlZYn+bhXpHRQu2621a5yYpkngf5nJQDlNfHo5EheUuAg+GB
rfAd2T/PMGRdaUBfZDQ0SYMFvgGEXBjOy/ytwT+K6XymeaIhz1IL5c6wUxeC0Zl39GCcQY7ZKhs/
uyc4TFCbm0e41xmrm6/oE3WsXLkcWTwLtMJMz4orAgRqriUdyEIYdrMB5sTsFK+CxDxIBifCmwHj
bBvqD5KHdP0NDogXorNEu2xuahiyDXrHCTnPHqyybz+IejOd2kk1ZmMpEwHFf8J8vgAArTjEz9hw
5aJGApMbvT1GpwVFAQ7/uiodkwrmyCOHdaBhjYVMKWgdGzatlF90lU40NwFBYWWbSDub93Ezx8ZL
k4/zuNLoYKNbFNJP2YTl0CXMSkoVbd9drQb+L7iv1D4MuzGJiBAEmheR+F59guW3ehUUTPwA+DED
+TAQ5fwKpeHJd7H9myWNPFYr6IRwE986dOrZsVJZbe6heHuKo4vZ2E0kAci5M3Fl7S3LRIuYhVcB
Ctb01Rxe5kN7nwW3xUupm6Iu3adw4Toesm8iqvJN2nJzV5Fl3eFguJlkaZT6R2A9ID/cPklK7S+X
/AkcOQGeac8CdVS5dfM2hLcZIXcOkcLgtEpkwEcdtJoXotB+Vp6XFh8EXffZzm5UHe1qse7UjecC
OBCMsRDxmWRPA0Kmhsp6ZmNCDycj6QcjatogBZGMj9V2VU0oiRlWOXI926MnXZWiT79gwCbzS+XY
VnDmEftntn2+56ub0VgxnkUd3h1aI+jTcBC8uvKzdoS1rjV2vWsOy19RCKrUWe3lDlVKxaeSdH8u
XpjKEgSoB79+5HYgEJswVogYQg02SBh4yIfhnT/HpRWVYUrNk7k3jeHI/EWAKUOYsItsqNTKvlSK
8AkVogKeVjcjBJATJZE0FRhAR4TVAeAR0SKcN59TsvXs8+5MPV6YCmFcdRpT22UpNfM4n3dh/vHZ
l+Gc/CVzOhkRTPcVfaroq40m11O8dVlTa+lWGDZIA+HK1hG7PBupnY2SozDGih8dj8BBlcaHq2Rl
ygbzblzsDnJjzIL73gwtCJnzizvpy+bsEj7TTpJpXcUqFa/u6MhGQcFLOyNskpGgpTC9x9qGteA6
9JfBAaHeBRbz2FtjOGvfdsynFOmPybYwZxOhfcEtvT5mceCR9dPTopolMpr3a3fOrb6VXKeIOVmw
CtEO4lGvVV0ObDPKe+5UZam0KboLAWiyqWt2Gs/jxrQ0mClMGrQitP7TEo/37PrqfxuqhWpbB1/0
7fRPl2i7JifudqZU1AGb3zhIkTjM66jYALWoPiZ0lQIzPtE6EED9Bx/F9CDNtyg/HhTdWvjf4+HB
q82jYkYdunYf9gypax4bWRm+VXCgD40r9k91s7yh3kC9a+46WkW+yYjoCd0mv+koVfzPiTudseUz
adyodb4AuRBooN5M2rM/rx+DoF1Llnom8KoWb0fdXy/vhN5YV/u+Pts3U42hcfIndnUgWCI8Mwj8
VvxTMIqCQ0XmBo5+xyb1bJ03BD6XwZsjt42bzXH5Zi3KN30Q6bpxw5/B9bCOUH+oCzmOIl7Xl2hM
gToME1ulAcbYWwWw9Mc55u7Y7OZcOTptNX+7+Znn1sps4QdRk1ZJGgQ=
`protect end_protected
