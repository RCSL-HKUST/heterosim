`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
md44ugCP+VD2NplSIgassxTlTWCGg82IsBUrhVNl/8EIJvImbHmHQ0qFtlOrCwcOzB2y64+VNGugUBlTPGt4IA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WuXqiGk8fga3/Q3ROOKQup6YiWONF7n9XeWY4XM+D8/Ikf3rKnHXLb/SgBCF48tdnFRgeFw96o2vlyCtkfYNHCXEF3n2nnKEMNQdeZUGkE1FNVvnZzDQNkFiNmmmxqJljgcDxByJ8CZyGTAah0YA50BqN1mVjMuPCz56A8a1VPg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Eje2U5uelEWM99CtxLTuBSiYMrKrTjAnAd1QqliVexqym2jZ7qUTRflu2BGWrC5WRIlKzweswg3FGrcPMjI72JH292fWh50P5qC6EFpF2muX12GM5eRrj/wy5v938MYX/9YAiGP2VFCKgbym3pP9/5acyumJ7dCILP6/kscbv5KltVS1ErFfqVoW16fdXRX9tkVqS67xY2PO5kqboGQRmVA7AlHrW6oldiJgdT+vam4nD3YM6CuXv90Bda+1J+CWDORvfVV+h1zhDXbpmHTCNYXGzHvUftJiUy7YlelrXy2+9hgmeGAhBUL6EqpFJ17I28HVuxE144ghEIkBna7X6Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ThU5lp5I/jx/YdPhNdpxR5lXfBxCSshikVpQT63Zuw5hhaP7bUBO4m0VPpOYWcBhCeL216rJ3Ap0RyWH61su5haAgILpZzzZVCQEErxHtOqZYvr520t2Ny3xeM5OzVEAMaKz7N5HIGrQEpCdwOFwKJn7dlQxpUwSA6PbnSAj3p0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T+vgqaJitMZDaV8yufow18uHhdn5vIeZo1GvlzmtRSAUwgGqCtXwC81yh5DfBdrpJeA0BAWbhoLGscDJ/Du/Kw/AsvJiCQKbtO7i6f0/4/OjpVZSLZxRGZm3NmxEOXVIHUObsQOUP0RuNT2NmLGb4tplFLRTqEGSeKCEsIqaXLj6SihE7LG7Dvww000Cfl3NiobswXjmKzxc/FGUYovFiulDh3qTVMsajsE+zDDxO2nYtWlY+2xGGHdn6rG1xZNkpSlu9n5dm8+de/A+P3+qgHUiDlbIpi/CbO/hjRieYDdoxGub3BjILkpCTYSWreqwaDGMzQ8oCgX0B8EPz8TQyg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24837)
`protect data_block
ZWJvLFr92uwQjycidHfvFapmF32oi4XCERhW5yNW45P8bPjKLU8Etd6yXohMSK9Pe81LszIQGmaS
Bqvt8mYnjntrwt4lTSbd6sViB8VXaIJDtUActz/kylZgIacXmOtwDvMVxEqW6n3yyzl6rbzGYRrl
xNGAcG7A8lSeiQxdscN7ieMYNOqC9dBvq2vutj84m9bkxsQarcJMZ3z7hYzoaKwq37iK04iYEaXp
N3F3sUxYBvzYBpSxGXyMtzDlL6TN9c+MzmAtQkSvKTs+LaeX9hlrld1e2NBiCX17FBCpSilJEWAS
Nyrj0ggpZawmWqADEbG9k+21HLloNo9/HykhLpvndyfeLwCiYus048/nqJhkq3Ua+8IOEEf/Alyg
HIPGb8pcB/F51rUzy4ZTqnIUa7YRUxc3eHAQytj/Od4vUC3eFtIhhfat8NLBxTuSiAC61nlHXmMK
mkJfIu7ySEds+qTzcU+XqQef3zDdD/2R9xj5qI6fY7c76uUa3NH9xgvDeu7Ptqsrcc7RhdBugxlQ
pfhQ961D2BlfeNwijab5cFg2ZwpW99hYRazIzLzyJ76c9Eu//DXt5u2U2RMiJlcBBaPH1Ryt2YmJ
6K9Nqkkx1/hB2gS2j3AIXSg7BeoFTliIo9MMk6/HGhgh68MAIqZBaD++e3TkZglMAv0ROBdf5s1g
r+AfQPdFwp9Iwy04/sWigkH4pI9/kBkr0XU0fTbtaJ4j4EpgBofJsjdMnkW1rs+O/Ll/Uebeh3y3
ujYfSAaaLgBn+utySTsyWOtBfHgNXDrc2D/ARz7SYE2blSt3mNd/S/QMrm5QWLewNTaSiokHkI5Y
9f1o6ncKSi2oU5X9M587IYzQTCBw+2ARplfVh+CFXPnlYL4xXAlhxj4jrwQDLPWFn1fTPLAia55s
F1wT8SxPTT173d3JNOY05Ei87wEx3R1ilAYoAqfH6VZgE/uzBauLEbaNfcPUjMhv9Sr13nmnWRvf
zNpVmmZ9p041DzrKZ8jtgy2/JsLzI2BMK77YM1KpTUHv/yuseYPxw93l02sLOaAIP8JK7mYa9TNv
sgpTUQoqEYdTXv6nBgGtEaQSqAmvhVt+NP2RlYxFy/Pl1Uj4C0aSgWOjv4SMopjVd2twsz3XRYHE
ePeiGhO5+RQOZv2aJgIOpl5B82pRt3G+d/dDRrbAXC6q+WWyAN7H5zA0x8fKVGlk1xadpdx83U+3
a90CnanOz/Mqv0Q60kl5ydmWJzWnzZwv0PAZmMbFWnUNTwrI7YIv0yC3df/JpIxO8L1Db/QieB0k
kWpMbGV162Jr5WLXnnIlmn/0rOCIWkmQo8vHyQ4Mo7jnEfXlh1XQ9ghfYSZY52yISREh9GOA4wPB
N7CZAejL4OYF1lKDbVqXf8vwL9zGzoWL4oO0BDruIniGEMLIFf+FhH6mqu+kibMzscKgf48Hqqs9
hIaWCscbsMRctINmFLbsQPO7EWIlc6bXdR45Qwf4ZOKcnue14UHn/sQ4pV7E3DoN+qdz7yWswzlG
bB5yA8ueHNrEqFFOFx/3cUOdpNf1WaCiWx6Er/TPNYZXnAp34C8ui6TrxvN8d4HUpN34qr6b0GUG
EmDcjKeWOjy+VQNd1tae8WqwdI0vBKvLrGtHm+8KrS7aSDgOFe2NFXLwU/VrX9Yz5FiCJBAmQsN/
+x848zS+9q4SjDC9joZDj1N31PzkxjpBWfV86hW2SJv0fvPCosfcZeKTZEi72vvXo+WU1ling4pS
Mj9k1ZnFSeC3oDfclpD0oEMKFcs8zknyfK2Xxh068F9Jsa2femMHbNHwFHpkoHLXY4LcrFn9i72q
NkJMvs2xt0fhWmAgLLQzs6okS6EKZIApGv6zsVzZiq/cdKUBUwuBV+AEFZILpw1Mq0hWG5LzPC2t
OknsoD+3c5qJOShM9RtTioFZr+nVUxFKlYr6IF/gm5SYoVEfavkyyAT4Y/+z7dFAEoEDZZroOw+q
3GIi+mW5HfebbvWazH1QRncPLS75oEiwCqMv13Xh8FSz8WALq9b8ub52kXunWfQopK83J2X7oBxd
Ri3BaaFKdyrqVWslxwsjDU6DgD+C1/yBIWuHigDMOJFY91pnSFpqpI70O+teaeRh0JuLdc21ssHO
kwWraVSTB/DGY8lr8s0DNycXS6kebjMpqjZcvnsaS2vPq/AqYf390UsUBOMZudUsD76fN98HWHas
jA0R3MTb2w1MtO2/ZSCYVz6NJTS1Izv2UlkBx7ez1aZ22b2gvUf1vdahbOeRwg5j//M2HwWCDsjs
xE8urfhrGe1tynHt02MKfAuHKWjoGhy5V9VLd8kmekBsFNzKlFOjJJU61zXUwVg9j9QrHEOYmqIr
C7gn3uc1UjH27gAO+pzS+Ny7jrBxfYk64RbNO9G/YiqFBsmy0A0qE0+ODfAl0eEIGV6RVBHvjtEw
XOLrhcI1yVfTIUd5LRJt1zFqYmUj0FUWHcx/+LIGRcHoj5pKNfGOajrfovJvQK8RLFvlHUnQu7bX
N9OXcqGNrynQpHx6APVxxaP7y/YuT7CZANGbhfIdsshd71U6sO/Ygimn74SMFdbys1HHxF6DKFOQ
wqHDYO/Tk87FgZfmSvg87Y0qB7+RpTTrI4kBcCCaz6W1G/hPyNF6jp3zXbK/rc/GqqvZrx/zgIwh
vndyjd5peia9SDCwuErgbpviwDajg7M6qYJvkVGd2al6TE6Yvj8L4ri00ILFVYCQXPkzBdyDz8MK
NH7gvNCZ2xW7FhbqFkX3KKVs57Ss8N7Zhd03wmWfntJJuQR0hQQ5aDAuMsCSIrK3SNFOkGv4ZhYn
p+csD0lFmtx0/ba9aNiujX71sNWvjfbbmWNglcbMV7qbEnkTE8ZVsGbD0UispJ9oJt+BPl2VCKhU
qYsKkKctJUf0uqpul+K1PEHfXojNeQ1IaCtnyVGfTeXGNQSd31thTsbzkybEVbRQxWl6aKB8PdPz
SJMMe/drqa0wVWJzjpGh2LHxKwHOh51MY7349uJyMRLZeZXyMQNehBdhHvNT+7YX6bit8mMTcafS
gSSaSV/A9CnImvqpOVGv/LnqgIk1OefvsWlSvQrna9YInIicINXNtfLRiD4wIzN9pp7Was1Oscgb
pZWqyceMMH/o00oUAmfA7QOtp5GcMBI9IcaesWYZkd9s6h8JtembKs63tJgaPDxn3KxxEOnJcQm+
qZnqQvw9/Z4NvnizezxxFE5BNhJKok/TZWItvz/AYMYFvGUKXa7Rmoysr07ZkXSM3Ib/MEKsDl3U
gqXvN4Ssl2kgeR4APRI65KquFgGGi5RLaoXvMf7u+5I+W9Axqt3BgK9upH/iM9hWRqsyhdiAhSIn
3LSRk96QeTogXG0wGI1xJpDYSpmOrrrG92+5RV1Xn92uk51BjzoX7WTTs+z/K6kJE8W3FVw4qVIq
kpRbNhFYFFMGvi2zAG8asE5ibA85xftu34BZYb91E2ky9IN8406rhQ84sVxUt3gkmKXX2AKxVSy5
OEoin9YzjjnavPioc9iHZ3p8c3nz5Mkn/cwSVX4uUQ+TZ8Lan6pzxc46RmaIXLvA3Qj7v5sxkFke
h8xfLnJB7jiVB4VOP1IA5RjyhMKLixjeU/594+/V7vQtmJXu1HKR24uqf0W0hZiaWVQgNWMOswi/
ym4d8RpLtmq2swx5GZgppO8JZhTKnzhm+vT7ntV9Ft/6TA6V9Qr0Mqphe1TQ2vhbsUSmA1iPFXkk
jKoOreC0Zy0RybI9ccFYATVW/22qYkTj7Zq0cw1LhrsYrjLtssH9b3m+Bk5nvYxPWcpWood7IOsG
JCxOSIMnxcYGMEhfH/HPVwB2oVmoyte4tCtYWdQBOuAIHzkOvwlfGVWMmTi8bLeBN8bKY89x/KIU
V6mR/Oq1nRXTE3IkODnjCuqoZ89Kl+PDl9blBefy5ZqBpXA5xFISo5H75HcFHZg4lexulGeX9kNE
iFrgU3zFS0dvxaKfefVTMVULlZQN7etBoi7ra2hmd6FvEvUEXFOyppOjPBMU7MUeFvyQUVQpobyC
o/lr82B26vCc/2EtyUOZeKSxxMX67x72g0qL5fOsZvx+7qNSt2GppyRprP3JlxTquALxIROYjH2u
opgZEkGboXweCvlWQ4JqFair1+eF1pO4V3pB5Mpo//qX+POHiumD5syIX3sQdatOf+asTfDAEtXU
GU2N4BMM96d+YESd5rgGyaQ3iBSbpHlBf3rX3OoVYlGSd6r7ZcImo+TsfiI0vjEsgyzz7txNL2lO
suGhfv42TEFfktvur6g4ipWLbpZLXufc/VgPosb/Km/9ZvzYQgiJmak34kPVYP8FGe/Q3yO0FfT6
vzErh877urc9yDgiX3XhyMcb5YxyLkHDPna9etRg11G8SMPSmLCQ09yPHXq/m2yIRJC19Xz3Rf9O
9cV5+i6FsuDh++F/Juwxc12sWnoQxV+lab+7u8LEjm3BVEEQQOBEHC59T19fOvjukOG80Fv0L4P+
LOGozzxucaiiHgXFBdNic2hV086oULdWnMVsSnRz0A2AH91e88WtHBlAYWMexrbnznXGfOKC9Wya
7FGIPhg2ILW4EcsEONmSop31oLnEiAGcVsOE++1E621BfrlVhrA8Aqxo3odtf6ZOQCS7JcwqiM58
TE60fIpLXY2JVUzP+V1riuCsBtGV8y2Qb5XBjGQrk1ohp35sXFX5WTlJyu/oijvFCrq4zGjTdrl6
s+6VE0jocu6STGQLXclAaXoRPK+6B3WweU18iK9ueeFsKSCviomZzx4/HlvkRbomDjaLY0n/rT1u
6U2lwOgdP6Rvq/6nQJLHU9eP2GrpEd1ijCjzApBSS9cnUpohAUlvwfFXbFmBI1X2EIfZ3LSBJYo6
H1VMMbc1RGUrm/DFIEk19vQETVVi4fqSKffbTkaY5KSiBwr3KakyVCB3pEq/0uB/mPCmAQEtksgB
etblyXY8JF/4TiGRVac6QH2W9k3FbohtbUJlK6T0ba8ikYS5w6cYRqh6DyUN4B3iWTrUN2l0guxU
Dm1S3hb4BJczZwYwXCStotlNbgQy9I3Q9hmMqiuk+zajHxtzh1fXIHRmr2o/u+X99rPcdqJ/hK36
fnKPQanb9SAksHAGlf1l4ukL2il8tRuzvU+E0Gm555IyfC1JHgmH9qzTu2nmev75+D2ITF/XBXca
XQ9Pbt6KvgepvuLYD18ppxQTEd1lQdwyRKfF8A2B2K/jhKmqCYcu/H1/qjkTCAlM7MeM2WH1rVal
1OGo1aAS3XGVt7x13PNcxPJp82XVkA6S9C0WvI5DgR0BXj0aepRtGx/HMvBQASRdZvwuEz5wjpnw
HUGc5PeuGkeF6xnIlO4LnZWnRX3/arLWOvhBgP3vN5q59B1nnP0Cv1WN3EtKTtN30G9qhOzmlUG8
XiE2BSIH6Y8gBSFGwSy4zYnHaRNZweCOV7pV0/Fc2WBPIrPcHhHD/W/m9UbonCf+aoyu+1SRCXG8
yc6PoqDnXxfpcV0VbrY3/0JqJGAeEHhn17l5hlyZM3K9STovmN8KXyqEsh2VH9LqQKXD1FC+SapG
NYoj7jJxYcQFZDxF4dAuZ3dgnz57TeXOJx3GDnw585MFPdV0pvp/j/OGQUCANS5q5nb7ZpmB6H37
hWmn2izfJQRqCgLhlKBaDi5LD4SxU3Vo/k8ufVIAEMVIgMwJyB8xs8zZS6GlFzsX/NSCXmlYPmbD
cJmQn+Bm2VlQtZl/bNrRBTLrSZSOJdSH+IJk0VWaUC1renCGkKfNAxFUwBLiOVD5nyoVeYSIzTi7
jMgerTVhQHFgh0SsDCb/RIYQ3EChyRiiUbyakpYeyBNpxHLZ+8OpGjvt+nCgHuTvEeG/us+LByEO
QuGF7zPjMKDeQciMgsduh/ngpEMYifr/lrraiRiInTreorqtPwc/wUIZBLXhhWpjT/T2gbFReW3Z
5VthHP+jib8FdGAh2+s6E6sVk0Bdz5lzTfGZnMXPNANlW/Y4rTLTlU7Jn2+wLxrYc3ir9joQyXCO
nKmZIpUSXMiKACowoveH6NphuZFqAzegoL9xR1IQijLwMgoWfKgM9xoKcqrs7W/kpE1CwhmpEbrA
YrkYcHeIwVUDx5x2m3YJ8r5k2xjPGvg9MGxrwcyKJ0T2Q9cgfJ2BhDmENDs2ZexbB0qy3fQTDDJa
fd8i3FSc1y0yjDXkP/RykU9A7CtjenfdcWnIhxVcG5uS8sMfug3QDbQBx8eTy0hi14l/uYaDk5Hr
MMcPESabN/N1qRsrNFtF8bzCPuxOJYp88eaZDYBR3rUBKYSmgt5i9LxKyII0GqW6QsFS1XSSoc7T
sBB4VwHGUEPV1leOdJjiIv9gvgH7W/aueJvA9GKBs6MZZU+9fhvj4KJVL/S9i85i6P4kdPt9tE4F
SAkICYg3IMSpajlw61Np6S27Ahm7pldSgLVOZEBZquzrd/Jb790r+oG+8qIvvLiNKyxof+UB2hnL
fma2j9/4XQu5pdcD2tNJBY0QQY1wU8A7SLfTy1lpZiWS/BGpTwTkSHz2cJArhgvHoFf1nSP5T12s
WWU7tWHaP9Vz0z3oAjPgsvTkzxeYrJErhM7UuZGv1Z0GmZVsKk1yKm06ga35Sklzp/ESDv3fXDRN
1cXsjRh4uMUrTn3VtXtAv8u3EI8Xrna6jKw26pQJ3mPVfYM+IroRNfhA0Qu3ETkpbs6WAm7m7N/d
OCiJGYTSH53nG4G2g1atpfrXHoeZLCVDpPOUoe3tNO+dId3Ks6+CoP0EIcUkWF7UrFSOUZaHZKsH
PQwol6KjWIMCX0UkilDewAOZ0iOHrGl8PXmGsseiUz7+ZOopb5R4kU/ITNseHICYHpep3kFsRvJz
b1SiQjrT2sfipXtq9rmlz2pAZt/qBaIh6UppRJIJy0xfsmLP1FvJskPrm1KT6cFkSOK0dI8Pag/F
/E9LlvFkM+LahclfbBcQmuSOhUR51Qj0HdN7y0wUFTZHaxaKALv57yIfiYtxAAscxJRBo9+2qwPa
PdDbNZ39npsSyBPRR8MBd2In2fr3xNvKGbehfjyC1tHItAN/5eGoUrtygK2hXH81Ih6ypgzHTODf
8Fc+/6iACanPd/L8xkIw2iK9Y/F1czDgcaIBm6K9B/hcLa1qApNTQcoMaC5k8uC6qeevkGJLh5oW
YiOOsxLa4FzY5xJ3/NMlxGM5Jz5dswvKUvPNXrIJeBRd8CUPYx2KwzI4WAFT4W1vEVrqB2Kl8Cdv
4lCZqfymlkuur0XPWeiII1c3FrJGYYMmvnXUlLaef9u6TW7QBJeTCzMPGdvivRfUCUDm2gyXw7vr
8eLrxQip8f6x8XHAAqQun1SlFHezhoCCcVqsoe4Xr2F2hwMhM+NABsC9pBWUsD36v6LBgUqC3oSb
WBk2Lih1BkwIwADLQs7Um6FyJ8ZyL8Zp432P1dal/ZPlO+OtOm4mEC6NhUQp7YF3uMkyhFWaGmLU
K+e5B4WKxEEmDThtQwY4GxwVHnZWENF3JNBwcAJk04xCV83S2DTEOC0Kz2OONns88LSK3OeOnt1X
MdIOxFfGimiFO1gJERQqrYYR9Smb7kq8aDzQhynAWSipgkm8PVuT5tHFuoe8F4pWBSkTh5yqAKLz
QVlAW7ms6lMkHDeUZea3Bn/5SOmdYi52/oQbUdIu/rLg1rnCifOGJCE4L06m3oFifVf3CiKqeiOZ
5mGH7iiRDMOVgYXWgDa0r5HfJiINxlXsEoJeO5pkhk09H4Sw+rxQnDtNBHyVueXpqL1qxADrzpcY
ahV2f5NYNHuMrYuFwT+uuFxle8kw1BDWKzBqWKmfQ94hbE77lENMMNFbp7qSQh6ekHw2wTlC8FKL
SdAOLsqh8DqGhEP+xOQ8gTpxye+gMMRGrzfFrjKwvJ/CIdMwvphE5V5vsWB88Hgx6es/LpgjQe5s
5M6dZMD3DodgxCvcw2wMF+AuJ6WhSUqweIaYDetBicGcUyaC0uS3yIrDnFM1uIkEvSFREMLO2M0E
OJJZLyCQ9PbszcMkaldy5DTnInXNjcEdNOznh/Z1VgkCQMAURvaHLWMEyDlsdaK76O7jW33cuPLe
Dw0GlaYN9Ve0krTPGZXB2hVZqk6ehlPLlx+0oOivDWGp7Lo36im8tVbfE788jfNMUDouLmJ89ZHx
nEUNg+CzNZ769V+yFKYqNCT3QPEyh6pThbp7C8TVcv3QBbOHnrIJn0g3u5528tWvwA0ddxmJEJDE
iSepV0Jf3+hxaegNw8ABJIewAsuLu12mfnktYV5ygpEiEzz/z/1YGw77pk/vBoBpFNcL472kCg1c
sU6PxEpmRUifMv4GVagzuaO04o/yoA9sB2sKypLZ9Jd759oZHcIYOFoXND+K4Wq49GkFNa/kewY0
U3izEB96SKbgtzyM2Be8aYeiq1zQsH6hV+7qIqgFZRYEyLiMy7Sq76BXsXbeKB4IIA262DvBkw/e
J8AgYUzDzBOx/Rgw9ZMWW2zjJxgfiFTLD2SdAX3p1QKGET2EuKce91mGtlVXFl/lTNGafiI18lAv
da+qGHS5k8bG8VFKkWutYfpXddP1SFrumZOF1Aml0aOAfV80yakrtBUQmmsHTFY617NTBk1yJVHq
PjMjmuD65kiCnoztl2A14eeL+Cr0OgyxOikNHGfXDpcbBrvn0qWOYxPH+E10IEpWlnv72oGT3eFk
sJm+baPdrR+qyP2mNKyqz4MMg2rbJsdV3EDW8ERARsLWFRyfUum0f/By6/FEzO+Yc+DpWKrjTC9K
tEQIB3tI/EIZegRyVf6nIRK48Rp8Dai3AiQFfRdy3iDvpYtA3SncMcbn6+f0g4K8hmEN4g+WIiAp
eExip+ViOdws5LUs+Rg8J10TxVzj37XK0oq5NquK09Nty8/PuhHAjGgEVvGECUSNy1GVpT1UXYIb
revDglZHj4WNms2qTrXtUw7NoMBvKU6eW0zTxi7s7jts/mcJoJWWu2WEJNtC9dAZF5cm3dUGBu1v
6eWxLB3RJiUTszNK5YYMVALQRCN5BEpEar6/PvLoIWpvNjtasIvaiaEa6yyBaKLdEKvlfN1c8yGP
MbQgwllL8i7TCJhetEksC83dagWTxn71tee5jgPWymz7UlPo5MAWn9zckZOoX70wO+/aDiPEF6W3
x786JWfBWA8//i9WvV8muqq3SmbhF205woNZSab1jadC32qNwRHWb0UDjOc5SGPTxv94JVo1EzI5
2RM0KB01A6bnjaFGCZFOTOLLlDCPUQ0/8LT82zxefQTHUGT44IaG3iJYDtdHV3JUdWYq/E8JXjk7
XCIkCGbeDhBOsBBnROKOxCef4134BFSKPvEzXQ2mkvWKiXhGDiyA/8iCYEuchMn/QXrds/19eiWe
WvVsm7Q3QTxVgOsxILObTN0RUhL7ApYy08yUJxM0HGbkiLKBuccI6LiwxPn6sJoCcWkBBU2ZyqwS
MYIF4O9ZFuUW9DoAIAa66uaWz87kXQE8ovyBPzJv+6KLT+hi7Du4AJbMflvCl/eGwQM4aRiXT1bs
V6SIJrTFGm94CmyCj1RYX4Wjw5A2zPcQH8E/4IuJPePd9sbE6uWulpZfi88bFIZDtJK9afuC+Esj
4Jpx+AChAq8/U0yjwmS0JJTpm+qzmBUzicdbigCQ/e0hao43tZxmmublL09/pA5sH0hRGOoHFObY
xULLW3Ba1psOtbqZXR+GdriSfKOmW0u+wvW2NIxAAUqv5YHNyzqbcTh1LlDZ4XTHlWHg/hZ7XfRN
JOBXyC5fXMiySVN7fuv6UcoJbeB3yGS2fXqGcmZJZ8Xw9rc8co1otbf+58eqiy6duSehV2QTdL0n
CQvZWdK6zMvI88veSKxoSLjO7Xwq2UfTOWvIRK//aU0xhQW3MZFAY+OYN6Axw5QT288LQBR7DFiP
KhkSqkObx70H2W+2/RzsA+AbRc/JvFcxkR6Nec2Cv40ui7h/lbWPORgL7IuNhtzFuxOoJVGBdb+U
plwFiU4SxbSOC1ujzhZYWaG+ZaOC85DDHAo87G8+BcslKGyhuouTpQxW6O7F/687LLpadBITQnc0
+FhVdMK+nypJcDog7zRDO6SRfyEOPb00I40oQpnPjBlCW0lvBj4mj5OD4PZrIpG1oNhH8H/30LjW
VD6vVxD3ezqY9ufoitI7xlQsA8+Wb42Sxs9TC9tIcX9O4M91bCBtUhs60IGvlW7iyOKeIs/C51bK
hvPyLHVnI5V2/lrM7aMcUo9QMCiv+mxqF2yrM1ksJBLVqGekBp7of1U8+JKcybY2uCFLmOTxVfLD
vv5KFgN5e44XSCG2TEMy4zlj5Oq0GGDBmzo1vsFNI7Bltv9ocgVk6R6r2S2HOcfagglu4oYv15tD
g4gm6jQOv5+L2F+fSzbXFEEFuIwqi9xJ+JwciXt/y4ctD0Xa9CcjwU7i/mx/CDpTl6Iy1it3dTgy
G6ytN0q5J/OJn5jlSqZ7xfYMQNY1Z4g6rfkb53BAz2l0f+zpStPvDLdZXm1SDa9C/s6pLOEUeVy3
+y35du9zu3lHOhTdO6GCtJSgXdp0S4Qr6G+YJREehWPVlgtMwSSqAKzatWBpTyH5YzqmzQiwoyMK
ck+F0q2XBJ1vxW63lOqx7dbvK7A6+c5t3EyIg9THRu8IC9C2lzY8rQAjIA3WJNOQw8SS8GAwkoXF
L6/zMaLFF+QXDcQBIWiiWBeRpSGjronYgVvORnQjS0whFb7nMNdwFV2G150as2jkxxDoGjK+P5ae
fQPTF/ngyciE0mlYE0AJ4z6V9Q6+7lzrKulFwCln40BbroP835iac5vydqWTHVcs0y4wny+fny+8
GK8AuolJJuooE/pMKytkCgr0s4GswOFqKsUy0yNGvhVqYQkdjocfvPAOvBsIjxobB+6KJCEa/y+P
E475cFV1VqgM5+ddeI6gd6SWRhPVbaaYSuKiYMqU4QhRrcZBjBvhADuPxUM7sQgX8/AWXZ/poolu
mLu83l5cXKRdY6Yu8EPQyp3JBOE4NtYNuB3b/1Gq0gpdacb6K7zwST645W1LIavdVnFO98geLCow
q3CmL2GmVzm7/+81BQhxZJsYM4XWsk7xjQ9k93LYsMNSPtOmuiqHnpKKWdUJa+mXi0uaD2z0bBno
oqyRfCHXP32caw3Qd9BM2vmbLIvU2F9woQBKJIiEfUWhwpzzYGbtiH0C4dqfLtHhzdQ5vwV+rr6+
yxtTPocN1UQjefCdaSuodh725IlZsGLa/1FmSMql/nhbzeTyC0MxE7yNbOcjGcJpbcTw9dH6lr0u
/bigzP9TA/Y30BfaQEiGhRLLWE6vnndE8U9dJQKT02BexKgchbpo9z+kjAgBPO5kvMfBbqRo8VD5
7LIw4vRgqT0Nfds+jVJge1Pr/dCrY5g6mGNzoEorMlbI6XxrWxa2fgXQPE4uvAacI5AadBCNPTl0
BJHvk4A8aqxEtjHxGihSkcO/Rp4SM56kjXPk9Adh2ivwakCWsDNRaXovQyMyFw5IQvx8Y5w9toKi
lBDd4cyPRZHmNmx5H1kR8usV6cq5yH9rt662bx42hQV6C0hGdJYXr+7fnqyfy8g8LPm8efYRHhaw
RjCYDiAtNkirUI89k8FNfa6guGAp/73Q6tabZXDLa0d8VtTbMg5Tdu1DNB00MF2v1tBoHhONyssN
AV6p6t0SmQK3+P8NDNex/7AalxcaxGJgqsbsj1CUojtnXDPtaXSTbEYk8zx6G9P76tRCWCQahkqx
9KWcg72liWSlP4r2R2UP9ym2jB40HGUWlvHqqJeLCfifXhLQwChx9dPK7rU/aIQlHatEDp/7bj8u
WMBTF95tjdr2rCY5oTHTDEcc8qWyQ2W6rcGws7jv5xzBhkobhMGrZhB7oWimWmz1U2Zz0iQPGvkj
4nw/ZENLMgXgXO39n20CelZ88eqC1Ed+rKDD36usk4vXZu+ZNGjxMGruf/mw/Et4bW+w7BOaxk6Z
PJOOcUCkjpY0J1LbsjT5qouHddOdxVjCQuFzW/f14zlwSKkQmOoaRW+AaLi2/z0ySAEnTcKwV2le
wKwu/+C/tz76w79eorOypHpmT907C6THisn+QilohpJGTmYTCyOcHdJz98f8cquj1DKxddEcqOpr
vSWhdJsZXOhD8qYYuOqqMIIpW+aGijG1VimfrEqW9Uew7+d6gL+QyEQKQxjnlwcwwmpgNS3fIbza
3Grn3CGx0/pViYX0HazCYzLqNfwxufVgQ3Rrlp/en9+5l3hsYEM8huINyCOzj5DSDTYwBh6Dnbs1
cgvj616/0+b+Pem9Vfpt57CRMzdLBB7GHhtTJaXo0nXIWBuj8h9zfoi5I4H4btGeZtgMpqWJ2TXH
XLOlm5Ay/ALYHApDjpfS6gjY0asA4Ot6qpp3Gg4VXrserZJNqHquIm/Ob72QhcyTbaXnvpkli4B1
OB0MhLmCUVYmVXtw2l/35Z4elW9t6DH0yVWpy2jyN9pUgucUmlLPlFsSJ7yCt+HwQoe9SiMopHtF
Nu9P3Je0jA9m2iegXlxc/xLejZxnDTQVvtFNkKMu7wRyMmwJWdDy3+zwdtcdd2m+Xns+AYSCrLqI
T+4eoRW283RahAFqq4GyaTDBBD7fXU5X5A8LgrAxlvA3ckbYOsGKLhPc9sejWVGq22xektba9dhH
3QsDKkYkMRrjI+1YWKcT4SWH4LUeDY+8jNDhuQyiSfgH3R7jeu+QMZ/uwtpXoE7z57RoAyt3PWeF
URB5Cu4uP3FODxLqq0fB/0c5H/oRKhxlgCY2GQOTzwNW8G3jzatLNr4K2kUkrCdIT50DlZp8RedZ
PrIq2aR/vUkeAbH2YbwuqIQJBnxFAzV6V3MrMN79Mqmblf6XR+OUWHJjPXBYIhQfTY2fj1+z0BiK
n8kTe9PglkHz996/togQBaB+csJqK4I0lj3TyNojRcQLVU/jgJ0mkY6I78XYFigGXKblW5RTGCku
eKnJmqP/opIyCCXmb/FZO1iYRpz36ASlKBSzeuexTZtiaa5NDJMphMS9Eeqj9u34bVhrPv+ppywA
0ex/cMKTsoOjW4tA/4ErhXVNlVGvnbokvihqGmnL4oGiJ2ZY9zFGFYp0Go8x779y+n8AlA2lG+Vv
U79E0HjCMiNA9c410PhiXgXr2hBCCarFV+rOHUMqfT98xqjFkczZSjmRTuA2XxTgEjNrHNyt2uH8
dlASNtuuo+JFLcx48qW9Whz5EpRR+Erc5Qvva1TezE0wsYyB0qTJUwYxanGUmwP//3wk6eU7AEpw
w/ychGeANOXZKr+HQYLgZBFVfkJIm9FjcAfkiHP/Ui/Im2+LbMpw0ay5P8ygd75daz32SQdtsXuW
48I807b87QJVXlz7bFAi58+mm14NMAYaD/aX5G1NjMmyDCaEc5uOH+/IKI1UzI1/0JafjjlbR9te
NYLW2dnOftMH7SuND1jfIkNoNSiLe3VdyItRiZgjOuoD3OgZr8fsSj8JfJ8WHxHnWUXCn5b9w1Vk
oznXEUxnC6TIz8dy6CyzsuLFzQFP2tKZDrmobGOVgBhJ/YW+9QmiqEDnu5VFZmBV5xST3UVRM7Ry
iYVXUsF82OBwMjt2USvquAB4n+Lr1aMvdrO9QqYoNHUbdzk9STbAQIGgyakMUEaBSaPmxU9dvN4r
LVNuQqUwMKKqYM0BaWocWDpcSZ0I3X2bpSKkqN8ECc/lwey/WE7bFNnNpgxo2h97S9Wwpe17K7WP
WjxR2fD+QU1c7azIHPuuz7+NROl/m653NqkTGTzq3IvoYBGuBQQBHCGesXEZUc0SKENsnAU4NxTL
aRUryaPwPqwxOi9izsrRXkwleyOPcIDIYBG6O/oSEeKR6YwW/wZtL3ho3Fr4YKKxM/fVDdyxwRjs
1fwAh3+cvLJ8uXMFvgSnhgwr6KjK64WaeQympDeTKNk0+fUmp1Vb4SSnoZh9HuV2q6BrLVom29MW
naYjI6yzQhQm6Vqn/cHACSLP9O68NSNG2tnckempRM805zC7GV5d5wiwnv941IRBcaxAM77YH6I7
409mFWZ1+UkVhrl7us2/cAyb22OqNSa5+uzZbbTzFZwwPrDIs7ndwFCRY47Z8ixGnsG6rSVwhzDB
r4I6+AKUwrw1o258zz1YuLK8xdH1ZNLIZY2NRJw+LIjnGqcfCP0p9dmGV7Z0q6m2/OKbnoZx9Jl8
YPWCGvgVoXKYlENZioTxW04vqrbb8lbMZSqswBg/pRbJKZK0EVkJ0svowHdLuaAUdZJ0GyWE1Vke
rWpFluoFiTXiDvx8HxT+z88VvhyBNVUZOa4/ld1zvyhRfFOudfjP4AEp1XodrW+fA4m/unp5Z3he
DmYVuQ9h/qSyfBjfJVbI4IXIEuFa/s2Dvfg62rASYraKJCspCmIdurUBBnwUK0diFh8oNyzGNKnw
UTn+BGZmC9kkJpyHyS1MQjbFuM1XOM/6vHoyWRHp1QVJJHJ+oJvYN1Iil9LbnWYasMfrVAD/sclE
KjiqfD1cPBtH2b8oBh7XM+61sS3FhT9u63a6OCI45pFScWo/jTBwwnKjwG68bmmUX18772Rwwy1+
zQUQhxaaw/sKLM8DSrdt5LEI2n0hu8HCI2G+4ruxbCkECBqM2vefOerrqjKUxNQ/uJyP4Uvcpve/
0rpmzOzhlBI2UG+bhvVDHhHrk9aM3zPbgc+E54cn3yAJ/LMlnQsXlMnTazaXwcklQht2BcJg3Ly4
/jtP6ETjYu/WeEWwRbqbXsttR85N7dDIuFSCe4GRmtNCP63r5lUawoYRwAqYVJfZI2TBqt1A3+EI
4lTrMg78cgbe/f0e/e1wPXtjZdTxJwhnh4Pv4e7qrdJL+cByhCUuU/4t27Is9MJMBHyKY4tZIkPV
p0oseYz7c4+kbpjw5qiLBPUnpPrPd6ZrBSinrz0cludAoXEdcGYxtWv+LXfgbiih1cU68Q7MDjsF
VxLMGS7dzHMH0maOsxcxarL5+cdMRTLnCK9g5NkiiHNU+in/Z2zuejufVZBHJpJa0Rj2ygIPLr7z
n8T8HL7otDZZ/8wktXBUEfZybYMPyPt8UfbjPVjsDW68QRK298WTCZidSi5wQVMQH0DPZB3bFDqh
eJUa1NqlIn2FjPRXg2SmNMjiy89Fxg0yKqajO/PI9chleQ+qKyOI+WGGbO7Nyri4J/XF7HxDe64y
GhsrkpRF7pPuvTgKYOUSqnNvgEhLtA3aIPoNfzKfnrawufs5KvNw7nCgT+npVynymGryrPXvgNa9
HWW1SNpfpg99y3Xne4k5bU8bFd2By+00Otjs5z+smhqRyvGBBNUHX+Dr2S8RZg/enZ0iLThtLGHj
KYlBbdrRqZUHsC4kHJHWWT6Anil8Ig4v5F/EUqAFPg3E0xq5ATrzRhE+7QPUQJwvyGyJAKgV+Lfm
ka0qZkVRaMIJDzj66ayYPpDJR52RlxMFSoNt9wcw8393+YWDLSet9EvAc4d2n/fbtB5nBQ3ho21n
b7SO1pZUeWVVqmwMJ/ZIG9OkcrNKJIMCgijMnp4f1ej6Yn1laXwcT8xA1zlw/b+tQSC1zJAlPP4N
ZZp0Ne/dq3wX3DkCdDTgCGg6YRVpB/RM5hvsRDR2ZNRLMDbQvk4w85B0L6/GIgnReTC1npMe9l/I
Jy/ygWGDh9zid/jTR/AwvZ8oM0jSGFUxk5plZPgQe+i3V0hhyC0UwGJ0yOUchDWzTO3nLYkoCk2H
I9QuLKRfDOJZqByGKGXVHYqLnwDVNo6OefRL6oDRh/Gs54sl0sEHcKHI+Y5aJwhj6cCikkifFo5A
Ywtr4auDgfVqF74BiPe1tWJMmOeCzJMwxjGIff3nh+yt4oBuM1NiZutzvwenLtf8A06GWTZ/YoyZ
b7zfm8L2X1T08nMWYEI29vXGqhp9wAdH51oVyXLoopxogqSCpIrrX03XU6lyN70XfcN0+QTVd3Y8
0o9Caf1IXh6obX1ds7UP5M5yldpDc+X6NQgsoa5Raj755madUa6ZQuL0mpXyDyPQ7yTcAa1j4Oun
SNSqa3Uv7xsnFKGS+ZlbPUaiVRtCHcHtlVgUnvqzJ1zH/KS7427dJk0681EwK6PbvlEWXUh4XyUf
7gHbE8rB95lVFxhJg1XFuDiLS5HEd37S+bC8cBYgNQ+Lg/lPQLnoOfOLEG0VJSgwV8a1klN9+cYa
hi32y+6vLCiw3gyOS4pn2UcwdIeqpiquDsAsL/LzNzQDvAEp4iqtA2EvJgcTOhJACNZ20nNIS6xg
lH1Ub57s526zgTcYLFtGB3qolyztdyQ2nVK/8sShV22GMpt+Z8QQ04eb/Qf5IYinTfIM5yLA8kKw
97F4UA1FXRfGZhhL7E6AtzA5m3lNtTSk2Bp985MvmdPpiP2RqrKRAfZmmg3HxdUfkMKXbaGtQ4XN
SG8C1enHAxi/mtLWKQPsa7g/RXLZqRgIXfxUcP7/W0pJ1jjZeQiInveM/bMI+lwHIfT+thwcd+YQ
oDyNQK8oGIbbQxwtZQnBSW5qRY+nvyh5wbYzUPLTGUySqOZrL4XhYBpdxiT01dc4mRKaK6Dw45CU
P8PUzBr7+exD8FpljjAsLi4uQt0Q3X0LVDGJdV2r/bvQZozXy08Bh63r051HCe4wAKQwxc0a/BpS
iNXSeZQCx7yZ4HnMCj99z1ErPngP+npNxBPhHuE4lntRb2KjIZuvt4YASI9Cbxa+JEeJj1xHQm5L
ScOc+miL1PfjtUpaCxMhuKGPNMPZBXp9Y52oRHl6V3nT6tIYeAzkzGKTP3YV+xU0dCAmG2/L8/pf
2kouMZVLYW9QaIOyEj0469Wjooeo6E4bGRJPG2/p0yLzbAkCJAB+ZtPW/HRKbb404JMgx1hRk/Yv
aC1sJH98SgE10qhQDvoVccILnYOKN1X+Trt7xWW8xy4Kw3/XCm/Zhe902NNaGm/AKvkRmySGmg3p
lixg6naRRkyR47QQld2XcWV50PgokxIZhml02asQXJavePiK2k2H6oXPThnENSuREEserxuACKL6
cqf7KRNj7hP8NB50L8LDfnnoVgb+1auNK0giNZEikEgH5dpMbaPX+Nsv5El6vpdmzrv5eiiA9CUU
G+0awaMhw0vMwofrtAWPkqQwXVNSy1YDCPx60cBBV7lPXzaYxw+AweTKWNAtRtwPG101RNw//PNL
NOaKTsS/ztv/cwCNzt1EjGr9kB+zZ+fqlT6rP4OF5Xh3rgEvRNxbpXtRziVeY0ejz3dr1m+qE59X
TsnKzP8Jq+KFQNNDnTxHXrcBMalPYApnsZDlJlHUrrOG+3nNsbZFQSxa1MgTmqDBpNsvbAHT0cuH
x/qre+V6xmJZTFW8NqrRQcS/q2lw46CRk0v9w4QUfzge4pPVQiRrpgLS7DpCxvxTrY/hPga4bthk
QO+n9o3LwbinG49pbPqEQawv1jFA2Z9yY7jpSW+bqn8hEJXr4CFGOXhLTW1FXwS7g8ozZUaLh4Px
uEfGVgvgwlw+QNwviyycX5ji6FPiKbGZvPyQ5xBCRHo3mLjyAPN2eu8dfjF8qhQgWCvBuc4EZPoQ
vS+QLn0ixgrjYIFNF0kxJB4ZplHSlF9vfpoxgWxSen4SxxQRJFXfkDYKxyuEaA70Tnaobk8Oxv03
yfFrMTi2dhrWJF+tHD3RBgu8LToZUV5KqbUXhCbFMgmtwTyyfnIvKSSZig7NjnHzm6GA26Nmyho4
jEJFWD+u+Bn/3aRdd41GajQillisTHY+LD/Ag89HUR7TuQ3hfGfhwWvlmeCWTYGKh6s+xUlkHdf9
OC1pZuizmnEXiZEuBOQE2tD7fz59HZ01WYKPVkm1hoPEGBQ3aX/6oKDCvzWmHCUdctdUmYPGSoIR
O2TXyqyMkt9r7Gzbtj3S8LaJ99PS2aLyIywx5dCwajWNacgoZmHa5M7HAfXVen9bp+ttUbVpxTXn
/CmcKRCQNBjnuUJczhLkStMWXn6XTI1UbS13My6QcRAn+Ym/8xsWGLx0QxZ0FmKecXreJ3LA/GAh
15qWtE3/6921IdrJ8qxDK3ofZ7a4aE0RCDmbafCQ536qo/tHDoUNgZ1uzqZaGOO5i9T4v4Gl7RDz
bPHoRqq+xUWQoVo48UkQ4dZcfT4I/VlpNBjEOAnlMTMWP0zrn4vPg9gSGEtITDNl2IoRlCObnDsG
mBR1wGaFZQIwIKNz8Aa2z3/hLKbXWgR7nzyi5Eq1x9n/41khiXH3P7e+VWC8qrZDGE91GpYqwGHU
6krZsyW6BiS62Sm2LvpGmRaJlBkwL+oW4gVsWygOn1PjvwJSeURcGTYgGOAdOl2mM2vT+7OkGRfj
k2x/0n/miHpES7fVE1ufvmPUymwfg6t3KDKVwvosz9LSzGkG2AOFvH9ZPFwgjF2SlIJez8t2yxzQ
+UDlBfBVDzkn1rL5LvYX9boMj+GFkHZpDIfKC6Dlqze/t78Lvo9wtCFS8qQxnlKevePQ8Q1b3GV+
9Yjx7O2upu8BukqAJou0SzVGzU3QdqKcS1wy0PkDcnMhoM1u7JHv1Ra4FSt4thzhggF7/7OpeJYl
UeTBDEO/IWc0vd5mJl3ACwCifX+y+7FZSn7gT0h8SetzTHFYFGeF02mUzHduNkDl9BPQ4E6IVUQj
Bz53p6Vv1EreaR6quz5f0Dy1aXGCDvRxNdmbOY/wfIXFoNTEmhH7mLL869qwAJeOsrEBBQBP1h0J
a6cOXj7BFxLUYsHvxFndjygq0IApp/TaqlnloRGix+sfHtclKoBuoleDfmtvT8djR4jMG9/OwvGT
uCNO5TTZfMgYr9SWOUGPqdMOjOYN5SCytmieWPsmQdyLhBwQxCKNv0944fZAReLRx1EDeV5FILye
GAlDF52S2+itB01FCVlNE/Cp+n0D3WAAeD9ps8Rep4oB/lgAuRbikHhInt7eDSxrw5Tn2RGEhrS+
bEhQiL3y8llqcpx8ZWdcvc3yybk2F/xbNaqkpVert4hZpQSbLpPGzOqrdl+9gyrWTZiLMCDCBkxu
ToVWEYkHL9CuRDmAFtz/G2DMqbIIiDq8Ops21msvjydbbOu2Maeb5XXwnsd9FBKVk0pVPPIbC9TQ
OT323U3e3UP/QKhGagb+ovOqXXelKgcZjTe78oZ9mE235DWLFT3TPjng2bMTy+zMTcoEbxRDHdos
t92Gp0WWUJJ4LlTM65bCuIIkVLVoz4h1gFRowG/ovy3x2kIEmVJ85HLF9hDn36N53S7GbpQlJ5Kb
xxcXxjdRK9Z46oBR0llbta/fkLsQdwy2mqdUAMF6kQ7WYaUq+TIFJk9Pbl0AWkrex+DCXd0rnHDo
MXqR/sdSVgalG+RW3kB2uQ4HYlXK35MZ8uCy5le7dv0uqgPDd+Y7eNRFPnk6d/EZDCASu4LuyD7p
wiNnlGIjAtvp6ZiT7pA8B5MFPGwPi+yDyIc96yLY7LcJ9QiX/UdmcuJan1qd+DuXHnzvXB8cQlzS
4uIp0dTxDs3WHLXs8T4m7P+FBxVJvmwRzeYR+0iW3bzDRlqjSxL2YkhcEKWquaw8W6jaMBNrwXL4
kEmGWa6qA0Vjx+XzfT877b7d3NNXRc4qrr/0cyeAe3k2/cutetMa0cX2T/0iT/IJCbxcp/mycRew
o1xp+vBV8lrMZ/1yNUVso8GW8lIEFEkjJw1k7jntfl9Wl5Hcwr4Vmju8eCCGBD5ITUzInG/rDnTo
EqA5H6bjfRu5RiMRMAseG0LVzcm6cFcFLcPlnK/uZrzCbbupnfatP0aFmCQmqcDm6jkZPekYmfCu
fVW5n2/jag1XmOPpB0nv7sx+++O5/Irr2amvT33238xumkTrJf3POBEvMDLMUA0nw9/WcORYmOBr
js4ENQVEbqt9dtuOyyBLGpc16SQvGfrYkSU8uFiW9KIviwqiuBfWKH08kc4LnwDU4s2J0QWtTBLz
Ju7Lx3B170P+SNTmK50QrLLlHx8DAkZ/rjXltnD3Rt2GDsJVOzC3R3eTud/s1/Wrlk0iVzXaEFfc
vTU5+IL4Ixl2VI0nRp5ARnwm59KPBU3KEvUzCfwbuEKFAZgfKSFFONAeglP3p+sKTbDMZVPplzIN
V89tcEl/IWYjW+z0cqmZNMIoBq8VCbRgTZ6webq4pgZsotNz7ckL24w8Hq9ZW0yc8c1f0NBmHKW8
/tAYnlJ8bcLqTBP9E+4mDQUngW67NT3QGGkeNvHlrxO/LNnqGpOUjoJVMsD5/PT1Q556iVewt1tO
dx+K8cTfJHYMlCgdekn8piv7/Me5c9e6uqh/OGr4gDYflkF7ALvIASrPU7605jM5CBAmQdBa94fO
IR3QWaE2XxwTRwnVhMBNUgV9z1yeMev7AG+ZMPLsPD+C0NctJRvcWvl34XeCza2DBAPhzx2VGASP
IfE0jTezzATh5nKPZmFgBjyfoaSe5PfqNIKi/0zM9PKzS6SaUdMobfHGrdD2veKklHqRihWcZhl3
Q1pE9ygEMVUQIN/iBefIjl9YfWkgKBPKhYCymQBlbzX+zft8TTwN+bsrntSBoAHTF3pbtMsxUgyj
fgd48gXpX8N69B2wLJ4Bk+qVGAfznMl3ArKfuWrLL2nAnyOCVtFBICP4+f+1BzsykwgPYDcgIgIR
uqFyPZrOj5ww2DBv9Cbb4nCaoCEL/pMvJJXBYirMYgj5rlBYS80qjS+zYjc8xMRPReAKbw7QoU/x
7JfXLqoF2x7SqGg51Kq6MtBa27niot/gmxG+rUz3WPaHOozYcM2cQo+W1KeGZDgzdwD6gAR2a8mv
u0rMufqcXAizUwCPWR69mGP2d69pqm9r8zAfGtqfRC+4TrGL14HXa5njGG41EFprl3pFNIXUD1S1
oWI3PJPEQu35WtlL//JKdSQZlDNhXjnmCoKuobyUoKDveh2oSKgYKfQIT3rjVj9gptaKJmG324Wa
N7EoaHT27+cSEhNvVp5BZkUCw6nR4PepFVFLLEbpvzuYzYY2aJJB1ZgcAMbhpXO/8hrXGJ3ledSY
SQRvgbmvB4YzfQejLcj5TiQgyHshbG2KQVaNIHaMf15/dFbcrP30u4jgw5GDM2P/QjE2Wrk6PoC7
dgyqg8iw8i3DBr+flXYG1oWhS+SV3hBpBpu9QQKWHweSAPSjOBQ+0aytITYRMnqPX4tj6gx2V58h
r9gnXQJKgyzW2JqDRGyXhn1YzTd7PUI/MykAMhscBl8LYW7qFMOQgRfWcx8KAuQZNCnEe2J1Ot1W
ptXm2GPjciIVJTUDqITcpbsR+tHaN72E63xbDmNh49jH1TNPyzVI8sDTsFsPKvOGhZEllSa4LOiY
VWfeYjPZzZN8WiacgNUJn20clwx1oXakntP3kNCYzLlN1zG0za+fZ5IR1MZMmpLHiRWQ+vrWX5a3
YDPZZLraTEcwZHNTu24SN6QZMzWyguuzdPfUfDvH6BC1QdewJogEMu7jl0JKGeZ+DjTqKwV0COMj
3SAXd47YMX42BEkSfyc6T2INFQkAjkMzRbgaHgQYlXhVjVyAXzsgtVa0xHEQuBraQQFsNvYzMvAc
RuJlOlZfKaSuFk/57mgO+6nUuvTOkZ4Ve7+fkvBXT+hyKa3MP4pvfc7mS+TCr67sYy1rCIpW8wgE
x6VkQlHJ6xlaYbbo9IwE7xX8rB6/BUrX3Ay/7M4NXKo6l0GVz9w3LPs/19zmtkHycG7qG/UEjwNw
gNHpnsYnVpA1ZaFTtdFbzGM9chs9E9ACJSntvhzR6dW1gYjzuXU4HlyuFERfevtIHCQrm6/cDNrV
clY3QvpeuT8ScyGpbhCOKEpEvSDAq6tlsbFQQ3rk86sExLIuwh24tmZu15GWr+3GgS9FVM+CYNeT
yR7txrsWTOJXUNwvsU0NpW2wPFxPlgU8rP7RMNOm4U/T5CneZSUE3dCyvTIMwRDU8qJgJ+5tqMcJ
7LwoQtBHTpsBFD66gwr1ir9tSeKF6CPExIYPJIZexFdnrxRKTueENGvwkG3Ku1yXIKa5sQFWnmge
3CHN/PBk4dw+JKyOIuTMKZht1MkrxMfBalcewvznVdyApGpnHzHeKu3Gt4GmXub+9S7NEumCyvsX
kZvzIqV4wXZ2VOGumwAcjseZa7UfqcBdLfYi5v44k/9yArtx5hl0FMfXN76XG53NjCyrhJ5YdZCk
voI4mqXfGzz9mun5vvh3I2m4tubnKgXcquEwu+QUvDtxbu6leyhXNXdgr3SvV9p/z7bJhlXzaXRK
nG3VF9oAMOTYTAheBc0tX7LquT9GhiCq27PIQPnI/NPEDl1muFK5icWbfoGHoncvjsxlGtzpdHZl
b2J6Ga1GaKWwsVfdXlrjH+Ow9YhOEnqSpmuI+SdLKOfCiib04taEqXiaPlQE/QfFZw1wMWrKK6CU
wkIq23H+DRHZvGLaEZSAPXP4sklnBuA02tHkoCm/et4iuWsLQt308wySdUifoC1KIV3dIpmIYW8M
I765RcGfb/ZQilgh2j9S2SfLoAnyk6wB2ISbOHfGPOv5ktwOfRaEiYGGU9b8rj9PpDJ6xzEv/a81
H4FAUkhmZiudf5G/pDAy1aciifZNGx8VEmxGvcAJSmZ6uHfHKh7BwS/TcqHwZQojdaQIeTs3lacH
XEk15+qbGJbxKEFWoFJxdj5uMBNCRwhpbhjrnxutqEaxjwxjRjRbo+cUf+voSkSxSn87SPgZ7T8x
ue0ZZFn+lE5Bi+/ggCIr+oiJ4qj8lp4wOhQzQ8pr9ZfXP3lz9ofhboY2iuQK1ftPJdH3ZsHbDg0y
K89n0K0/e05P0aa0BXjJip6+EMYsMBQ9QJWY2cAxUULkdLHDKh24/JvzbwM2OfVzrd9BtvtZsxWk
tN1/2PZIvEKcc9JZMA6V4YlSk/4svdLj2NqwNHALZKgvAyvLtIA0juHVJobvhnAWSOWGyMH9vpTA
fldk8FDJYyXO9ZnXFpaMxphM338L7zHIn4I9AIPTsgX47NTHDBN2zTPfgVVyUzcfNMexkSKZVzq6
I4Fq4zJKSelPfbmML1lx2IF27YAZWXitPnAGtc3zjT4VIfgJOb4jeHliNRtZzCJwYGljJx9XRe9c
pJFxgqRGSoapCd3kl1776FFWAxXvqCW67CYbMhqUi0ciSVsqmT7IDQ6qYkMhT/MM551KmppnJ6ek
6LELnlyGdDjjzL9qZMjrRmgjW15zqBT1apZiZCOeLZIq2m23pehJb9z70JxLtairSNTA5V3VmliF
Dix2M4g6+lTgUyoj/AIbtp9hIIuOS54b4qCCcOLf7iu06T8Nt/ln3rcOQwGqtp9u8RjzjG9ClMm1
DEVMRottY0m3LqJkBgGG4L6X/IcQD4G4+t8huSOqdCUOYalNmAJAWAJeCJnTxY4bgiCVacSIGipa
JvBp+Oc2LZd2rvKa3T9uniLLubNtkD9LV+QEq9fL53OUmArFxs0/G4+M0a2T+XwTgp46NKaGmmri
IqPcaFBaFJtdttuxWI1frkCZjroskKzn53SOB+yR6tQ/w7ws+Od7oap4uqD8mJHYSxHlrS1Nqqsl
Tmp709yvwm8lupc+tpq2WgpGShSkRMkf4rXE8+ZYFXgOp+gRByREa4Zzhb91davs5UGNfF+LA7Vv
PS69LTJyulP/itZrosLr2mprz2Q5F2rHDWnT/k+TZb3smaMwptn12AqHpFIAEePOQ+BUFOZHHS0/
5AJXwsJAOjb5heXGX+gMCE1dU2Qta84xjlAA75XgP5IPomb+ZmyJ9xKG+At9PuRcVy2C1C23Ce8E
hAtOFMwfkL2hiExFz07FFfjbqelpkJziNxB84OszyACy1DNUYLCy/L/ZvUK9s8CbjplZaOiaFQbx
i3SttzoY+aj4WZHVrsaQ++kcjpTG0iJ2gVWsSl+2819TY7DrbV2OrKDd+/nVwuwNajaozP5Ei9AI
CNh3X/3IRViill5WlnL9su89wTEUJEUMdCWLaD3QXF9T9EYnE5zteDUQbA1zPySZL6THK6k1ugMr
uof/flpir2tmR1jerKjfDCx3hKK/7Orf9izUxjzrjX9UAjAgxnKCSu22Kht6guNcAlvHWA1n/2nq
5KTI3xvRDgT9ZjLMIDAecnOPQ0BLc1TPvlrN2nzhyG6kCUdSWXZMz4JiUWdEkYLWrMdUKF0yuo5s
A84JBrucJHKQwkRA29s169C462Eht943oQulAJhVEYGAmh47H1kikWd0mPTBcpJ5qhSM0ET3Pde+
DPm5mioMuqjlGIKhXgmk+mzf+VaDIpj9zqTQ4C6cLVoY6OxooY1xM3FruUp2QWn0Fj6epdaB85xN
bwTUsIvG3z/kpF8XZDVMKW5uJHdHpxsZEt6MPDaMXuxzOtgDvmx/+ceRqv3YmP+yx2cxWw87K1sx
/QUcqd/QIJXGMao7qygRm2UvS37KewnzcdrRkcd/Tr1e4Ekh5JJi7sFGMRET0qj6HllojumwrZAU
D1Ai1CTNhttrQog0jg811NVNZKPCtB6xywAIZygrRiboNX9ngyiw2NY8knO3T929kzd1WNQPPOGt
jEeiUozC0+a2cQeN1eELzgG2gmGuuVSk1wkbVNeJ+/ZpkgfZLrurRrSHmChAa5QqqO5+Fa1aq3JP
5vPd0h7JEDteSlO0QlJV6kk3eVHhho+E1WMVUzZI8zoTMV0xXkzyEYeRcS4DbzIkyBilIq/D0tce
bl/+QL6DxGOzUwzgRwWtg329AW+Wp4bu2Me4LGx3Xqy4yRMHQVs2W0vtU5NsMWjFRYwb451x2h7V
BAi/lO6WAzsFaMnXExLWkfQa2N88bABpgBP3X3fGLWHpFJdFu4fvA3CNMe6cwCMzMnQodLBA1gfj
7FWe/tPtpDv2uIvZDMxcg1l31i53Q0lpiAPTTWDzKmCCAwLCBP94silYl5cJqq0k1x3ZPP+9LGo6
OTf9mJL/uesC/aHbpkOBzFb8hsATXppr2UzwLHJHtgd8DYCC/yYHPah8ae3YEEZAU/HJzo52ohCV
U3VamnLo6mrIFBubMCBuDyBOiVirAbESrNfCVgRp5zJPLSCJji8jX/EciJ2fFbY/5sz7LBvgNlFr
QFYwCSihQJTNFUJFm1DgIPSJnddnUrA7hucpohiBUusDDshk+VkPnCmPk2Okdtay6+CKchwesNHU
UJyHdKiZgGMjs2cyACQEqtyU/HhgPO1SKx8I4meEgK2TifoZTXQApwih/yfRu8fq/iDOhDx90qK3
EKZalGTDzsDZmhsPD4Hvg4k/J8iTCZpjIpBjvv3wXl+k7sbzjjmfpB0IUGaf41xrVgxbqM7THNnK
deuW7iGbhDoS7+bUmhYIRjMG2pFVvsHHuT50VsOJUteo8OdY4xWwhVmCHRliiJ2sCOsHQKVjSexa
3meQSVwzPaQVypEf3vom5Y+YqI57J3FeWcCMRhYTBU9m4RnMXEzlmUmynKBPBOnNNcv2mJ/oxi/H
8xW4Tlrza1C2d6A1aZaGYZYUc5/Uc5WDwNmylEEG7R5MEJTW25d8kyo18ekZJMcWpfkC7hZ9qlZB
4eBII19ezwLj2+pEw0xlGnj7sqY3M0Hw3ljUZzSe3Z6z90HcKFC4UYFTcDeucamfwx5JrhjNx6kC
RQuWz/zNipQRMO+LFCSE5EtQgG8Xye0M8ksg6+jTIBzjPoWPIryIf+2HNndhEdfKPAszNYNXAps0
EXFsnDjbq6dpNgWyad+ZlqfEfcOiw2KwHv0l5y7Xrm+rmovqWv4X+BxT/jR4Sknxa/8EykH2ou00
HmL9k/uVYdlkHPHAB4JYcNmhZxMJhgasbHYgEB92Z+bkWGVEdDCvLxPKG1SRg7yJhibnJDcyatpo
TJTEvAVFkio07OjN7td3/wsucAO/VgbUSqcwhsYqhE/KFq3vCY/vM2y5FykyJ6A4baOtnTSF5643
8FI504Ft1fW47MnieCQskkfN4uVLh2idpMSB09TmnbUAk3mFJrg089eTtc2qBiwX6bTGWXlGzSm4
vyzQ/7xJyLP8fdNdw8gM80p2drsVX1MP6HJjlU6eUxqjFB2TjIu5kOahP7y1IqHOogmtlO5imwbL
Y73/8OLAIYEqMuyVEpSfZ8vF8koFsl1b2fq9OZt7HGFMBp9r7TUNCnW6w5vS/D7nSwoszDyT7b/p
M7SPoQhtKgaI33wRFfpLRhn4zStKEcEFKr4Cj2uTVUHuGxKE7QKVQJjJ9pnsvw9w/sjoGwMxAyxs
IF/VFC8sQuDYCm9aumtlxjmkv86xoTWHIcfRJzdMRwTBKOdMBS57KkOUBL0RNGbmvtuawUsf3tEm
NBw14mv27XyXvaNKp8xJy7fLoY4Zi6Ct+FG4rbwf6CLlGM5mxkOGmZ9ZHpYSTwUK7Fnpk2Rh/54y
gmDtFyFnS4WGiH+OGXKl0PTqvWszdnXUssisLj4qOxDlOxP9hvFOhdOFbsc1F5hDW/fxgMDge0jk
BZh5Tw7mobdj0XpW28RjTCLxuv3k0cI822pf1dgBZwoy6BheGvHUyWR4TG9OvT5orSP0mvJdrb2m
m+LvBur358LeRy0ZFSS0wIPLXqs3ERx/P2WCxjYznL1z4JZjWFqdWynF862L7uHU12K4Y/m4TlQ4
x5kOK11TtHDTeEOBFYUBRzrQqAgS3Qka+50nMpkbGOdpnxWyYErK65nW+fpXSwScjir//2tK8Qfd
LYha38jaS6kKbR12tvwe8QBI+jMKwqvCVH3yT5VB7yjCOYJ29mYGvGhWgiK11rvFxTl5e0qRFpe9
hPfafoeLl3JnqAeBQUvoHIk/yIrrDeoeiCqf5JK7udL0aObeSCNd55KVWQpEy8sAvQxxUkID5PUH
poPSxEWUi/lSnR3xdpr6OwDGfCoL71hL1pPcyxojRHA4c9E0Ox3CNzRHG3GCiRz2aRdleH3UqbQc
l5BYlBlhat+5X/128fK4nLGEvS1waPx138VKPEYNtv4ARGkc+V2OIEBCYAzXdRrS68/i9csXMAhB
4i/8uNd0YZ+owi4Gw4q3VU+tTTsxbW920zEMp9A+kEtVE9Xrfq7up5280ZJo+eCvqPN/wqP9T+Sj
ShB7t3rAnrrjm64qhU3uZs6I2FRiXbi1KSZAIu8cHT19RcZWE8A8vSChHsOAptVpj199LavvER4v
9LtwkeLpzH7lRdlFRtu34SO920TR3Q4qIpE4wvo9F/iAMnqnTBO4mb8qNDd/NBbCNGC9m8llzoDX
/kI1OW55HbvOv6FnV1HRdWBUnh28XIA4NVCA7ZQcNaBCgQ852pk+/fEky7pLQiQOYw/iJKfdhmAg
QqMXqq+Z69aC25O17w0kCJ7l9P7XSycklZF6KLgi+S/c3HMjnRBkKCHOoZJxYq5XRlHmkBkTBsJA
zGmV8ru7laJ0qw9QSSXmF8nY4uiHXib2/0KJpuBymrcrjA+fQOvttJ4Tmuze5ERgzlZKarKrYeIX
4lVtYyexLBooaCip794S0LzK5UdSSCDjG/sgJLfKvEY7jGrpwePul72jxcfTStArNCjktfQbRyUL
qsIoLbkMP2S+N8LygJ25S261paoAwmYFGjiII2/6FQRv2znf/l+VXGWZbWV8jsz1WktLwHZ7mj05
GeuHdbV/rW15HNbaxH1G5KVXzgaleS8YxTl7vQUU60SjCb8XyoFh20LEklPDOSApSnPTP81k5AZ4
+uE5eQ191Xpd2N+l/Mcc/+boB1KWZNxNdsd+NTsfomuFwE0wlUuVuOKHdKeVpglFlsyDDErfCq4G
jsk+wTmqWy/H15vaAKigpi0AjjEyDi26zfOBWAUUq9NNdjRwWPEC3sG1t+0fATMIOKTUrBblhwWI
LmLH8StnfXv4RqmtjTwoymruGwrlLQjgswcN9tlVv5vQbtjy81CWL7udblsPOXdtkBMqYAH5Cx0g
icn43dgTGIfiBGAFI3ox7q6QLGxlUmthdIjmxMIGvhgTQNLVkpfvNKE6acxex2EcQgx5rZbfBwHg
vbZsoVo1W47NVjHOz+VklVhTMKcW/Kd46yuvtHKTBXlRcBAWnBQDeh4H2htuZqHcV+C30VKmvv+4
5ZklECiP7phmU1gLZgTE7wt4X8/PiO8Xjg5k5yQm9It1p+JhwDEZcI0J6jCJrIQlDIGMxO+1u8u0
rSpnVVMfT7JoKWgWghBdvPPEcuxmAxLI/G1jaWKm2qC8lYm6n2WVkp563cQzGouE0nRhWQe1JzqV
bKyUjT4a7KVpjbuYzQsiV9toRNeVhquXM9PqXrVuDcmuOzaVtbYFzM3kQcDyxHWj0SukrYvrHLfX
B5MxmWr0PyjLaUN+H+JCS+5GlJTYCwoN7ShZZK5iduekVLIpnH5ZAML1ODJpYvL1lWkC2HFnsoRY
3HwX93n8aoDGqKc4u+Yv8064Bjo4FH0WQ6/f4iuR798r1jurjdPY7c2yy+md5OU+xse+j5p+ozn+
bFoHwnWkwA8sl3Bayq5Z44vwHCPrGXeZl6dRgcUldSrUxfGtzg7Zr5TNO5tMzg/WSx3UusVE3BcV
BGvtrIX9OlV2AuCfKigleYt/tRmGM7tS67Y8ZbgFb9i9CwPjZ8t0LbpnE1IRNlPC/zDO7PmdR0HQ
7dOf6UCyJzl9XC4xCITfM+4aXbhXOt//Nh1GOtt3QJ22E2SH/cHNTxEF/ufDJufDIvM2V5fv3Fyj
6uVliS2cOgYP9QtR+R5bI1SwpKgD172fDyNWTR4FZa6SvRsjMXqHARsejhBctsZp+ijQQDO2/xbu
IaMLOyPT/etd+yiRtytc/xZVdMPtd6o8ujbAoRXWg3AXhjVinBud34dhkZFhHsPagIbT+wOxW6UW
LN92B3BqmLqZhVSvO1iIvVYSnRuHvoRO6S3UkyFOmh0RAOkk1smHFA3491JsKShS71AWiqvkLBrx
VCpGSuiPq81qPVXm+wLJamEnX2gUIm7ewm2Zo39aIvPqJsHzDn6uv22FcTJbMxPEoBvPr5GsL1TX
fVCEUnw419GJk6e77Q96+FqsxBQLq3gfH4uixztfLJaM6fs4FSgjt6ssSU8qSluS/1EgsH4FU2tf
IPb0WrgBDZGSKTg2ED6DlauqlHxgJXeMJKqcX5JLQcTp1XpI+ciiDuIJqndQU0w7fqWPb54K8Y9K
f0WS5I44kVoH1mii04IE8MLp9UDg615pGE/ODXwSyi0WA+wf9vwi5Jjvy4gRQQUCXOjR+3zRgkE3
rOIll3Iuedqb6FigC/ZeXQH8PLyqqZXO0WMPIECTjDmievr2hYXarJe+VT71sf3jzFuHoC0ODzF/
ChHcxsXLM29ChXzc+Jhd59AVzoFKOcqzP9LVVZKqpRkXElREZfayutEXMNoOHBKyhnQgFSpb1sNI
xDx4xA5gQgwozR1HJ1dSd0Tgcy8PQEqdBhHAicQaIWOcF4PqDRMiQLweoi0fbbeZ35nvFoTkY/mQ
Lcdj3wscO0Cxix/X9tq3kCwZ03+ihVgGds/X5XB+ssV8eldfioxpZoIPwnevyvXeXK2SxM1AULhO
yLPs6ICFh7SIPfgPI1lO4Qt4i+dsb1KZH1zI7oG+//64dbRFKrwIZvlFop2TkE9wqMwC6HmpguTi
09xZvCwsdAz08HNssSnfHYsS0WwwbOkLmQQ7ueaYf44beAc+wtxiqCNYS+xdNOYNVcJGc3DMGp2/
QTspIobxVBUny/w5ANBcsBRH6MjwaBfv6+iZWncITKZCzXsIHrzN4wFgQFb5cvHxpblOli8fSCEg
Nrgqoa+gE4mFAF5JQT0iyhaXMjNgzlx7p2/B8M7Q/h/IGVjd99B3vVghN0dkwztNF5BEjQAwVVr9
VFd3/PEYFQEZoF0ipHeQnfnEDfI1RiMY5Y6O4stLW+2lJhk9gLD74Dm38GYUkCK3a81AiCepclD0
chohevGQ9iPFVyc8NTSimkZv55tm7NjJboLGGd67mbpMGK+jMlShrVktTDgaRWBZ46pnqy61GXwG
q9qh52UeZhKSscERXuF/J2i6QXTlEPkdJ9p2pKK6OZeQbswN7dw7LZNjmlH9FCsJ2N3R3yy0QK/h
9g7oLyN2aOhVuD2TcyXHq7UkIkT3XJhYycSPz6FM3xRqD6CbB/+QKcG7Mpo1tgow1bUT5x60ihXa
Se3FyVlDDiybloc+G5lJ76Gurgj1fgfn2nygLKfqXeCXGvRyOOcm7e5SbCyYhIUK+3WZNVJXx7W8
wm68wMksX5VycE8/6b9NVMRYRimnHQdydmx6yKxXielWKOKlYR/JkBPPZd551zwDGw9KaayKkPfF
2vPfFfgIceDGyc4Va1c38vWNG4YGYMTs4ZeUlaaDy+z+jbCpPqFLkLm0OUDj2H3m7lBMWjUPXDCy
Gjh0s2HQ03mWtDUIyt+tjPHDa3vSARq6d9VqkvKeb2zvq1v7jM6SfxajeeM3syZ/PLjiC2w3D64D
QNQXOI8zRTyR/O0AObNfaZ/hi4eMOybZbfXeYM+HrNWK6dxXEKUq5kNv6T7mL/7UiBWWU6s5LRqb
/uDD5KlbjJkKUzvv9IMG5iYieYCXazzCbKfpj85fz+6o669mt4ntqqMctT+JqaWkgyUw/IYqSRau
VHSKdFxGXWmE/C3B9FBo3khxguPPVEeD8SbU7sM4RgRtfi5jgWHhQR7HPuCNnJuWOAktB9/tdNtp
8BovNrf9FF4p8qyKLIaqLBKCOdTSv8v//ehmuDmUU891hg0piYlbqB4WD/euPbj3roWl9NQqLq1O
7UOj47ENKlsClucy8ZghDTH/qog0F4+8aVr38KZhF/kH/SdYAX1S3TWpVOu179lKNpaoRW3SZAlu
2JpgpZRgZMJov9QKuOCkgqTHyqownBdX8FFiYxtO4I/c07zdiDkGw7pi3HEd6hZ/k/pyICb73/XP
Vv9V/+k+nr0exMcJWIs5TwPQhkzOfYSHRTlhz02QUyJ7HZo5GcSoGpqa3MPypvZvi1bHfEK8bQi5
tmugA87hQoBBrxbpMXSvg8CE9B7RBwsCD8koPtq/YOghv1jFAw4EXKc1kblSfpvCu3I0cGeR5DAN
ab9TsvWgmwRqr+4eFCn1WNI3UxjtYRMSnjEU10pUDURFicNkRcZJSbTBrsTz9swdtnrStHVKiS7K
43YTAtskEDWApFGw6f0gtLQceVoCDUGaHqshUuKEJOOP+hSs9teXJEsi34ekCZWQMN8PiE466XSJ
6DKdcOqsaWqfm3cGTsSUljTgxbV4z2imxDdX76xXNZnqq3OxFHjV1c1f87W8Fribm7yPyrqeI6gK
Q9lp9OsPqvm7oYfadsQI79dCKyg/JD4feFb4NFdU4Hze+n0Y0H7MTeK8ZY/QvwkNdHqoUMGXs99Z
/WaEyJwCJtyLKfM6xyy30zOfWskU2itBMOhwsIGsO6J6zuerpEvFrPh8Fqqy9OTddH2hNuUoO5ot
pWYGQoO6FG+PKBPz+QW3xJVRe8UwfkLAXD9Hd8IDq96rrXhDTJNsFMJ8u2xKfZgkaEU/Tg961/7t
nRUKkrtARfMHxWjFLTDbt+Dc9lzS21hJH5yfwqtQIdPviECk3PtoDn5CAsQs5cAgyzeaJYUPrqxp
79qOTAoIA8mQXZCn+C1WOrvsSnk1T+heX2UCdQEBVZnL/g5wVEjHZgUiSEODPB4lwqchMjiqBaxA
Y3mlNgkXpg6Eh+N2Xr1aVXUgJdIUVFLq6mA9s+qICr6ahc0ecRKGwPKKJsJhT90dps8c59bMT0A/
ZkJ1qRD+7qfhW+iUsl6IF69l5BzVMkahXgroF7fWvV7fuNgjlsMxS8kr2erQOcIfB6qU20BlJbe/
CJ27lHRxmpljmWytSEg1Y67F2uzObdcFlOMWO2mUZOWocQALZqg0e9xpueoW60PNIjbZwDRPo5dm
7/BZXiVO43FuIVjJPwzkzO/4669EThL/dKVAxUfGR8upH10JmZfOn0iIxfi1gZWKBJxyTYM0VhXP
ZB9AsiX13tUgkq+nkJBVJIMJMULrpFmXZhaT/alzJ8QV0vWaZdwvGwJiTuMu0PbXhW8pqSjB8BFc
oNYas6f4OheAjBxLq5lrS9AYph+vhblnfRll5AxuBSUcOrU06E7p4uzD1f0L0tRz+KWvCSWAxn/o
W/B0bj5b3TwtqYftXTF9P3GH8xTfgoISX0MZLHfDL2/nDM3eYZXrfkMatWV/NEllyO5RqKYweqe3
g2BUv6IHudJGQqQunxM/+x6kB3jrYplr92kYVkHCaS1Q7Gx0RQ1OqK8nxkolvkvHtup9DFABlhod
u6xCcXl44mpbd1ZAF9EEsFSZAoKOHUJDdWd2N4wO9Enjx8vIA7z0vhhjkqGyfuIbKDlWry1W3XC7
41oIg+OrI6nBxBIfI+EM5CCxdrX3NeAILzkZdr3DIQkfa0Hu6ohclvjp0qq0twY7NEn5PgNN547h
f/D205iZxOXqt/WGCmOE4BXa6cIsqtcBN6dXEhzIo+AO6fk2QJK0AOTz9bIaxHgcNbiJoYO7MaeM
EGPkQ3tIogbNt+LhRC64z5xQeWTUeyBAbYPpLQ5vyjTODm5Y7m9FnAEhx5io8KuBY67z3wLpT+e1
Ppgmd+xd8Mfs0iRgEZrQqeW+zzjR94fAnXW7gk+7jUWvnT7Rzdpr1ywaSwUk/2HrIoB+t+ubAG7r
T53ATB26tG/JM2rnVrzT/Vf7sN5Imh+9/IokNDhVEqWNOXN/1p59T6bzzQ4i2CdXb5AHue2qVHxe
Ghi9Vk6wiEjrrluOi5uV1BzMEuAZrKnIAZSwOnt9Bcjqlcq29eGgxOmraRa/UxU0YHtHl+58fFFC
A5IC7tlTWi9rxlshHYNGoZHyRxtes6Rs7Joz2ZxIw70S0W+ngumN5ieV+gncoQZJPNKjLzNym2wk
pwB+Ctydi1jvqNIFE/Eq7pPMDJUuI6eDzpDjrzIvLn4TsRnC/7RRYso35ZxM3nwjXm4xA8sTmE/U
HpjRZo4nCnFd9YCnkFaB4UErQ2b2A3fp/7w0lBeMsVIWB0ZjJdOxJqD+Wm9l+luie2Zs4HtnFodP
YjTX0HyKzhlnjdO73km+EVX0S8y2sQBXAlfPB7Q+7IUI4U7Ggf0CreYD6ahOXza42ctkwiYTs/eZ
pAeN+iYNS2uoKWDBobfBBLF4TNZxuKHeY6itMNJSXTkIKySSICn2NDp+XdRfAnBaB7FIZoFgfV/W
7tRuXr4tYO+teJ6cUNV+Z4+NPeVvpjkXzFU9Pc+DB5Wlgcl5PmVrm9Vd1an4+HUzUvJFKdq9Gep3
q7A0TwLHHo+sb/3llBtrP4+FzqdE10N+R3p5VmwyH6mQjMIoba1vbPEJhohtURif/tAVc8rfuMLY
y+Jh3dupVmzh6urq
`protect end_protected
