`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
J4eOYqNYPAIizwR4vrfbiub9YoxukFQfS36BwMKMqLaqUJqFSKIMpjhdOPLsVPy+6e8asbXlWn5qT3jr12dgcA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c99gY2C5B6oLqO+vCXdv4hcVCrrA5qOJkVE55c2FyuoharC6SCvGcMikuOaAWErum9pEH99x1Tb6DGt9r1Z6bJQAeKVQ8jLC+OxVI1sdLmMfHD31V8Ib6Dezo9ucbvVZesCCuJNs7faCIxNmeamFC6fDReXBDhS/R+SMORGmCC4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1Kb++sGVQ0QrEvXFG5cSq/cVI8R3E4rX/Gs2KbYshFwYpuWxoHTc/RvqgF2b6txNVyNUPHyIc0YqkVARDFuLXnXUJmWMxaySthFCPtay/vtDeHgFAzyzLFjR1lH870AxfWOW7auMVwr3FVciOQsER14bTaCuN3UO7tCOcYcOs599+lxIcHZvu0V8i8bBvdfsYrwsXTJqd664O6cjl5YSV3RDOn+MmWkajiu1t65/Slm8zzD7TkNwVCJP3Spwh12+UBXnTUBYmb0pALFxcoFQ2j/+hlMYHdiSdjOfu7tzOPS+5UO5KWWchGc+wzAG0+Ijn2kyonk0NFnCbiyPLCk1Jw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2auvFXw7WnpSgEh3wRlMKqAGzPlxKalxe+QrwsRbxQA+oPRwHNO8trS34HZevcAttUsZgQs818bZ43zgKZ9YSC/B5yi/oZHbdQYWFyiB+FEEIXfSYBV5BI+m+1omR6FjkEVaTQGFoscqbv2yL+htfw7KLuPnVYudw9xy7bfcMIo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AuSptVdW7tT9d/C1LiHm6eNfduj9grFPC5Fin6L/aQb1l/uvC5tdCoGtSoYNBjt8sIPwIMeAg9UP/ZWu08v2sdlfecTqN1WX7PNIZG0mVbNsGs9IVj2Vsd8Kudt4vmEjBJtOBOE+Mph49ouV8qlZA1e8MwehErcne3EotK3U+iUSDAjOtSQFaixt/PCnWcxMAlul5lunQj53+601+F/y6sqXKxNWwfH7QcJhiuwaZLFLNt3YXXDyDmcfy83nD07CGkxd5BDGurIMQg12+VYctnopsJJHyc2s27JSDESEzR6YZVP/8OX3K88am3LBCEB7X8n1o4McoZ2lKU6J7GpjWg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98604)
`protect data_block
0Y2HF7N5DT4ZECEFzKmgfFWT8IHYZX17KqoLgb4S0zvRMxbMd0J4DL1dIAGXInUX490DDLgmTiSV
RbM1kiUK0/MCB0Em4n//8ndmvfqxlHB51m8PqBJ8RbL6tOeZ7WXnLmzS7TBa1P+JdT2Pe+VdOK26
K1t3cLeXMgmDFf6QGE1xHgQ/iICOmnW8oCpR7oJQrKB0W+Isgrw0yr0GZetkYjsAhVbjJ6KQAJom
N5BCw5kR/emJN2LxJBsHKjnMIFbB4GJQr95eo+/U/eIy+v8rkOyO19dKOrgjrwMgo5yeIAkDzlDS
5GntZFcek7gp1fSvrkNUiQiGiyxJ4BJnVjecixlv2XOC4JtTOIwmUixm9lx6dcHOY0n+3CIgyMSx
xEtUm9w9WcB98VjnOv4o+iCS0oZStiQxfn+R/uF4jdVWJy5JeIcvsT7MD/cLdAlzeAFQVIUfRy7I
UjDdJX33WkUnBv2WzFF+Ko3hqKiEplf1yu2HqfhxER/5dCIYb5ln9YDl1u/fRA/XdYVj9WAHNsew
4j8+w2PeLYouXVKBltRQf1TEmVEceTx+dKzuI8tekZRdzrU2EjJqowpM0DQq8Xf52BNoY+PNWWb1
2udOe+blOS2w/zdGcucR+HsbgSmwi+G31sWwfYjy1oF25sECtaQGzyUp29P1iNkPinL+7XzW+26W
cXEmQ9HNoCSKQUAS//go0Fy7q3pnTgWmmKfPATf2m4c0RrF7xqdEV8wlkiNjHE4W59AquGDJba8f
UpVIZnfr+46g33zfqutInmiwm5huKwn6pA46Ccxlu+H//z+bzus0/tgbX8thq9sqbrhovLB+Ql2G
eh90KY7fOKvSUp3O9ySnn3WdBQpcd//dLUAVekeShJWmVrkIJxpxzYJJXEyHTY/zexQX3VVseOIt
g7If6wTBDF+73FCH+Vo4HogsQRiPl1jj2r0LMBSvRkqXmiTearf35tiTmpk5+OJabwR8DjW8BOFf
IaMln3XfBo4zMesGUxrczg48omEul6za1cqbhTMscLHXJ9UW61+XgwgT4uwLU3BATpPFHiWG0sP8
hdvsDX3AuiepKtE/VBIqaa7CtWWd7cOPtbDMuj2uNEx67nD6HrSvfHVKfR3w+Vkqs/uwmAMmxBYU
T19fgxFDAM0evKNsLUrXtuCbshdX/4Ew1nc4Y/crGJH4d5x1M7Daolys16j9+VXsOH/WTTvKZcQH
U/m+GbxFAg9YdjY9mxv6g4ZMCjBzZ8zEM+LYj2F4Rnml82HgjApL0n+M2/8wXbYb3Gx63I8MQNVt
WDTIV1INQWGgNQ2e8hHb8D9Mbd7m+rpFCVf7G8t0r+R9haG2jslyqGL8ZdHEkVRSI9RYr46BD6Ej
0YOervbIBoJq+OsldYqiyxbJVJw2L4OG4/KqFATEyPH79Wy+RWU/Z2XZOhhj2xGy7O5223I9fdfi
ntMB1OwR1xFT3ZMoF7p7mycCEiOnR6ZfzUt1IXLmVVrCa7B6Y+LDVKu9dRAHy5ZrFSiv7VQLFcPo
nJW6P6x9GOPoFGD5aiXrId9uPtr4JPmg0curNWcLO3OpnK3pCA/LREJbf+lt4ohzUCVqwhPfCzsf
817BqavXJOeJx6FkhmjL7NpOVfG0Z2nVLuqOH/HXKw8ix7e+d30jIglwu0G5imv0/2PhwffNaeZG
Sy7D3O//fAsP6zgkTfszXUq3QQ1LmCkf2R3Po7hlJy18WXSMVFCwakEplRBZUgOALCLXbG0vQmSQ
unACmrNAoD/Glxbkwv/x24NxlaD4Juz37o5NBR8wutZ11hV038iQACBSP7ZcZGhF/4PuQqE2dj+k
J55o04NJTj4iBxzIRe1jsSsPFXvBsMggd9ZzzLdpxB8QYoZQVRmy94P/uk3owP8DikYoAnKlYArn
wQrY+IuvUY1A4pcN7tq86G6Zra9bM+HhrR+YKAX3pu/R0MDsuCbEl/OtpVqfonomiu50rn01JpZU
6BZ2OgqLXUG1JABqby5aP/7vTCgqbqJ07uTyLbfB/WXaiEGQUHa8iC/sJR3jQWYlfr9BNTJvXQrn
P3NZBdQl9IDYnpwd1yLfN+apkJRumGK41geLM/bfDNY02vax76MPvORDdg5BMIYh4GExcqIy315Y
CvUFl3EO7ZbpLfGoHsvp4SOUXqGhx9XDod+ApJre18IZPvhCCyZ5STlWaBVY+nvYezNaZzEndwJq
FY99vKWWSt5yvS/ku/EB7CLJY+lUDPKwVGWXfL1hAo3ZneoV+Cc44ZfmNLF6JwJNJ5b7PeuBQo1/
RbilK8PlIsHwP7uNrBs4nik/nzNurK9SPh5z9cMDUqcASsd8iJug5Cel+Gqgg8WX5giazX+ciWo9
dSbfifffVWOOo3p+8RGo1jqAXNJw2tgUE68AZfER1CS7LSiEh/4PwcKyB0EYuhzMfj4UawHieWa4
USfa8fh7jDD2sqCVNNeQf+pXmytF30lgXFZjjbsbjk2rl7gEDT/byLb0siY+9KK3QWie+QrFj0h4
oD5qEhZHsQ3GuHteEUcht3/Gb83EadgjoIICkg/8wW2+EcT4chwj9H/XTmOr5wT5LMC5mmHW/uGS
2cFtV1VbqozcCrCrZqwPsixLyLz589G/uORbvH1Rl9i6mc2Aoa+TzX7/9LOhRCoPx2ddvRMZvvWi
3+TfYj1+NueZjiEHAj029kH71L7pkNwMyIFgfV7hgQ1NjEi4CKm0yDkPDCcyCc0QKWjRwSplA6LS
xFlJF7Gmu2OKYl/HOsx2N62QqPntJpQE8khiNBusOv0ndFnMpgHqWMYf57/zGbgCUs56RlGPVgfL
eJeXyLSJinGs0aJMTFlFyGUhUzfpZaz0qykcrVa52K0hxsTiBUcKPOKy46oEx9N2OQYqlNLJhuFU
xcXSsO3wuMvrBi8p+60Tw01BzG9k00fbAaQHIfkir2uISNowHMS7Z4Pmz3bN7CAWU3X5z7LALxJ4
9GmSwZbARrLQifjLE3l5Xyq9vvOkZKb/7ad6VvoE5lvZAgQQbahb6XxlbOjCiiw3LKwux8VEAkqy
2XmJYJqW/5OzzsIJfgBem2nsjR+ImelP3evkl/u1ReysHdFqgrjBXojLjOunYfCRgPoeKNnss7hu
J+ZfkC9jvcJb3u9ghlvxti9QvNCLzyn/IVfX5oYl9h7GXMotkY0HVJR462nZl7diKEsRIrLBlCeb
6Q/wzikAnyZ0IIuzOgM3CsSJCFtHksTQe7dol91RPMNp89NOpmkaG47kp7GFrN4iGEQlbmn2PnP5
nlCphgSO38ZppKvJwhLm0acBJoj+rn3o6uqBtPKWctddHAhbbgoG4RuBAO2CaHxeT+tiXeoI8QqM
I14kUQXyJD6J4gTYVxHLZrkViSYEPVoc4jrre/RqhYET0aLw//DtVowDKQMgJgateQcZCO3SK1jQ
FfgxAaiG/NY0HS8wBnmkmPewwdWI0kOmWENMOY59cZXayrwnf7UOSbENTZDbpBYqVmZpZ10qyyK7
PPomgSK5kVbq45DNz0mLAVXm9E9jc9KQ2mu0sSxkG+lKanaR7dPLupfIarxwtjYKPnnbuZ+aIqQ+
DR4oOQPhYw/4OLI08Nuy1ivlfL7lW37RCAmrKvcaYREOqagSa0V0kkCXtl6vNELj0UNrnlfOb/kW
3kiv8U873dRZWBulQ91d31KXgG1lj0i6dr0ZC5TK6tF5J2UGFaehFl5FpHst466wJuINtTv83ykq
u4S/oX4DPJbRVcnvOuBJB8zhVQA2Ey/lN1CKlNavxwlrzcgumzkQUNELoJHaZWenJ3HoA/iAJ+Wl
WMH/PdCiFkBhC+hMTi1R5HCGgB9d/+blEJtPH2iXNaXPQZ3dbOWx+W0XXsgTjFZU1lEqhAlNbzdI
D8KcWX/HzQg39cT15uNRGFkwPX0h97TmWciE8I00lST0df8PGETE2NvmPn9LiTGz1qN2PqAz9sOk
RXIPVJQ43DPPcJfKsbIfcmOkDpWmUfu3p3/Fhr8b7fZE9J1FO5LNtDcBrMzuIEp0K6mfXwLCFcA9
5vc1mpl3gAUnHPLKnEZXtkU6dYr1Eo4WrY79xTo9IDZK8zdZhfCMk6ARbPlPxztCS/tQ/1Y08WmB
d6AJYyK22Tqbk8dwWTqnWuXH8u30EAKOJAUe6EOBZP1Lua6QXnQ0MahkLZKdTGYMcPNUgrPDmICM
FcKwThBp1mh07aY+1+YjWOLdzf6q6nB2Dd5CQKZkl6uJIQJGEbQ/gNzKq7K8EtYQASq+8HIieqd/
BbCL8PMpozxVIizQNelJLWOxEsb03bKTPkdyOv/sNbwo3UVstXj0JbSAZRCalBNNvFifGezlvvMS
DTnWJt/p9MAYBgZZNW7fw+lAm7v/qSDOIumYdWYDyron4iWZTQ7UiRLxivUY6+kMSwBQ7t+1BYWI
t5ZcpnfCtzcaRtbahYy5Mu4BIBXTs7qx9Z6SKkiPQz4tnYSt+iVPfoZTXANoU6A+h//lWt73yINQ
1j9V5y7hvqWKuB1q+qFzqyShdy08VZ2Kb0j9SrMfzkIEoaVBM5VordfOWkBYMvnmbGi5LCN+v4aU
uEVHMh6g1B6ZMJR2nytoY4nLfOmC8nlQd96i9cGjALXrZWsT6qZGdZ1DESYFvwdc7ecSyKMLPM7X
fRzDDtoP/NNpCdE+qGYfl7MBjIDuJtHrkgA49nGqCKoaIDRicj66IVBByfT+KF4nJZu98pYNp6hT
J6MRrcfY/qchWDLd3Y3Ajocwk6AeeJVy99UJMzM5O50t0FUX2RZ0cJ4d51Ai779jBl51tWncNrYT
sI6lSsnjSEZKsy5Zm/OD7+xq4LJKinbBBZVOjCKtD1RmsGRhXiFYq24mzlIPuCzEj3KBnsnOEZtK
zuVPXssI+2CpfjYSgxvz5FE7Ug+HI4uSHNOaofB0jtdZ3L1dAjEWDz+GPdtwM6zj9nLugToZYgcF
V2m3kr7VNMe9U35WeSdeXZQOqILp7eerHI2gjN8CaEL9FcJAwQ+0HKxauVEc1IbiLeEpy2xk1DSr
9KXj60Zpga2Ou59clT6f15pktZvnzBrqvgSxSyfgHISPCtAdpivakOrtdCxfBTkUtU/hNAttEdKk
s4BD5GZzzL6aDsST3uKJx8juZB0YdTgfNO3KzcoIMeXLs3Blv8p7OzHoC3AjvwjNm4m1dL6yvhrN
Wz32EDOxWnAlimQNnASjFrV3w3i79aRJMRaxPPy43QodipF7uaaVK56Rznb8cYhHgJn5cMHZdBSV
XrBZJy4Mh7ILUt8q8q4Y10FUpXv+0I18aX8CD0XSm53em7UHsEpk+KatcIZ38aqi0d35h2bWYqcb
8BFiWUyiuOV/X+GWo+76pKTEQW4nFr0ke0SAMcmw/dmUy3rpKLEacBEECk6zpFNu+Uwvd0V3BBh9
MVO3pg04h5K9Hs3PXUf9vCzQ0GBAVM/bIy34Mvez42TutjfamNbcPBKpeIfOJCxfNWxd0OK/lZmC
pQGTgWdHrPp+SQgCGdAIphGR14S7R376TxxW2LoxSrMWUGtGvBTzHEkivm+ZLLWu4dWz1VDQP6aT
Uz6QBlh9pZyO92mpRYNkXGiLSB0wl/Cm9+PAFsIliJQ5Xpx0qOk6n6k8SOs/IsGIZctrG5LPgkwl
yyrOS0ShvcxTHl9o0RFySYXUEzQsfCysy+5sqLgK5i++M6tG/hDLtw2W0wlUW+NiLbO9aJeQQ/ed
MPzmnwhNjBAsrShbLvgGE8Kry3EScuUnI71bkc2FLEe2xywOXrgic5/tCNO8XXIlCrwxGmr1jR2T
0d+JnLAGxLaw41qp5XAUYYxQ+Ad4Lnp1IkyA3VUky50lANm1cQTkXRs4r+UYzuyJhGY7y6CzbUo+
Eu1Qp4WKgwzjSsdYliPYaE1Y30wHHVH9l12qX092NMkWxmzsa8VWMRmhcpgKCGS3Ik5FLAAxlC4i
cCaVruBR+hgEDCssrVYZWDnYxq84r+x4pOnxlsvlZvLzMXH30ComcTBW4tuAw6M08FLFmj4BXl18
4dRFxOtqV59lqjOLWSVhTAq6B9Xn2tabaAd1IMqeLAUMHL7KfNqSuCMJVot1CmSGP4Aj9ofVU+M9
T93w+++O5xih/GdZOwzoaxNQpLXSp/vg++Lv2DM2AouQNKTRBFe0IAmK26Oa8BBF9K9/klD+JS37
Nx3coyf+S6aFidXFfP21WER1w/y2ZVIxfj/0I8u3AZF6/OF7SgN1IhAfj3IxhSkNd22KpKEq0Ada
IdNQYfLi6D7vuz61C/GZBKdl/8ZiHzsHMVUmmznb6zKwgiwGKKj6Vr2mh3ZMVMbzyWpzeMJdpDyk
jqzTPp2OfXFCSWlTyfQy3KNIAz0+1BUIz3oOxdM85COCm/jplSrIb3//zjnNz9FXRDH8/IfQmdVS
788ok0BXZaJF5nt4VfndCsmcml3xzEqNwWhDveR2tp6LmzmOMRwLJYRWvTtiunOeulkYKFhT/gng
Dz4OjmeAC0lDv2ul2wp0H2mzwKwW7hJUW/+FLoL6Ne3m9Z7YMgq9llb/LwFP7B3/aqTzarZS2Oop
MgcBo2SOlu8TViK4Hl4JMC9ox3SJZ1Tl43LjzkEIr78KnLRB9ODS5YPS7hrI7Iyefu/BjT4AqM/Y
Z8xx1sbyHWGH5hnpgNSLP5Z5lAmQeMOhGEehqzA8LuNEjoxKbAWXozbO06vHkNSeT5l/Ry1iE3Bn
Ri0yzSQXjieTwRzdLzvM0Yzl+3iNDV4wPMOSNdWq15/fv27G4pwNdcTAxBJCQu7p4WzAc4TFtK9J
bXl1r1kbAdnbPOwDcno/0+QiNjCTOrav6vRGJD2lg3m9xhC9Kxy43ZNRBcSpRpVvC45BMWJOKRav
iLKpXO7LTRHuzNYKhRgltXSBJD021UI5sunApNMQ3LPOe0jQApUnCUqtPyQCjleDeKbzlcqqQZSA
V7NfYKLqnglpOOB558805InWuR2PLF+4ryThv0BX75UEb/BbOQilUVDGRYbnmZwV6WCk6UjRQPMO
qFoPDjni/iXZeV7hILh0iAw6bkViOMDlwJBDl30gjIHhPfPcD/gaVY+osyUHc/1LjV3BOrHezHJ5
f6qJ8YEpwR7HlibJD++DC3KX+7lFWTBdNMWkAtIIko29Uy/NqUu6DfOx3y5ps9A40hgY83T7CWGh
dXdFE1VgTAwyOZcvAW8CGo5vXDNIJERgf/gQ0c8J6L7WtmcSdEdk+wmyg0NWKWN7TaO4xiy18tyZ
Uz8EaqJ3pVRM3kcnYzOxpkbT1Q2rZ2PMgf47nCkWsITu1FnGjjYrnxtu01EnXyxtL4BTB3yFaTRP
Vh4VoiMZvwGxbSO1IPEamJGXoQeTn9/uIq1FOIaOYpgFcgz1ccC5zCthrBQDmJsxC8oamwt1mRXn
oAxZdHhDtjVdsHbR3nnZ62ABAiwNXcuDFp/S6f223G9LZdj2bwjkMW4URJ+bjNoYCpYQ7AbKn0BT
8uLZq5sZ//Osriu3G8EyE5HnE4tm6gVouO+T6v3w/v2WFkPuKrEFcJf6rnJX/AVtGo9dNiFcEZDG
bGQA+lJOkV8Xt292GyDOZ3ofm7G5ec7R3NUkXewwN3Oz8mcMpP6aM8YY8VwOEx+yRXY7Id3niNmh
ycGT9T5C/LItYrBkOQmrasG2Auhxs8F44sjv8e7FLAqixW2kSpYxUudOAHaw1XFPfAAXaiAgUFpV
73g4N/B6fHf7pWad0E7DRq0NV+HSG/8oUVPU6xx3CWdyBSyDbcKi8nC7XU/FAFraxPWCpas1DcN0
4tXDnKHCrOErXKnDCs24XFAhmI31pbrZPdFQlFuroaLOlC/wD89dRT0P6sr2i08pT6npX1YShrES
WupH8Fi52cHOsVwuUAbP6Fzf9ml0JrhqxfDk9tpXHZUg8N24+SdvFyZlUmzTL60HV/5v89U4TSty
Q7J73o4HeeLCIlSSk4Ffal9j3Qlg8t7FRxxX0652Prfb88JX5d12aYqGwFf8Rvq5/SBP2DTFzZXP
XhTwEb+BL8jXvj1Ul1BOINsgMJoS9zjn3g82QAIB3z84+soa77VUJvNFGABqNj8RelBLVj2t6Xru
fEi8GVLKQ8hmEvd7L85gExPNYf8E2tkJxsQdOtrF4t42L3novLT1DnsK7CPkBhlgnYOQx9fZUSmX
lX7cBTsD98wk+VvAfKXF5lH7+GpLxBM06mgyv0mjHwM22p9bNHxmyQDhimJ9v5qg47y4eRti3WLr
bocZSUl+wFWRBPnGgwkErk4jy11UwCx3xYOBG0EyWziDR74vE834mCZa6SzH72mRqP7r5rX6gm8A
6QgrNY+d4NIFeoLWmO7BNM6h2eKmp70Nr8qlEvKQ+cfzL8DUNPTwI13+6c3GMNNd9ikwcYj6MoOq
Okc9bVVJJ2DrQ8DJt+dqzPsIPR7fZPqZJFqxNknSstyRd1GH76+Jv3zmNOyUaJ/0zFM/JeP2PBJ1
AJ4fT/TO5UNNse20myTPSO0m0950QxWJ+Q9M+pwUfVriTIowoipRklWFjHFHhCfL1dPvdPaHhuzp
GdtLjAjdV518WoJii6Un/+RqBhVioF2aRoONg5ntntZ5mNSD9n9EjKtyC6Ut8dI4JeMr+jKPda71
iEKESGiC3LHECKVlsqgXPFk/iVtCtq/S0vXU5D7DVz0CmL3NlurwMYJ/IO2gwIfHO/2AncWT9d1Q
xqhzSIjWLCd/Zy0cdAuHAffoIooUjT+fdOmtgFckJsL0sMnUbAGPWQQrmZ1dApFpLzvqx3rWDuOx
gQP7N215FPDQ+KYwnpLVpzKCumsUEpcPPv0kUPJr1PCU0YrnDHR5NT9OuC96c1KtPYXrBQA+sRFH
28g3xqjWjui4EU7Q8VGERwpsYTiYnmB3G20aA2vj1zpjJ3DLKE9EcMwu643CsMhIVNoSpqJ7+rd7
EKwjuy6rrgDt8q0xYf7MwNIOaxQi7L59ZIcqfRL4KCh/FxNSdRXMMNuvfZdzyN+UkxFsYICuBsmJ
XT3YYYwdetQKEjSc+5fRmrASYPQumeDSjVQ5ZJV7plZ+Dh9GqfrGGnLM0Zea0dwpf0bcouTlXS/0
SjH/0VFWpoqSf5x6oghWG7L9OXahiRwpFqfefsstlrZHdMf4RHYRUEqGYTIHcQxWsUdbqCLfKxC4
bJu0iEkXW1m+eADK1NTD6EOdRpwnnxaMAv8pm4njnA01n+iLT6mffxP2lA1Ay7F+G8w1SJc1vj3j
E+b4YN6DuYKv4nq2RcK2JXFGn3HqzFt5IvwJr0cNpBmBLsd8c8bkaHaDhKSHCNMrDBKmknGJpsxd
kWwNUFQfvIbUdXbbzK+gNoxRaCaudtLgOdLnPlxSiqiqUg9ExQpor9hiNzvlYRdafEGRv1sdnSUv
9bAR7OkNRbak01iAfIY+qVuoFp1pQ6ueUFZg8+mNueKWmiwso6mPbYybvyjC4+PDwRuUCUTt1ntb
7g9IJ4RQRi4+Ig3aIOnUlZhs7oJRgmaXPnHcT5Yzx0gQAR9J1/zYhwug62LPBQO3ZiCAq9BvXSCh
eOmRwpfnXlog1bh+lahsoUptPu2kppyL3rE5oIZxmZ+q515snMOuusN7dlQLcpjrcKh3qfa3kv1C
SSehRQjLUIZz7aq0PwnPRdAlJWDAK1KbMskN7J8DjPlH2ypVD18bt4TsQSnzg73yfL4uiunm8AWJ
LAz26h3vpxnQv7M9svwJAraIDHl+QNLC8xg8sFi/OXoRdbgpIMXqc96onIiv2SoU/S3xPx9Wwd0K
Jcda+jq6CoQsPBHFvfe5CLMzH9KMhcu8gByke9IgHrql/KFGWn048zkRux0P6AISmax1gjUT+TvL
/vSC7aJOPRN8RkuFH0i4Q/3f5MquhRnQ3d2OW8tksmIsFrBl61Vvf6CqShGJvB3QOAGHrt2yl0iy
NIgugCKDok3eWB9MxfbH6vq/LwHhnLLh00J8+BOQS5lL5OVFW/nEEqmAMFZ+gnO8FceG4xtGPdN+
2VrC9iJ6VxkiUkRE/l4pXg2fJnngb5MCoYgcNBREWzM1GzLOMqwl268Oj8bZdJOf5iv3xhM60vkS
xzi5lxvN1FAp3ZZyc2tzWIwwGlAA9HHgA3RHTjMujhV00NFZgaRMUNH5n3DoSdTgcOnrx8sr4R37
UP37RbIfxtA+Kslb1+CylYzlVqyyqPSGn/uxs+2r4gv5RsGW5OPairiuol+f2Nir/6D3HPmuYkAz
2dFMsWKMENdz4NT30mdPiva6FwfK94FcvYJnTRefg4j2Qa/BHKPupIXAczm3N8plx2lQkLaQRC2B
Tfn1fmMG7QesMjQU/3U4zxofvDrPBlgw4LrZA1w594KXyj4EyM1vIIfaOSODNKFZBmB0GepKBow2
mbXBPuMVOqGtgqzF++/3Waab3aXZmRXnxuYq0VEnaGnfdqH/0fq4EV9H0gGS+CIc7avGsby5tXzL
SGKCpwHSnrHVgJKN3TWCepkAnf55f8AVSF0EHoEzzsUczJ/wBK40rqMvlGqmaAJC+/fAnMiCItbN
8Fb275hL7Vlt5Hc25E/uQ2cn7BA+/f2xN2HE0oQz0avGorOGdhJ2Pf0Hr5bYuJVTBnxONFfy8adJ
a5iuDaB62V78jWjNsMSzMPHrknaL35Yt/PUQpaToF/2bnER2xHpDGw2tMo5nzTElXJz9U82sXfUT
vURvHZKeyLsQaKu/YE/BNooPTcBJ8sVXiAq6KBpMKKYPXyLMy5XCl1Wk83f8hNRlO7C/LIZy6qmv
vJiNq7sjcOdsug5EMx0RG6RsFO3ZJjPIQCIvOIahn3HfP3W52DEeGvmLVFE0xKxk/f6zbN2kbeBk
CeSXSa2hDQlFewI1WNKqjKi36m1D6hmVQq0w8TdICCbhG2nCJeYTeqDjhoRXbhxD/psOdetGq74z
IypjrdabZtSj7SZ6YVeWA/kZI8MNkHENVb43q90UAP4C40gQ8SZFxXC/YGfRm25Vt4a3KzUfJVrW
13lPF9XxjmOL6LMADLCl7DfJ7W3gnCMgHQzJVJSvyA3qT8kP8SNXx91a6ynoEH8rNcbEJyyHcTAj
ps7jcWAiRyRrPUf2iKvkIEsrQ1szjCyDvCH/q9PKokmH0ebkgBX2iN0BS1PKAVIvC6QbRU6VPGax
QEK3clsCeyjoQxETkHFuUIZkQeela0ol9p144/qDX49PDnRTyJvbeCNOAewu74xKI7uJ6ORgK91w
+BbQVOeLa4DrnJpSjpocqZAuOYRgTpd+O43GfFyNNr2oLlRanSpcGekBvle0giTDONUKck8ZzMIY
AjLGLeJ/pubjKIRTKtNR5j0lJMYNfdRkxXF/P9H+ckEYS3VrhioxRDpJZItor5HCPBsZurybYO7i
f1l1KKHNpGOGH1rAWl9VXpCFed5roOyHDtVgEtR94+E8F1JqJ8C/C9ea38GUvtbIGcUWAgUeIqnO
6f1NCREZEgZ3SQjX7S4wONbrWl7HrcrzAQIBtQ036QHblLZwqHZ8H2wWkrDeJB4AHRv8kYhpNQRN
fqZjR3VhgxeRaFee0Ag5FjgUlgxufU2xAY6NwpFKU/n+uRuQPZ885PWJn38LkuPS5Xk3oA71j9fq
Ijb30X9Cio9cIk/A7w7m9w9rBtGjIdxW0h/QD7YI0ttTIQeHnT0UADYgGHxdyZc1d4sCY+Ia5DEq
rYRJB8tTzmGrM6C7krxOV4Df1zuf3WUMs5rV7l/0fbQwMQVtt2WUmdLtgvNwpaIGi/9ap3boLrHQ
06LEhXGdOy8GwCcnBXJA4KbGe3PqyxK6nHNzUGeJo5LyeFhiGtDHlcU7NMnXuuZ3J4aJhNAWsXtA
lL/D++kap2cDg8cfxnnaT4C173TW6k/FclSek+NWKU/MzyUD7Z/6Z6/hoigFrfF2V5s40KMPnCjp
Rd132e8hJ/vHh6eoE3J+rVA2aSSoEzU3si/GkkzIYVJBQ+Ocd+drLhQYRWGoIbuD2WenQnFpPHnR
r1yoPmTGr+MObWcSWvVaNDozktAQ44PDTHwi/ZedSQxcxwPfdIXVY3WTiLv9q5HQqIdZZ7BXDnAN
TYfogdCfeKKzaBp5LtC7CmjSbM8GOym0Q98ZUb/u0XdYp6bVdfU4dSlcZQG+WV/5xRj1srDRq0FS
mqYGBYTlLHEVva+b2GKYzEFjIrEXNB82QW/ZoaNLrUnTnatvaUHo/sAW32SBPLlrxa64PhqqOieI
Lot0J8zF/VxoS0TbbkkNvbWxl3bvQRYmDhjM4+GgWgX13fpCYiQB/pndMZEdh/4SEJTXynyYnQn4
8kRA83vm7Kd86LKB4LAL5szmBkF4N08dYaSHuLEXXcEyWa6NSvn2jV16aA0X902uyskE1Y+kIZmG
xFbgwpfRCPsLjmAvQ2k92TYldGBaz/wNTjxCWrc1xSXSMIkNZaO4e6B/TvM4VqwLuHbMZ6Zom6bh
y6kLiUdpJcnjYfVTLUj+Be8A5oX7OWUJxV3BeqvtSIfZVDaji+YO7ySCqKrVM4O1P+w//bhAYrxN
9YPhLuDXOxHrWNK+aqsKMgB3sJKJx0aYHHituRi6PWft6mh1WJt4u9nMd5dc8ZnNwZB9M/1T5Di2
99Pfl9TzRbBkfM6X/D1upatpyw018L4g8nTkhffP/qzREbC67iaMgEGEWnMdvecVSDSqlmNxLJed
M79D1z6t4k1fr1IKdvMLQJjf2zdAR0qwon1CYvME0CjVL4WjHyulIPBem80QkW+fsWni7oCOzXOC
YvpP5u2c0Ie+M6v60bZBZ97WeW4xHIAck7s1dg+bcS5Lta49jCbDqcHB856TTUOvfuuSCM5pL59c
TTC11JlIbY++ZqN9BgeWVp3WIMIjLk1F3qUkKTpi3DEXkKbby3dFXu5/4qHnGknrVK54l49Vk9p9
0eLDu5YttV+PS4qEbCt6UPV0eYWksxjub2X8CjGi+t53n3yZz/Drc7pDm/Ztvtytiiu1ymsdEE7W
Jjfpdmz7DHJhIioL0bnUn2riEqzfUgyEr9t98EDMtvls4NE6IXbgfh3S9LkFR5HTEdRuQsyRAfDT
cUmrlIeEJlxbKvCs2iJUwkJHmLTRqZFodkotLMCICfgRy1ffjYrKU8lxU/5/TK7AwJUoRv+q5nto
6LfRlRwsojKnbrEZfJ/Ehb/x5/SZkZgXqs6tBe1QJsietRdq6L+awp8MGQyH4MqPICGIGTkgGoBU
ngVoAnbgRGabkxWjVUTCG4Ysq99zZ0ZiEfYErhDR4BOXIAFdfVA0tpYMm8bkhgC4C/LKkgCyHjzC
RRgK3R/C5S3So3RQlKs+Oy1kJNpBmy3khAaJeOXTW6xEBWxQwEpjZ69G2BE2SVHPaYRdE0qOobkt
vMokdAZ4XK04qE/Vb46OOAuf72vlkeNKLsozpOymUKKS+6VOIJ/kTQZeSerIq4WvKtp/8zgpk6Wl
ocYjBchqn5vPUxo5O2RicuGka3yLf7Wfpx4xMedM89aIdGAvK6xpEmuczTd4rESdSXUl56sU+S+3
nQPfhUwJJ1GCknOwtXS24lwNr2jOkvwWGMyyIjFKIpRxbcevswwxRx9QMZab3z5SOygZ7XHHW340
ocLV9hM+JNIVySCxskZzf1kyA2APST7yqUrNKYUqk8ViurlvTsMy8OrRwgfUdh6S7mMVz+Cfm2B5
a73yzHV9ET6Oib4W0G+qTo1PN/vwPTZha6abIG95g3ITSQcQDUKtZuREWNULi3SHDQPK81SJspRw
52zc9rufZG9EvfiaZwJA8iXcKEw8HYh3AecNrOCfIh41ZfwJq2Bp3x0plAL4GoIp3GWNbBKjdchy
WCafLRErfOH3lpZKWmaIBYGUHV3uJQvyuQXWz1MucP6LDsBWdQHyNr+sotJ/M57lAa7NFizsy1OG
vFK/Ec/+UPfqqjcsDCjHYUpe+APqgMewc+rVzK9T4qM0pubdWUGTwv5xNtmc1VnnZC3ICvb/fc53
q0dWyuNoOefDbpuqA9MCwjii7qWsIIm1+OqgFMQVjI9NoFz+3v+8eRLZlzgYHlhHTmMGIVjpLAIx
MYLE8hHK83vT/dyxuzDQSx5Kodq+Y63gsQzfWqJuBKCu+H2fEgHvKu2cx1Ab6p1GRw6eUU4ANnQp
8bZj8jjXh9QeTfKA6/DL3F3xNaqw772hao6mP78MiSPiByJwN68TLMHfvSbS5SUR9LkcgHxxwuqj
OOTBdBeZ51TSspQzcBvMld65tx+IBoWyLYZ3RjdlsZs0YioH35XHivsWwW+HWfr0hXY3MIjtRm9a
QhyKhcrj421tkTg2xeQse/GTCjwpMQva4TUXTuLbF82A1+5idwtN7lNb5ojZHEk+ZnLJYBONM+4U
kdLxz3LKjqrInW0KAi21lCS6HRDzNkEzIEmUyIXVZxOe5ROZqkSg+DW2nwAKvBX8DhU6Q0xcTfEP
e+48RoHXKoFgZD0Eway2/q4Ji06DytmAjge1IvQMIPObkx33Uby4cVRI33N8qM5jAt5Xo+wVFeJZ
ctZ32E+lx/QvpkaJbJdASvZRCLL5alR40F1uYAYt7Gmzi1imsxzQAZEX3PYM6g351iL9KLWb2PGd
5JgBwVfz/8SuZTFhU3vDax3RwUFMo2UVWEnkZNjIm1WWfzWm8XKAA8WpnpvZLdaQBoEjDev5Ar3P
io5hM9ZvsUcap0l9K5yrxeNmODQ/fj6qaTQFhPfFMk0r3LgVrJy94y/BuW2VeujUT4hm/E5rO0e4
9twoj2QbwTODSAJV0He1MwQNW57bdpo0KrdEj9n7kPfdZtK4SEpBQ4Ih6IOtgynCap6gO+L9dgA9
lhp0chi6MWhf0K3cODfFiSMmf78jVyWpRaOyKaWD8A0Mc8rGD3v6NJWvTnvcaRkjx+Fkzr50pVkk
f1eIzyCd2KJdV+Lj7QqjAaph5Rvg0bnVEbjYZjZw3VcEWttUiv/KJODAF9eTDVCUaWwQxGSxBwEt
M5o2iEFv3sPc3uRgec6TFI1xUJvL3fdbTBTaRG2Og8zwh1Yr0fPRDejZLsSFooReHzyiPCuDCTE1
LunodYiU0Pu0RqW6rK5EUAhj8WQmorz0xjZqUpzwB6GE0GEg+buEZN/rBCuI75c6LMD3ZZsOnYQ4
mLS2rVX4HDJ82tPBXXuzY0v9qA4D1Ik5zMh0x4DiD9GR9Cg70KuoHVsl16QkdGIHbCuCnUa8vKMT
5KLaSM6ioOunc8vMZ4/eCHAhdmXorz93u6bWFE9sZcSaSc7v4tf9sm2wKPXNvRlvzDuCrMDVUHbb
VxzIsBpKbB0X604AYeJvB8aBpDjm37Qpsc/O6ZiKwTpBMEbUpJlSgkHUXCGhU4SbwNB/7Y6NtTvX
OKbbygRZlckLVdow/nOdpS2WFqATvhVLTfxtxZL/kxaSXqV1aPKzUQ2fatxuj9sQaLwi3OWyzt9n
MqNtC6B7705hPUKXFhEQqIYM8p2rIYuRDXsKnB7Xb/wKVuMHR90pxe/oWfn7zIjeoMr+esaX0RgP
Wod30odJjVI2rhpdmXT47JDjze6Xs9FNDwM8A4LdcnnqxteKB4WBWa8b/iWSGBs71UmQ3EouojVc
bSCTqOMLFuCCskfkk387Cdam8ClzoQUS4vKCw3rCj4YF60/GahAFWQaIBGCJm9gkymLisDoFYLEg
58oKi8dWpe9hy8y2TyxtYTFgFU13dGk01EpvMUGSZ1tecf7Vp9AevCPPXvmkOo/2km6C7VPqu2lB
oyYJ4qaLDdprY+XrLnb3/cLR7ZilblTpFpSVqMWXY3c7b7pJqYg7xnqj9dY5+fE6wSFHeNU9nmHt
TNXShqWri324k4JdKaY0hbezTtVurQpvYd7Vg1lDHzOiQLN1SreFPxdsgpJDZ2CZw7kvcaHOPqCZ
bD1/7STBZfwMKsrre5u+PRP54J6dkov8Dj7z+pWfRQ/ZMz/qi3wDophNOcMgq891Vsno7pAS1SBs
tZvvuoKlgl5abLZHG4cLOONXOs70LE3uAqXD1TSH2ma/Ww1m9Wyy750MLLGS+EgwZmvERIYeH3wB
z3j0LSmlxu5BYWvhzhiGdnjvh15HJvHR0KGVeldykJBxylJ5+WRto++iRtuVhKR/u3ti1szpAVCC
Vt0NJ+wfalPG7zLaQZbubE4tII+nWvp4B+4dpfHsM4KKnvfcHwKCC0u13GyfmjENNmWe0Acf5jac
IVfV4e2J6j0vMCJ+EWNiaCvjgVtTUj014WjZ5Tm0OT0oaQFc7bmZHHkF5tWtMFt4iLZrIiSQ2KyD
IOUorbsmnu73Gij9w0ADUM6rSw4pG+iMJpbAbiNVSJPnv42u7rtoN4NXXwkVPxqRQTO1rk6L/onp
AWlVNh2OIj2QYoo92HO5tCugYE3YuaG8GjJc/j2xsrzzqC+cTt9E/x+eaVS53csfQ8JH8kE/3CT2
1XJd7gWABDizwX2biOYx/tgKeSsakyi0XjgaGjjS5RpR9g9kSAKofmRK+W9qmmRvFGquVZHVBF+g
8WR4MzlA6N1WY36XxjRRCCxrUshWg8cqFmnxlkZX280L2ka3P8ruYRcxHjam5JkfSPvHqxgAjkXx
ZOq5grzCX1b+vF9qZ85C9rBJYSqjf/3884qg9rMPrk27M/RsfJMdYqsYtqVnWP+Hn1GCtOUD2xqY
pq9ZenHePeS6cfl3L4cx5ur29KO+xYlZz3zH3ac8H9LqRgwZfUUBRM6PHWE74GDBKTotenIvWgMd
NqgF/q0bCYlZzvAEY7TQyIcZh+9gRJmJWnQrcI52aah1Ob7HOwCYpmuiKwV1Bf+ynLs6OhpxR3kZ
LFPPVdLivaisw8kcc+Qzq5/60zSRSY4a3fu52spJjmt9a03AOsVJcUAWmYX6nLlubXYmYUHa/x4S
435XCoD97SCG0dz03gLwjNQt6QPeTP7sEfqHqhWja3kj2v9WyoXaHXOVsPDgEEpsFYwgJwA73XjE
UO0v28E3GNYvPt3QyOIVXg3Q6QhYCZNxRiHqp6U+URvBJbLsvPSc4ElnyYA4yTurRbNOBImSAOpO
VhHXsHyv977be4YwFWw5Ysi5P0RpEn9frEG5r7kaQmorY8tBaq8Z96ctiEkh+P4vCsUYDxEuLS8Z
ZXX76o7GxlnEYgXSAbfpBfE0Y70TLJMpCW6NRUUil6OH5Gfun/ie9xhzuuzszzZTR/FwKKFcmrGX
roK5/UnPaz7Wh4v+rq//BcAXyJI+4FJwd9E3fLqf+K0NF01SWXfD79rn3GyNN8OU3tdCOqnI5LbS
SCVHeUJyDeEViFY1UsoCLCvJTnhnI584rJIZsRcPcHph/RyoUK/NzCkaavIILwbA8T3aPe9d8FO9
LF6krDCy7TfPxk9gO6abuCUQj5ceF/Mcdzj6KLY1pWEHJFTDh+0oy24S4WEZKug6YOZ4UvkRmbS6
Y5qkmgMJIXCNcQ0hMMbxuP4vuOsRMxTxlpZK8mz7M76HUN46h2mUW5eCwrIyIHDFt2jufYcQcl28
3TCmDdptpc6e+X+sVAi0LycW5scNteiq6LLvQ3Z+3FbSLYz+Uyuim50IhP+m/uVjVTmMebpdlwEx
RDDc4BkWm6Hqct1BWA6IIEFlDPzv4gDxIFVxgx8PAH3nKE/pYUdqLOw+Ak+evZBP16qYSX0HW+Wi
TGHzRy0/UPmYrYsk2E+mYPDU+ZIENvbDQ/vd61HYw+4ODDIi78OqKpoIbjJ4H6MQWjz4CeMMpC+y
m1NfgOQmV1/guGHdqTldX+IZbUFtYcNHP5uDbdBr4LJJ8WCmm7urjgFabN9iTS6Ns08++ldMvwff
nJC9a6Xi5pnV9+bJnlEq5Jyqse4gmYwGxrBBFhe6QOHYb2OAvWHDM/kRCShJQSTnQNjg41a1KwM9
OH/rCLjptSVI91HoD+k/LNcrgWOWdxvBm9uoUY08ZcrN0qt2CTMxZp5kFVOUSYGwjOYhOJ9Unh7r
mnaps0s0QNvAB4JvSnj/Jfo2JnMqtgcjJwJz0GDw4JnqdY7SNpfPAEAC5xkut8d08KzQEBERezPo
bgxsRZ2PvhTjhR3JpChJ1K5jlKdABESIqufEXS1ejycwFBcfnhla/0rqsAEL58l8zo1CxOQ4wkcL
VA934596Ax6Yc2cE1yPbEefxZexhZaV7nPw/Xvxc/GGNjY6K72Mr7/yii7lZ7ahSBTXDoqN1nRox
MPdyHcs9n6nlE4Z+71631PlYeeaEed/kljNYI+Ddg2jqN7krgzvwMoMkYBf9AzhTBniSEhTx6Hnq
x3aqC20vVWvUJIv9s0k6QxYVdbCAOYjH6+GO0cR+y9K3WO29OxvTp9z7C9owPR+5Zz+NWg3ZWdDA
k/V9Q+T7fx8QwzZ3OO5ht/uie5xZh8RqxgxoX8YN38aAPDJFqMc7/kZg37V0a/ewdzg5Xr/QyoQ6
eUw/VAFawkOt2H/kIJw+xN6qtCkoN+5YUUF+fHxlef5HtITVVMy7zKwPUVaJ2+jL160ZtpydO3Xb
ojwE+NZC+lZdRoS677pgvaxFUuMy9m7qsFuAIDlNKsDCsn37dWtazJ5EU8iRN8ZpfUODmTmHybAE
4Rh/Rj70q/o+okUQ0sCsswHWQML8owpCZ3cKkWw7Y1gqyBvjOy3sr8d794dMb9Ae1+SiBF8BMh+r
L+J8Qr9uSRs2deSMawliTpRt+HIZTcjwsojHuaoO1ItbzFULjPq3xl9ozyYLIr837zupHevV/9TB
Vyb+Vyp9+6UBLS/TWC/9mr+pkHNQYOpIAlfoaRacONgmZ+YMeA7E95VdsHMdUdwWCh9n/VVTrWtm
LnpXTHTt5nL5/pix73TA4Z4m0F0npklmVJIycfILoYHVhI7U9bicj7F7uvOtl8CZlbY92BI3QJbp
mvV0Yt27v2v4Hm/CMYWc7IJIbjhBvPcgxTQ2OEkXGhbx7U8CR8OUcUH+TooBwieKZVdx46Ans1XB
Mwa6iH5ZXIyaygM04Flkhlf3vacAWwL5D7KsYkH2fJpNrhFqLIJ8w+fzlrNIV/TVFiIDcndtCBSr
B8eoWOKBffvViteL0r2ZZkY9hThxqD+oCnLzFn+2oqEmzvZ+FSWjC/bPg8F08w1N5y2c+wyQVjAG
pDIMPopi059dHPzFLjzBt/f/RKg+qgcfr13fVHtV00dY2tuQMpfjGE9mM/KLhF0g1pUxcEazpPdr
C012LXgmOnGgQd8y5cPd+ociaYUCqf67a8666zUBGEQPF1UkhEU5BK+Jz1u0Wy8h95HCi0V8/EzA
tbrB+QVxVHzQaTSEWTICWd1lh9FZ0vN2czixHijGrLmU/khDEZDRvpNu6CkSijkI3EcjedrppJ45
w3LZzzNfiva7MtvfLlpoJ+oS17ZjiXTsjYOApk6Y8mOFlL0ka7cV3AduTK2rdL6U/CpqWwr2yqEh
sCYvF+XUXBafEW94xldTmEzx3gXlWThaQ7TpB2UoKJR57q+ddhycPgD2iZ/HLQfGT9IZXrxKLQIK
nOOxFumGkCF0xPL748rqsol4OAWXQOOrVcCgzACe9VFH8zx5Jlq7CnMuN2Jvv4xGO5IT0+Nommz4
QZs9q3llujTn9WQTW+Pq9Rwm2z3rftHMvr/FiX7SpkkRIUInSfwBuyvKUZUxjeTZMYGM4S2JoqtD
a2bQZMfUY7pqUrDm+5sNJiGDYd72JS15HpgyvEh952ARntd3tcO06/ZRUPrwMJ7te2yuFG4AjawO
h/DxBl8feeKAbjnaWWcLo7kCRKGIV0wQn2RYvGtReZMCMNHlRrFggzW/mjt+lzOuPeu0ecnL3KUu
NJY1bzufQ8yt1ffi8rD1cvgBzEj7gM77Hte9eLrGXjU3d735EejM09B9RJNuea9O1nebVppAI3ui
e8lvXwa/7Iewmj1x7X+Ei2nS49ftCM6yqVYTkPixM/Umuj/i9mp3H10ZtjRdFyryVyb6ZNa8WcDf
aDxGZVLHGkl79xiw/0WPppTrwQxBMh0OoKVZ5qDYNub7ozM3pxx5mvQ96yEaN0IG4n7tLh1a1frK
bFhPtqCgko8AUt6ZGubfrKl8aN/o/z8aChwXTdjlSQ0PzFO1X5yvQh3tKjbAoBvQRQcVU30e0xcL
lm0jLNaskefiwQ2VM6MX8ICt59IKpPwQxQ9DYVt9xUZGx7h8Mvt0TxOb+RpQm4quDpixc9+tRehv
1aXnFcHRSdJt6O09H+dzQFQP8soccTNXXyVLaX6ZF3zuHxn1ERPvoM3VvsID4bVCJPPDqLSDaZmz
hVRyuWeUYJgKZoISjznMI8t8vREjGKyUX8+VudF04VeYDaHaJYQFBIkRcdN15XWUettXGgcWU+5j
Ur534SHEj02RYBdTU52WTuGomyzNsb+6tfIbMFwcj87Fd0PCZyqd0JJ4ptY5DnO6Myxpj3aQkRVy
MAz++/Joj/s/RqGtdyIT7vv9O2c63tkpT5/5AEETGruJXORe8t6aT4OpSZPjyPQ/ByrWS5UXuJKA
v20DH74jzKt5pKiCl1uhAOSin++RbqvflEfmeJ5jM0QaUEs8I6z2/YUApcaWW+A1BMiveQeZDYFM
U6bpy3pzb4opKIqtcxYmrKEv1Xh7nicGkH2MBiLg6gClyEv09eddTX6Li7cib7iS3vMp09ltMTlK
R2xZ11xUwhEu9Dkf+mYJqu8HXXSB7yOCFs5ZwBYzxJ/Yh2LYFRr6oY5TPiC/8I2MwubxmtFUwwAx
xZoq28PGqy0rBUlKbYfNmCg7f5N1j3A7GwFYeW1NRr/4rfsyNU2bhUZp6f0+n1f82Xf22TLmwZWZ
liCQiIOAzyS7eKsU8ewDLcvaHHw701XzKhfoVCuveuEAT327nuTLUDoorb5L4FyncLm5sd0C8TKU
HrhpXoL+fWVYBYhwgFqLX3AyI+1M3or8OqHotUSVEmxMg+w2/HemY5ggaI8micNR2fLkZpFdL2jj
Y7mt5ffqZcIdAzciDZNt/u+fw1P+u8/wKeccmKN/wI8VAzvI9v06nxOTZYLwqsv5kHBpsz34XX5H
jJwfnn08vY/e9wx17MA1OsTXoQjd0nrAMAMomdXvAty67B+683e9rdYMIZDYb2YidfGE+mGimN6R
Q6Pysx+FWkcdIAtFH8ygjoGec1hyD7HQeXGNsUmuEE6gekhzWLqBDGS0hVvqcRLbmxd1vqka3tZ8
n25eNeV+nKxFwG6mmTHuDmT+tnBqHBpuMjyvxvrJ4D+J+Oz1HeuS9xEegdbOh5nlh0GaMLhchNwL
8KqaoNZbxgisHxwom1TWWkD46mxHsx+xA+Q7x3WMa8yo7HFatrNySyA2kVENJCBWxh/02iJOs/XZ
MPWaaduf/G8GG2QvOZh+kRgyayOOHu0G1uWnnZmEu2Bnrdtkt1c5FLerPr5QvIlEe85ZjoRbRZt4
FXG0OYp0pAtcfqEZqf//EG9tpafRzSUvL3qLFfch/oY6l+XCsyZcffKi6JWTaWvPIVNF/k4F5rpD
f4HRXFEfNu8dZ17HOFtr6UIlz7e4cK0ec9HFdlekaY9AADW/123sQAxQWu5RBXb1TgfMtE3UX01x
d900LlNB0D07EDGVT334P459zxhvaTjeEcuKY0yCVm6C0Il/uj5WsW8HH+rH1b2X13chlA2hn3+q
xO2KVdES3Q9ZYDQWBRLgtw3q7ZGkytDXwBAmeC9VzrqlER4kOMu3JfyyldFsoXW8RLJZjbupN5YB
t1/0jy5FDGtK4yyTjXv+8p7CaqtN6A2XjXiMCUzhpYzTQJ+zXGAP4IW2okwfqRdRqm5j3tuCZSEL
gQykW6X9tSIBmJCEs4lyzdSvCjKbwCEFaGmz0i74gXoiRbnpw3X1P2+aJHqJMpxPb6Te5bfYouDb
qwOVUpRw2VCVqyJuvNlRHS4XusKRj1sai5Ol77MrddSzlks10+iZq/pco2lBexJ4fPY6DEZE02IW
36XtqGB55Hq8xZ2k+OERYnSb1NcAzvP8HSAkx9OiMryuTM2E1nVZB7fhrPjBNFGUmb9F3WuuzhT0
9fIEjNHsYJlioqBxW6jl9x8ZSxelTFm5t/W5GzULo4DYK6K+ALHEAeR7ZDQgot00yQ4VWJ2mn08C
iUIwj5xZ/hlFVCJijY4oFgYHRNYnauHGq4MZaQ7qC2iQoFP8CHKIFNQOeg2kFAotXO0jaXmgcWt9
57LhtR+PO0p0eUX9jYE5ZkwNWSGmBSNYumUGqSws/fzX4/Z1SM7zHt0YFyLsFsZ8Ek6mzX1HBU/z
CKPK+siPe+FMOps7zPYrr996F4vSNxQP2Jas62WR2luX3sRT0F3ZDY1pSR5jnrgPSrE2lBoT5UBx
3HjDgPZ5bpz1l1S93MFV8yQaourkKsbGgGDXFUVInjbsYdw1wB1o4JbghyvlLOn4SalStQw3FhUw
4hbY9Jp2PWXXfQklKg5pYC5V4dmy1hV8WHX6UrTyTvfjMSHIKVxxum06MgoU6yYqAAzMAUpPnNV9
ueNhTTasvxdHMZMUnMLKExPD40gOQq6CVxMOsNBpsiLcatTMhdZBGEThXtvchnamh6DOm+czXDAo
dLkhVz8hhbP84q2RrrOP+/R+2hQJjUCW2XeIBdwcMvp/ulcixs+W8FYK90j7KCWFRSkawB4WMj+H
Vao9iKBSNpZLxd68bndW1jTxb+LIee+wpDfFDHPnS4G2Tmqaj8+gGgqa02uvYfhqDhMW/8FADH4s
YwQa511WOreNROHl+Zvp8f4KqAVqLZcB+KLMmhZk5+9e/aQrRDzOSCW509H7cFxrnvZRcd6Sww3w
XIy3I6JhWHth78nuywBvbg/NvgxoEJ5FvkDjMrNefSopcMgmnuygGYS7iQnZhblUn92X6Bg7qc1K
cRMT96Uq3DXkvbMFOeRJaX5xzUOqdqpOYpzIXRZlJeY/4uhforDppFGrriZOziQOE+RRgZ1u4iVb
ojvJ/Y6DgsnAkgnvuDU/mBbMGRlJp7VrdFWEgPTKZryQKx3HHhh5wOEJt9RojfNkNT4nmFdU2AJ0
GEp1iJwLXzPdZjT9nUZRMKSH1y8aQUIPBL5QujlYU5pypm7gdYq3KMQ/0MlexUvrk21sVWE15gze
3JZD4XvVc7Kl46VvMfWvBLvLW8HH4H+6tEfPluRHLEEHNuJ+SkBlSDcF6uNtrDmI0HuGWSiPCrPF
z+tNMv8Nw3VKQuoXDkZnrJ9yyHZ4JIhnEmRC6dTrmCWWh/g9EYosCu1BYWMTqKlcMMc2+7dRSfvG
Xd2x7Pq81+0I0KiepeYYETnzW4Rg2aRX/mtGqHtIHg/EH5E4m4bighUq93d2yyJABYP7tfosAUZL
I+fF73/w0Qu+ejjZ/oK0KwvXXtqrI8H03vb9dI1a9icGCCSM8OZD6gwmUK8oe93j/hyENyuF174S
4croNn1sxz1A8dAWr3YzDP8HQnudnjqdDdWljAcj+fHnkqXRfNLh7wPjsNV1w9j9JjtwXTqM6sv6
DQckJmOAEnxmf5LWwj2SWClteh+rzag3vKkY30FHS7rbghcniOUHgn/BxRD4/V5SIMG4MXkd3PNN
gLKl6RbQYbM8GyCDnDmDrsFdwNniMfgef9yvmaRRQ9CxRIH2B1hb8QKmvbZAI9+0wxG6CZZpB2eL
kX9sEc9dTXPPetDQ9h8RZhUAuZVclF+QMVWC9CWaGBdq7n38VOsqeXsaLk9gg0hgGwUmb/nZLLQo
5QxrrFBrsvZ6Lg17NMcEgEQDmyPnHqfDF1LB82flV8z6YIMabWTgz6ME8jJE2nkoPgTvC5EqCBPz
jtjeDwVyt9OvcJE/Z845aBOKhGB+oi53TOUQNsCxAiqg8VORNQggm8BI49V59FuSGajiMJflcaH/
JL0Dxlew3/0C6cmYx5sXnaEcFT7RIGnSDPSDryJwcHg00Pttab1PFDDwHTz8zMGizM72pQvAguqB
UDBNVLjDudbmbdq1jxQSQiuBzjTFYjrlWREHDkNuzEqJtrsFl7eFdOieCOx1GwU1JJjK3U76/fD6
0MEd5M1wYfU1U36d61IZANdmDSBb4BXYeWXkjwC18VJRANUGUhIa+y/jGH+uwk3n102aCVG75u0H
W0/uE0LJ9C5fUyBRvq8PJCMFnlewS+2ekKYcY69BH3ePaMmZDvBxG9wXOKTSJQGsPA+IkQ+ttQJk
mGpnt4JGVRBzJm0osJhL+iksAXqXMsTNjd8+xxblj2BtIqEn32yiSWLLM1B/5bavqXV4VXiT3j31
CQZT1FafvrY7HexgkUNZjXrIp+70Iyrk8jJ9ur8rFybLiWv+/yEgHWb3SY44BvhqF+8LGONQnXTD
+S3OtrUKRZyNYWjOsha2sAEkLU1m5S/r6wtVxEzXkgC3xEzW5A6+NUvrzZbD0H6gwyY17z+07gbW
Hbou3o697A5j/UR2YCzRE7Tg7OTM6/T1W3ouAyBuFeEFAHHYCHYlSMKBZj2gEm/rUGyEcqcJs3SP
0fU8MmbEFa/uOebHdzF9DWIz45p9e55+VvHFYGPUAQh8zANe4Adt2y257Hpqyz/zfhYNvDsNWWAq
YyGO0xCWMtKiAQOJ6ScKvq8L2CVS4hD8mqiae4sDZUi8LrvZbVF5PAmyEeQG1uK45cYK+HKILEWj
I+w2RzU3HiUvHs5S/RJ65n743xymnvFJosRmEYyZKubR/TvwW3wGlMkZ8FMlVQuxEXwofImHpyNO
pdPy7cvZsHC4If7sW61Doi7tCocJ9Hxmqa24+cZSiz+EAcB/L2Vi9pFQ+t2aqzITak2OMB3I7H1a
2q+BpHQFC1JcuPgwiBSs3LHy9ghYqv6oulTtlPG35DFz9YdKTGsIN6rewZRb9QJLu0qjhF2gfq2r
z1hWih4/NfY0dvRszgbm5r09jdGUA+YM0v/ecDhj2ZB8WE6JSDvGVpnDtp+oNU/yGGnT6hof49TW
72sqPf4YnVTLJTtrIpa/A9BPUatg3EITw/d9O60GRT8waU9t52uBr6by4UEXdRT19n2ufT87sjUj
xFBV+m2dEA6ciEvhjp8l88usfFAfLOz4QxiLm2R+BOb00K6g2Ujg7eWIzAd+BhVNIs2lMYZZhRl+
q+TOhlJAQ2tmeIEMFUKCKfzFSkMGmsmS/eFd28luePNk+DOOC47QCs+LtIJbB3V3BGHdyOx1DK9p
CRfkDeJVb+FzWUctunPmfDIrz2KcTmk6ntmygiiFamw7iaNFX5axqe1hq5+xLgOXLWEvhbLgaT/r
bXynWUEK71HCGzUftXi8pqgZ+NvfeRomxF9fwIL/WFQgPn8d/6Uqh4720Bcb3WaYPpQZutYh0lIz
bLAJMih9ucIWKDo2D5+COg9257x2QRZP8+4r0NMLK7zc/a0tjG21hPqkYgBkG3Fr6+7EldsFJTxI
7jELBfInsjmoI4gdNiSoNdNuDbROhUUNwXXQqeFLjxTVtcZVIiWnwmeirfEbk+ljx9A5TsVvqEE8
BFLOgd2pbrDCs866x9rtLmj884z9qjM2jiTUjIywzBb5zIwvxI+AA/pMeDQZ94aXQeU38QgFbdc3
b13Eb7Kq9n9gcY1aNeXdgh5C/Agvhr7JNfCDzT/2kJ44DTTORuzUhSw2HwQqSilQXkJ4uvPclKbj
nSwpFq4QqqKdy2dvcSrR8CTJ0FiwLdWV2FIuhcopQoa1KLg8lApJ+xA4iAWFKjJD+rhGSz3/CqfP
kh6yyunBUehnnDWzatuoAHXVWLe/x5OE+BNKjBcvGgBRmcn9zU9FiegvEGBg/spIiRjW3u7BP9OG
D3BpmCqd5DngQpCys91NyZ5InZr+/kvNLBGYWJI3bf0x/N+MULphP7YClNS+27O1lhfzh3HJnRyV
Kg9KftBzWD8hzVFrN/bf/eVDVV3ME8D8WiusOeC9nfJb+Z8n+QIGR1OOgi5Q/iO/mKgWV8rgQh5f
bAIyYreqApRWw39+w8ZQm4zaXMmOQSgX7vJIaUMyGgLPVK8hpwCQplX86hvFxhGFXcwsKOrq+7EP
6MkWMQaYpi5dOLIS4AZ5na9QLXrIlteC68DB0w8h1OxGPP80Te2h5N1Grk9/P1KDpOb6BThT9ezO
HcCwWwuT2VOeQc5Cn9T6y4snDZIunzlJZB033BZ33h2kbkCCoa8maJvuYcQ2orIfcjnNjvJwtvTT
f+fsnCFkWNHkjzmCBjGx9YHO+RQundKQVGFn42V/avRgMUmRVPOJLPKmhn0Fb7iAAV971ezsv2gp
LxgS0H5BP1/WR6k03k43Nl+rJ04pEnI1Rl0s605NBs515cxblpbj/4gdZ/0k6POL+vhz5pE53RE5
mc/B7kChizWshdn2NlrR5dF11ycYzT9bnqQ2d+bqrpwRv/xJZh+s/9TkJ4ULeIVsTwQDsMJNF3xi
33VvhT/wyPFaKKFeO8EpJdPn0WOy6IiimoPThUu+KnCngWImfqATxZfejuh28fLqFdxLoOm+lvIJ
fT4UI07RVoD8xeoMXEcgGwfBC7tmV/3VhgYieKwufF9zhmlBdd9npaEXYqG3jJ0EGlWBR1gcoB76
mX5C3X/7Vyr+owE/HkreET387NzAdPHfzCkYmwrhyEfXCpbqkt2+MJEungrBibPY4YGPTNk6LyuM
sfGELA9/jsRDQLVCzLFrN7yYF4dxXEFuxwN1Jbr+UOAYddkLAM37kcaxqOiylUF+ILgjKB1WkpqD
mEMhBre0dl64kfLudU+6JyrB5DCjT5Akz0pZ4zrYaavVaTWzOyds+UV2kXmBeBhL3qkMhfmQ3etK
xP9RlDsTiWHQwSkhnQ7RPoU+0bjMqpDHd5mvHq4WVxlv/vDYUHUzJYwruxnFKm+Qr1lSWg32ARIr
jq/kM3FTgyapV+C1Y8OpKxjDcV2Gzf8oBzj8hYfS9u8YppLUVSsor5RGAzugVpiw68zhLQ7IBh8P
Gx5WCxJOQgApVFvFp3fQJwZlwY0+w1SmpRFt/YRHTNuckH7R3Broye0uoNnVLLxC4QecPH5wDgbW
AITwndNnduepMu1ChbMMFKMY9I1FeeicS3DrgU+LINnHa8XH9AwNH16OtGlqb9thUSSwCizoGacW
vU+MPs4AEbVMr8Q9GP1PZdTU844mdiLX/rH+03nON6evCvg0oMzqIDXRmX6D1x8qle7Rp5tXLoXj
XOhGqksYq0dV5B1lfJepwZpcSj9JSX0c7zs4cqQ3fLagVNK8XJfdjF8rPqmb/WSzkxMYuW+xl0lS
PYJXvM9Dvdpz0WFmt6HQD/Q66yhqHjV2LcLyr70Y87AO1noM3ouex+j3xE9WpEpOKUMpYjJhkG7a
siRm9ts5B3XU7j4JjCNHzj4gEdkKJkVlqMct7HJ8um3kMm9bhDNRGXJPO2oayemtVa+tOpAY4Agx
6cvWzkKX9cYx0YE8vdpGJwXa4J2xsk2ubCvJAzOpKQoOQFFRCeLcvw2baC7nVupmPSsNONgSfFQA
uBDgb8jE/rcWJ19NhRjUHcMR/x2bDANp94TToNEE4/3fPNmkAMrmCAdsO3ArFn2mkjrR55TybZd+
eAVdMMgwOBZiPDGesdNBAKgqpZCod3seOxoDzevY9zVUH5V9rZFJ39xJxSMQ89bC5HW3LQi6vJW5
xCQMd9mxZzXDpyiz5xT+tUXlNnkuhupB0hDPen1DCft8wQNzsWO0gXBAGi3Vcgzw7yoCrDf5EWXr
bQulXHZP1hmYcPS94RKBsw77L7Qg9ovnFjO+0XnIcZjk64SJlVnosTtdDRbz5a9Ccc/WpgaGdRKo
rpP+ToOyK/nyyQukFWd5csydnDwQQujYon8RFfYngzmvXd6Y3A8f983dzbFkBl+nq519N2PDK/tx
B6DY4xVuEP+qMGFA3lwGvzc7Q+6YAJTjKunUCimNWDzrlBtgMY2vkVOA3OdAWdl3nZsY79gEtX0Y
kbQ+k0BGT9Rbt11bE8PZ3IddPM8xh5h16rqUNRd/gGIsdoUmBAyS4xgxUYJCYg9plFvfLsZxInu5
NvCK5yqGzJemQTYlSxQd4KiNiNntvtphpAu2P+Xw5YwVdHEeZ04yZA8GiPR1z6gvBb4o9N/ZMp3D
/y9fXGa6W3RD/+yDIRqQ1js/XA9F25s/XflfOuRYb2HmOFSUT4fWradOQmfEpMusLr6k3XEwU1yW
kubyGHMekcI2wMLsp4/t74KFGX93MhKcxKC5aOsKFfeeG+39JY5HDjm+xeGNIoGpoQFLkgpOt/yv
ySpxgA7T1jElX4iNGXo0RSobxw6jWLSAuW3NOsnT/68IuZVBvn6YEPw+S14BaXdUU2vRvBlbIUj+
DsL6q8mr11GSY3100cB0IAo1+eRS42UWPZYEBotktULMV7RrpBEKR835z2Mhe+EzD62xa2G5mZkT
/0zrbNwydMW6QQAaoa7H5xFNFlzJtUvZGx/CY7cI/6wT/ufi1ThKEoOTimX0KmqBp3/KaJrgmRBe
AAa1M/9ftqNqLEn6+CEh1oiGdmjjYjHgpew4MTXr2RXwEm0tQf4y00IufV8x7mCB20QqKC+rtmrO
MiN+wqziRlA0JqRka33G5hQJWJ4tILRAtNGcLQoOJFlnwQfh5dI+f5MAHa2vfDlFaHfe4xntHczZ
B00yjeAGtYrf7xeX7zE3wGZfFAhI2W2Eb7HnVlfcDFiMM2RAOMZayxWWt231GdT7oMP0w0Ik7GMV
DLRtjYFojPhCEXURtTrgGQiIFJl5UM+k5432HeCSs9zr8eOCKW5VOhvzOcmVl9v3bawxX0fSFsyC
CmKkJqTziba+zhAPwA6pKkbc0eBBjDZNk9A8ebFZMyzSKTb02QKCdkQb8gDsYJ/r7J8LtEdkXTYf
+2TSdgcIndytfhmYV98ox2S5uBhPTBUWUxout8VG5hkxpK4cgehX3Z+H2PNtjfNUrP54qqz6dW3S
4GSr7AB7iPFApo3x/SVaVuGiphSfV3Wa23lfHoor/pKh03sfrcGEja3ocvKm7ZzTla4eR8vhmvZc
OddZJJOzOldcw07eJaI8GL7/Xv+VYDwesiFlEHG2MoLJo6hxxrIWhdQxfXwhKTj/k66d8cKVzTgG
BvW4/285OzZn5jvAZJZs1UqJ9INymq2RhCR5UkZYeeEiML/hQXA+KxvggZDHa3URXXWjUkZN3PTz
EaInmRe6+iWzjuEvd2IU+ixXraEzkJyjYa7CQX9sCnYcBl8aNZ9yFRO91WWdAyfiJzbxanWm5Tl1
Iqo+znFhQacmHofQ8zQYhIa0orqsxv57fQklGwGheac1MbmAXNc3gTNLsfkyNj3m8kMZBUg2FSYD
yrEzfiCDJGCqkT8Shw7X+OcI9QCQUv8/p05kvAUvM2ucPm6pZ9ffRLxDcSztcZDE/xx+xRFc+AnD
SSQQ4mDJ8mZrAv1j3Rk4p9ijJrIH9Z7eCVYfU4p3b9GbFETq+P1M9tWKTjMEj41k0YutVLkzKK9B
jvqRdYBadjW2aWhxKa8MBwEg/XLCO05RNUTPdtRuXvsasjHQSTd17O3IysDO6Jmzwc221Ky+fEB0
ruLAGyt4tPO6iNgDRZXWKXbN2t2cKG1BWhdf0nGIy2YAKqojQbToZ1GTkdYPAZCohYOOPynbavVW
ysBZ/y7o/hk1zGW5v+8C4WZZixM6p8xqrgKx11zm0CDxA9WjD4hnBR0yYlgXlygF3U503wqkRZkO
koEgLI7SYUxO7zr49tYRUeT7awk+RLakAXr7ImoNzwnHBztViviTXhaVs0deAfEjhU1589vcqzod
RGLTG71vtVWYG3mG17OdRXwhxYJawgc2+yl0LngZ3ZB3w5mIoidqjIrL5yyCkAsp0sc0qFUpgv0T
YK/Qs+n6wBUORq4lC+wT13pjNZeluJ6mnPumTrGhRBqYnS87gNrGXvBuonjKwQmJqA9CJmOpgBaK
DlZNbsUvb4W3At1/OCuBZT1qInBNoBgDjYp1zbiKpf6k7sVC1Dy+QzL5w4Ok88+WsvzDLOZtNtvc
VsGb2rPtAvODPU6uXP8I7txABzBOsJttScFE3OMwBX84j4QkX75VvkURIYWb3f8s/5pZvfimiHFt
A2tl6DnsAWj5EeaTK+rI7ntXpn9EY/zQPDp1zsyy9mnOenPpc278XkW641j/eTxBEO0qo8UYn6jQ
hqlULrHFVU0vJhZoMRarrBfXhZU7gZjyDRTiAuLX9++A0+zsyxnnuRw2vPaadirb0WU+hWJ8RvT4
sL+CJ8Xdnb0xeEFubBfOj9SiCcj8pK07jeRGPznWe6Hu3sO8MGTOfjgLHnSxAQYZDh5o5Rs8fy9m
nP/M+0HPkSG8ZvuFzkoo+5jQ1e/jNSYWy2YmjzyXAmZzY68XpXafVYDr8Hcp7sI8zTarxItsSYDZ
j+y7wAGRF28DuFWM2wWK9N6892mBvhYP9NHphT+gAbaf/ULm4vjQB3mYqNIjV1fTXZoQoRGcuzOh
XM6274HKZeRm5bpx2hy7rNUQ1xyH7kDKYfOTN7uT6ZsHsuo958ipSvOBD+WiMxkxXQwAf1EAfxHC
YoaJVAKlLg2Y3dBhiP7IKw85vw5NE5l4mEIh0357bQvE9FfzU8VJiBd3nUBU+VW0KBACReIb+9fS
J4CWIN1k00J86c0/aF7RgxAR67iTKKlwqB8JK9SRAZrJK9q3ggyuOasESo7ZKNdBo9hKBvLAbJGO
9Fi3iFO7Z7Z/W4dxW1tdhKEU31zIXtDIm5c4Ygf2QSQmL4eg01ImEBEW8V8/3FYXFypFOWbt6fYr
hw17RG3u9TYsfSmwsr9t58l4BqMrxO0FkipImrBP9dQTO9sqPERsq5nouP3oYNtq4VKqxps5n+9z
vp9PHfT+RkFWBAp93FY71tcypNCrByDC4f1cY8nm+G9eOk45mq85b+xQ8XktZMKTqP8sm15InfCQ
inONeX08zOmL1HCjMWlNqrPM8EeIfXsoDFrU5r5D+q+XZLw77fB2kL9EYk1SFre/jKJD68vQsXvT
rZxX9+WFbrzjny4EA8INAHL0hXkLxfR+OkoYAYlJoCm8adkaQc/r6cTa4vhPLc7z4KYqO6gxWA5L
t0ONUB/sz5ifAkBLLKpbpz0AnbrCrR8ojlF4osz3ZWoSr94NUhOXfGz/L3cXimD3nKQzOF6okWXb
RUCEGPhkWv3GJKXZBsSTxuvwlJ7bDkZNAl5WBfgbRTZJVfOh5OlTTxg/zbcT3g3LElM4enWbfLTT
CMvF25xRHpdTprFXaVcEY4y+XzPsanc5iBMDsFw7Zgh9IeO+wk/LNfq2hR5h1PEzMFEhLQsm4c03
S2cDLtrF/lhPDG++1LwD+AI4tQcNcTppuhn5DWcCy/cKBBXbtl3UJ0SIvUF4obJ6iskVe53xn1Wf
ETRMZvqKPbZEP8+8IZsh0FXklx2j/zVNE8wcbwEAG9P5VywC4lS68/s9plOAJ+BSgWkyfvInBIoN
qif+ux8ZGXjOcbAB9HLDCRpVVe6uNWzF/v1LXSfeng2B6QgEKFaMwFQn3vzNNcU+iBCXxm3PJaBv
ZrT3+FFKUW/1Tw2wCqI/BpfF1rLa3Ng4HCR4Qm8ym4FOUVKlp6YZukRfLrNwkbTiBlY8kHqVZJaH
lGdQVGQxrLQEWISkPX3+qbNvO6Rnkl99+2mizzoyYgg7OccXdTZcgQPtzGWilWVFrEiV04z2M3Im
+cnP3qS/64sSbKfUAXFvFzc6Q+8AwGXipzITWWm0+K2GvLu2ZuAFIPnrY/PoprC1QgJpjQeM5pJS
0ki9+PqnC/K4jMWn9fsNGeaCmhaodK6Xo3LvqN1jCQc7dfVTnqTbwwZpTI81wfSFpFG/1cqaEU0S
lN0jR9hw6x5Y19sxn+Bd+nTIZdi0DQxMblcPi4VgWhBD19G9F+4RBCWo80IJGW8yVZTwIVmyzHVW
tKzYz9Z7J98Me5HPqqfkAGtL0mgk9eXrPUK9kTrV4vXWc7quKYEzYQxyZ0lsD3uyrUogTGk1314j
3Nl+6hKMuFa9nwV1yhwln3/xXV2ZQ8PP+77Jxs5fR6ggI5WnuHmCdkjsNRNAihWM0dh9eCYmg73N
3420jQMaGjqd1cV3ZI8fTTiobRkSjMwQII0pSSo/4D3QYs4OJTIRGLoA9StOG3l1mSwOTEgn3+Ta
XqrjPlCczd6Ih9NFjZ5pt8KaujSwN96Ydv3f7YtmdngkeYB8Y9SW7sSpL5zRzaYM6fd6QT1hYvXl
ASBdb8Ut0ClnwAE0A2d7N99V3KqZZwUl0i2c6GwUcgV3ULPA/d3OZWMb5nMtKkqWOa3TlGczOHG5
HCyN3Ld3mzl/eugut+TNqw9/riwd3YqsbcNogm3KXMdq/B246QmDH1yrx+/arAwIod97ZVWHqKDe
dAJCweuEIW+3Nvdiy2ytRP+ZEVKtdTvR+dIA0Cz7pVFuBGie1aU+uJHCK6m7One9odwiwLbZpgEz
9EzYyHWZ0+MsPGUQApq+G4hJrGTsqDC7gWAcpfB6suvfnWdsjCk/0ixTBx8saJ+pzbpgLdhZfDdg
NX0uaNjpU4YKmmu9H6PjN7npEekWKkk8oEgvNTy/njqOscFVFwnEdnF4ctXjU9KwNuR7HQXBpZbG
JaZZNi8C/fh/Vs04qoOtFWjRGvitmRfY/WB8UVlt+veVw0fnR+2UoOVuqD10yT8CJdMsnk3gtWqD
RcxByrrZY2djGgjudsmYqbAM7S3EKaFc+mcsaoBAFi2J3mSAL1w3bnyGCp46S8l1q9c5bK138CJU
V+Plq5/38VJvDPmB6znkTUEV1cpbMWMRXz8AZrwMKKeqG9l1f8HteYPXrCIG4HcD1qNR9MaPt9eZ
Olv7sMH0zfEDHhr4eIoGne358OtrcMpz4E90RLlwEJODiisx2NMnC0o/SIhazFAkd0InAqD35CU+
1Yfy2NUjLZqg5r8opmgqKbtp7TDzfBK6qCejx1hseonkWq/G+JjRhgD0ZX11x5Eo2ooQ9qgd+Pnb
AGP6SYjL4UF0wij4LSp8YmLTD/sT1K6wevjLViL2cGOXIOtQ0ysHBJsNDlvK3rwTG5pRAD1Ec52z
+ZJfSYeCtwVdaTd/IN7VFGISI2eN2VfTPrRbHzPNbWCS2GJkPdStBFn8Q9N72ic4ZNri6CpuuWwl
BujETYFCyCz/uyE/Oi73PkZ9NpKcLfhEnOcZvdV1Nu6U92XW3Xsf9Gu7IfuuADX9bgmM8OxR47J7
sVekVppUlQ6ax/4fQcG7oHGXgQ/HhCaL6JBrNumpzdJ3IlqCpGV4sqQBt2KSP6vIZgzQScj9+1kb
XiBKf4A61220jEXqLOQR9gKfem9bP9ECWqNZwOxQPYcfUP/BZI61+xEowuWoHx2HBuc5fET9d168
3rTD/jOKVz+zV91XGTFWeVoyBg07V/s/5ER2Qx65j2PbjWXMY1zXLBFuE+6pJ+JlRsps5mXfbQnF
H19aA1Yb6h72/K3gcO8CE+mhlSo87DxvsrNm61VXrGb4g1TV6/ycsuhqI542qfdMrVt7sBYeTsQT
gxfx8AGTR0fYUPhnrpJy4wVgufcSJ7lF59B2ErJjiL2lji7nNNuQV0IC1PTuIcgTMdBY8fzwd48C
VjH7yokuR7RA3ro8w+FQRAT8d7K/F8aanfxv2TnFrr+1UMg0EHFcA7C676hecGcBzZlLFn7FOP1P
f5dkHi/HOcZQMzOrXTJbqBtIvl6Tyk7UiLcl7knXSSNXQWB/vpEAehxRsUnQ3uEzmvSF9q6XGeDi
I2UqymyoUuNphA9SqK6x+6xqXVit/ogp5KQjDR7Vp7BLTJ7HU35/hBTVT3bNRAqUGzVGjvL5opSG
t5YyVi6V//vd1XvKLLlEJesoVYujUEjXP6uxOYZfP99RPNsotkvkfoz7vAMGh+U/NX5+PEXE5ttS
1Z4deZEdfObFBKX4ChL9+psoJIpns7Rw0vO8vy3Npq8EVvAepFefhy0TMOxA9Uc+qKuu6oTmvVdo
dq7ICEX6LC34K1AvtkB07HAursB0FnuFvAU9YNSB1Pp6AKboOrPBnRqHPLg73Kp6JAHGpHDR+5AM
qJPf5O81ymCgqX79yLquLLVjga4idw6j04+FNw/BkiLtX4nSYWc7E/znib6LBfAUnA7Pi9qrbXa0
ny570yO525Njzy3puPSAevZ5mUJ0Tjh67Xh4AO6BoVLwXHaETM4tSPNEhnxSjvuHNvw8kG0hoMRJ
MDz8yXXk1+SQLTtQXqBH5QjV6jjcPern9NOCZSlKgzAmfyGgJSToSGc4QmJ1tsUxu8SzkqI310Ww
/DX3H5ck1tB0p9l0TRTtQcOaXobE5jTuyGgJc7Rtzv+7SAU8qhGwBTRg7sIr4owkw2x50+qtVPQ3
6nO9pqx0VgQvAhbtRKAXhHTGF9pM5OY99IRocMve+TQn8nXqKY2nPnhR8+GSwCCImznSMPw7T1c1
vDEOBN6BK59rg0kr9rUsleGjlsoCEXJ+N7h6Keh70TlQ/mXTCOKRDTfucIjLKZFe0XEis7hQcsqP
d6UU7QUHdrLnKu0gbeyI+HEQGKvnrpBoMNXEPJl5vVExXuKX9mLpBUqEdycNs19bk5NMMr32DBMH
BRC/oaUECpkw7HXjJx2cuz+13Z8YDGHwXfTM03MjBE9y4EgDLG9Vf+i2C4emLbxqIX3LIlEFwDXy
QISezuSBB+NuHdShYJ0Fi6BVTUacxXG7ohYiF5rUUqt4l4ZiRsooE4Pa9H4K15K11TEu9Bd5lN1H
YkXawbqw8nJ9WsGemif9I4qMMmFhVrU7t/x3DgHqpvih5oOdLBtoph8+qFRR2SJ2vk3e9IJS3GsN
ze92+fUtjd6YBD8+5JPDfAPXKm70SdYZu0wQWeyUSpw6RDO6Br+NVHIydA+qVCthBYPjocPnZKpN
5XGdF5cl11Tz2T2sYmuVU632XIuiURQw1C7CRsrGAnSFSgFgNBRdXsISa+a2wPw0EIMfKHjPrpwD
Rorpfv/BHWm0lJ3HZ0O/2BOTsUq6714ig27McXHT+YolLqsbv/LC5+6mBspFYddsi+7CCduYIYZH
qGVnpRGgGF9q8jaOh5Zt4+ks/vMuVTSkb8R8D4dpHhgliHPxu9rbf2FH+gw9auKpQBq+U4goTve7
Wd1hWBgHHqZ0FSMgVd0OjERzyXTA2M7gsrLIq4Qhliv21uNYohoFxp+ZCfB6yPkH8L2zayJn72hS
T+DM5Lfgy0k76ey1isCQK5jSATju5ehJKx9D2siIYZ6hmDTmv0nzBlrX/ozjly5QNPQ+Sh50yjNw
DDlBl6D+EaoAEfMt2OfmXtYXhx+UJgXcZJlktzqKng03CQfqfbtgA+KGxDCv/wc12H1KhdSCsvKi
liFoZCznVIZRk3NEcl4bnkTfRmsdIsW4MxxlfpguuSBhoU3BOA0C1p76hqL2VyMCgh2UNmI/ML5F
WLEb0fvtX1BzBoD8QtppMtLwkK6h3HEqWZkm4lL6BID5oeGNM+onX9mKoGyJenZH5niBRig6h+cN
avPIMuYorEnARYZLgeJCWHuKtTZ6zARwqJO/X50d72KC7+lsdtKF4SWQOJkAxKYgSPLr5HwwG1zT
jlFsdbbDSZd7aXUIiPbOACFGUoGgvWzQOrtbd3/jsfZLoc2+fzw2i2QtfbAXlMh2UwQyg8w0dBDS
6RSdK/GufLg/a87vjQCRepMtdinoA2213XEgjWRn/BUYzntl/0tLqBo4dUMPa2J930NHtCX7BdVl
l9l65jyzkHHejQASy3jM/4Gj0/GWn3gfc3y3izrfP03Cx1i+uil3xUogw4byqQ5tBjzVLAy2BiYS
+d6P46ovQnOOK3+52BZemrhesYz90rNnJOy9Xof1c/6FH2ZW4BR/S7UuNtQA7eWoMSN5IQxAO/AA
BxtlSdPPfKMVyEREzjwJpBB2LHdlJtf6GgUwAU29QJ4+5VgLrf6J4Ry6+TsnBzWFefwp4JuM04se
yeSPPIXv6Gd3nFKvlavJNxMlWuc/ORftyWBxOrMFIizw0QH9YSu5CfKovDgIo7bSshMNAJZ4WxAO
Cudw5EnqlDbdWDpziW4ddjTxi6tO1da14B3Iv9dLhsVwuxDdn24Tx0evr5dl6rf8hAYYhv88B74o
9fAjSstdpqyyPToOqNUKHR76DJrMvdhX/PeoPPCYnj02CdeKmqEQCfwbWv5LD+E2BiMylQEj4ceP
+ydbrA0zxHUzKKSw1ykQp0LBNq+Os4GEEhOgZtF1zaECsWs7Vy9xaD8uW8MYbtabbRuZMygXk0Mu
ihibPo9taP9bDIzgEjRev5yOWnPsnsk5rgdufezoEH4aTfeEEaPkE0sfDj04Ofjq/0nyvbO75T/o
8Ybu+PhZC8FzEmuJl4Q2J1gJ/iqnR8WzF+UtwFFN1ZPsy1pJEJNNSDCNjmanQmuWvn3mUkyg801y
LM/PONsJEsFGMWkqZn8lK+K7TVgGsRSdDUVGRLZRj7P26H0ziDIhZqeif3e2SL4LthQSD/65Tmng
SYj574WatzaSClCtJnYIgSQnAS51GJFSIRcz8vmsELlFBWx6TqNJrmopPh01KKHAN4+3OD45FH11
lQ/6sQS3SSouKvUhgdlWc1YRB7W31a2FPQ5F96U83mXjZyNg9+0SYJZaPZiak2Jj5DmeFjdrpkfY
Mcac7sK+kqM1IahnfDP85tVrvr5YDbw7RfWRW6YauDcxhgRvVtLNpsdijPkpkHBn8YoP1kb0FAYa
6UqdccD+gUK9vHMdpolt3xa6cw6WV30/IO1rg3R/ZcxHcqmDbTLLhwY/JHC5cTAB18Pe+9H7yS3j
8R2cVFjemZOhGSeslsnWWp58nTzOIXSyKu07kImSpqTR2bHvHjuotXhOPTmTnqhHsYlhRzZB2AJs
k0aNw8FylYEOfTAEnDvGGJg+X1Qnmigcuu9K1L03b9Bx4lpwvKQUNonocHgxDEQP/vbVxY9ZVX/N
j7h6/KD3Fi/pUJazBQssvy+pFMf3McUkkUhrgR8InA21DpGvjIylQ/ORxoBunvjhm0Ras2mVeT0v
YPEAlnSBC80sn1K5EalQYJQzKWzwwUMzIwElmPYlE8lJNgHMiUvdhQ0uhaxxODJS9uO3pliOQq/o
4iVof1DCOcxPpTCYK14X958hGoFzMPLDLjMvZ3g+bn/zMvI1l3Sie1NIMSmHDhV01ZkOAhZZs4oj
nqThlomoKB6UqPr14mPhO1bDsEvYeM+wJZO/M+l3eSntB2AQ0IaOpkBoyoMrRO3S9deCxHzyAi/n
89Aq5FkAtKJi9YiwiJfSxj+DPRxokz8Z4ejJx8aFoCy/Hrw5JqfRckT+eGkZnN83yy0FkVy89ugz
vsuaceiXJ3CYGoie5jha558nDxnGJZtJ2L0zHy/XiowdffjzS76jZbMt4AlA+dkVVrZyyN0YKoXm
hNR6zN62lWwi3guJMaNpgNfac2e/FjlbnMe/XJKp3I7J2B0uFD/AmTxtUL3mkekNl5Jq2z8jlxif
gA9wJwv6lTfVYQOYKwzjlbfOYD0qebZmgslNrMZpTqpH4/KmfBd9JKTDumjzN7HwCy+3ps0TVNdC
A7cFIbqJS386oFJ2wmLxpGrYkqPDPnWlv4nacHt8zz4BjqfBW58tJ15wGqnwMIkVZAg2CG9zTqg9
yU/vgT8/i6A+fFxONAj3ZjYLPaPb4cg0APBbmHCxmXaWU8suRJITIK+QSDAjGiSgKQ4UInw3b8X5
WTTZogbz+mSvefZpmVioSThoQOpq5VDKXkXw0c0I86x4emtzgq719Dh7XGa+5Tqpfal4vlWl+poy
futkrB+kMIa62AZF8W25nvyZOGVrz+Bkylx6iDDmX4XtbLWLwvkaWA+Gw0EJGw3aux4JCcB5vixn
bNAQlk6cM7I/ctHcr3s31Cfb6hmbm4TLOjuUy2/APSURefLnS877wxDmkPgpz4IGAnMwz+BvQ3xC
W/5/TvPWE4htnUw9tokQCkCP7gPVPS7ZHjs5AYJU0+hbakMLUXOE6V3J/QS+gadadaigP2IMvP72
J35+cs5EiwqEnnNdeZOptKaQkg/4JMYHN2DOAD2TX76o4kD0+JNRmAW3CvK0pnlB2mb+Ms1PYt97
H20phQ/MkZJaNdNS6ihHyZYb7J/mzWtgdxGZ+dYkJ67OIBdM7NR0ClcQH1XnRiESoLutfwgglAhs
rYhQlEPS2XcWnNgLTibJUWmPqnn9N33p27qJs+nqJrJocx4vDS/HWNUiMlTzi3rjIgfQ0DEwPnIb
+YMvj3/TzUcxkwSSRCa+d3pFD8ivcFEayf38joYCLsuukF812OSoKetH1LwKUEnc6mGdoGfMs3vR
wt5KHu474vDF4gdKyvz7eSq+tF4aP2UZl13U8QIebt4tLwnkvSIKXcEuAycpon5jOJWcfPSYepST
7UQ5TswseTQ7Heb8dm69kB+YaIwMjLuo6B2F/ZdOeU7o7iA2ac8LyYye6Ok3ZBso4gVWPnvwjJil
8kdkSGXwJRw+e5dtEIj9kA2jfgRJHDzbIdIRaMYJxLwor8Vqmjoefdxo7dMBF43L7LYbDWt3Vxcx
Z0UuEIQ9IbefcQJRQhS3a5nbPDKuL9HO1IbPbh2I2y3A4a41AAFjvfX+6oNJ0seY5JPl0/LGn6fO
A+d5CesLLM6guV9DQE8hVdATME1LjocD2swX3+lfHwdldM2R8ntpmevh824JCLIKIRL2QWKvUy9b
iSIpmofLwIFUufR5Qpln4PD8C9vuTanzkZ8WYYIOGMysoxmCuoi6DyWcZbyB8+eJqDW2yTwX8vCL
AvEd9i4D5fB4ajEf79x5GRWwkLoME/OW0tVRMDgJ12hUnOjRE9CoR8+BbX7n72BbsIbL7wCY2Zm7
3xzBT2wWQpxg7aT1UeAlTZjCERCoRFcGafh8ZBRs176BIo6sj5T1LIKP5wkzPTkBGY/crWULE7As
FBc+YeN36HoeD4HBxTu/DU1UfTJr/wDi/0xeiDKGXHPRBIQna6AQOKuDdTKXrtYDoSa54ELrp1pP
lk6knzstJak4B0bacbTEr3lyAuIPjDAn3kN+VmzKXRfy/xnP+4cS1m4k9NbWEunHgj9/GR/dgxqx
cIO6WQNCTMkAZHjvSkcs9nELq8T3sbnh7kDp1fSGt/rh0dKKIWJh1WXp8JBhjHDzviJdSQ9i0N18
AVdfl9sW6miE66BBW55oA81M0YAIcu5izsJZx1MAwTy7KfKUpuV9S7mdsIlSSKOq4Uxq4SV1T2EP
1ZrV+JC+QzX29I+4Q3Vvysyx5tAJjtJXyEHnOZFLSOM6c7ZWrV1mOasAq7OkpZA4Rhynegs2n8IA
6U+49kZoOZTvZQg+DguemPoJ620XSe/wb/OVR9nQgsBXkGxHPBbvcNIp/5J6okW6Oa6KYB7II4En
R9LiL2ctRjx5k/7pOQxdeUFT+kTH+G4qjC8w7LL2D7WIATqgU8qG+CSNyQI8Q6RpH6I4JEqtT6kt
+Iim+Fy+pMRc19MWQA3UJRjEnenE228QQBuVvZeMZ8Fr0U4HyKAZ1d4FT+RCFCMMkxWwny9N16LN
Zcn13vqtAVDT9OXo1kn4DX3n2+Euc2MGHeaaYCXup+hR3QEX2zIl/p0RJcPVB1xhtHeHjOXyoYH/
sUGd65idfV9YgWBt0PHPP0vNcvX08rQFLe8YYEwx0tyawGKdW8QSjMjUzIOEjA8LSifUp7E+MPKX
I8X3zdHFWjJMwwGb+GhZxl3oCjsL+2jrROe0jZ1eU86O55W7Z4svZVYCWkLLeMlbEbYhrL3guhyb
L2LAZMnmRx3pWe+GS/KPY68ArdKgU8dCdooMXOtw17VzDi8pXmEa7AB7vhpyNsyELpjFJZ2WR5Gl
++LTCbhuigqM0TLeB2jWsjVhgCmyEW6Gc7IncfPMfJpyaAIqsR3BTUgmIrdSjnMJ5GFYi/yoqzOi
mTzWTt8YIGvgkKsDKGtM4mphIYbnqzK2vGURsl59E+HwdGRkmMJ5fRCtpgYzSaYBobEAnJzjPdhz
tmwnJ1JM4MT6RMp56w8lYvhLyk6VrdrMybOUbiKYr5VHPn9ttCrJIlS76vbDXQ4xzlhYpWn3xGOw
7bKJLHaYt06mSSxnY6GMbbHJX4x9hjx+sDdQf9c0DcWfTSIuFyfxG+lbEvHuOGodOQ6JOl++HIPO
t3US0NKM+BDEAp+np3mqH6VilzFcPUCi54g/0v6edFwlM0OlJ9Ck4JAfSH/Ulaw75s6KO5gHTzwJ
GIt2hw65i5EP/3eIlBfh3xfA61pTndMjnrFDFBW3GXXnUGvWKtqbWgH2dhN5XGrjXKOMU3ZCXJfo
26HvOtkeMLkwaiBtRJqCU68wryBPsb5Fsd4XeXVu9f50yubn5IVW4fHEcA21EQaw4rz9sS/nJwAP
yrxbg6YIGti+Mx8yQGzby5OEKm+eEJ3fTjgAUkvGybclmQsWAXMHpvIV5t8s0Sq4kVkiLpogvrPQ
j+N754aMCGM2c1Oo9xZYKujgItMhCPsvRi0uFMKCHIsT+pUp76vlW8Q18Ws0Vm57/nLA4PDNY4PU
hP/9I1Gt2nrBtU+lKHYX4UCQrnI6VucoPv3Wz/Vq1gQSlhJmjhDnJTDfEfwrelK5aGFinec5qbQ9
OaC3KxByFxQGjIiNyuo4YEcoDhZH2xGykp0uz/HLZY437RSU8ejJMJOw6Ezw0ebUS6ys3chJIqrk
UAmnX70Jl5DsUSiccrQcbv+fMvPJBvddjgTKLrLkf78jEy5idCWGYOw8B0e2ui7YKUKDATXEZglw
FXXdRRrgC2MJpfI/NKRApvk+alXyQbs/guVDMWZVDtGkww/WH8hhp1l0/EUKsOhGND/9jkFXvKTv
pUXUv5G/cDKSYeBHupj/hMRdiv4UU1r//jvtTfjISWliQzIlvURBImaJc1YLbO65jjZYedAnY9G7
c5nIAczOHq4lky8459Zry7jmtzdCg5eKt3zERkturxx7wsqxDKsenj1q3gCW+Eodzjusiw3liSGd
gx6HwLnYpxv5PlNpz2Q1qgt2EZ1ibLf7uA/pMG3FTq6mXTwGYYzaY0nrIaLp769K/FxXLjWl49vw
VNU3sSyxBNTJBuBPw8zfinHLkS1GXkL8nlx4t1vnxidtcO+7HLmsXUQKOXDgyOfLf9x+CLx+7+VT
JSB24eGKIXlyphAqF5+9NlfDTmxqhiYeQG7XXvY3Hic5Cd1urhZQ9m/Rkd7z5p3ZKX0YVnOG4DKg
2Wjg9CwfOtZTRilWXdKsLlJWJtFjUJuxblN+sKBvORlDXn18NL4gJWUnYu5WMCvNWzT4DqF8J0Sp
q+prc9C6F0f37gk5Jo5QwQ43OKkClP4XdoeJa5cwbwG2oDQDb5Mzh6HToy8LGuMp67wpqDkFIO97
0+3zv/CZmM/uwHtU41LyFiH7fZrawtPYqXNzJnjshREgH6L+XqXQ7DNAbT5XeE2g3ESvRWMn0lqd
zQuoZTwZaL5ajokTW+r3WbfCYLoGxQiZiD3zppiYkB/l0k6YAZNDIC6um7sj275+dxI7mRvF7+68
s6laLROQWRqSbPZ3wmsfSG9bQAxl9X2qh2wy+bNBMDRwUbOY15JEGz4elKrtF7OqsA5B7zBSstME
om97VMDxxZLPEh1Oj1qwrPVMpiXo10IcXobylp0cS2hxfjyoW/+OR5DS1HyAKJqVcTIgLXm0wrCt
PW0MZEJ8ZE3vZ+LSm8Lx6kHMHP7JOabwOnZhPryB+EOhtIyD5f9j3RIuMt3qu2H14HbcskPcGZVm
rr79EpvxH+rz+qOH6ZJsDjOMwW0aOg+yK9b/HymdPzMt1wXPelXkWBrxqRcBKf50MzEtUuREOKA9
LWjjxcHxA9nVvF9Hhp14zVA90SdEi/xnt25D6CWJ3qnARSoXkRrsuybolMRo59fASCauPVkR9uPW
Mpy7JXl+l7GKJpficPZbfxR374xcE94y8M9EK/XYJV6zvs/kHTQ8c3xJvyqFvNvJZYmttmJSEu5o
IpqpYAjnIpxTdcEFX9WCjnOnPK95WV304iRR/+ZUwuivE4Lt8n+qPhVjyVS0TM9eZBkpYnddvSwk
gJmLZ8TQyBxJ1HGc6ECm+9+6Nh+dDsxj3rP4Mzzjl0abP+4LylYkHAEHW/emB9Mp0HfG2F2Pfe1a
ULzhG1NfZTUXetpU0su0cfEWyFaX4Ri8fDoRkSAidg6cvBtIS0tIpUS4vlEsPzqtjhaHmQT/E+Sd
olC3qNXyNQmB+zNONiJdYczFqb/BuMRyRYceAgs1tUKssiJgLFpeafoWHgPdxYGBaMrFGL5eo+/2
DiLxPnXRX5ll+CdTnhnE6yNHsCaTeUm3wUzhg+dpe8sYVfbsHJDjNqQ25/4UJgW8N0Jh7cmjiwzT
ZvWd0aKkpyxsVoG7Q+R7C2PMLSMWmr3V5M7p4z99k/YWu73ynA5P4lw8KQz0qRZ3TT4Z/JwRqWaY
GyanwwcGc0hignwF+qVJnbBr/QPvT8LRSdMjViLNyCIUpn1sfUGpS6C3weT2EJC4BP7V0s7ICM0u
7ifCqVMICwO+/UZD0yOwOiGIOprDgrvY3Q1THFAdUhhFEw+b0PC585ArvqWvDSMEYvlybywV95wT
K5A0VHO56np0ctvYwGqas5DDAR/QaqnvVGGd924UoEoX/sgHi8/8G2QXgBeDFyLo1aR9RNTpdiQq
MEXMEwWVIJEc0TFnZPPwPjNFNXhykPM7bWNKlHMY9E2wCmKwEg7Mgc2IQFZo/KiITNmqnnSpcQhV
eZvqH3BXK+IFmPkxlPwHMVDcgl9XXHx+zm0NgaEedQcZvFIRs31ZyLTCkN2yU9SDWHc6I/DTJPz4
ixdit46XBMeeTEmjkyID650t8g1SgxSeNb55xCs2FWgEWMisovZTSubKHQ/ecff4cJF8G/QnCg57
JlqoLRAMybkeLP3PcnY2F0NHETpVson0hT36BDVSDODCzHyz0TBP5g4zvpj9HwynYfitz+CWatV0
znBt49pyTduY5evce/P070klxB2SRdbi2Xf2Sfu55mZNy5Ct6OBT4eunzFOwpfuhKa0J51+8n0sI
6pcPN60ehMy0znovqiG9itQfWIuq21sAuNT7mDYHjvizHmc3btETA1gobjKcFfqnLn4z3YD8djNa
vdlnEMXnR//oHTB0wZGKXbY/UljVE/F2cZ0zBVTGNK4adFHuPB5O1r9u9KP1ne+vb9ExAbFT/de2
51eMhV6ftdmlTKPxa7Rw4C9QBTGWDNt+0dn6Op08Vqdwes3mi0RZSxhfFeT6WDCftfxKyj2liW+N
it4YhLaIX+sritZ34S/+Icb1YSpaM0Imh0m2V/o5Cord3fFbhcV6h8RjbNVQY7zsklGex6C7hYMB
frxUXq/YFy6Yp2uvQETVoC1gQVlkN3Ur0EKHEv3cq5ho6t3k311PAaT6J0YMc34s9NtpSbNVR/MP
kQqL+iOaKJ3zL+PxxE9A2A5rLPRebXFd80NT1PWMyMTw7T1Z5G7539UBiY5BRSIAT1C98fR6iPnE
n+UDzlaWLvjUMS5SnWiXnayJAKacG2qblpaLc0EZE3ZXCfwsyay4Ly4UaU3S5203kuxAhLcy0OeE
gYfR6gvU3g8hLUx/Ab7e1YbGY85a89dRC1tFZoc7dY63qFfybTSjFisHfGE+BjpsSFqJA3HvuJZA
uvNE71EsFJyPZmW18XZRkMlDcsnm/Cpdn3xUkkAfL/0dnFSiG2E1Fu7T6geC5mjuX/Ge8UWVQers
leqni52ZvzMGEjBm70U80/SQiA0nrFTjwNilR/AnUY91tu0v9TTuQZE+wMB7wGuv6gR6arj9qvV1
SUHNYo1/+9mA8PQArv8I2Hjw04AF0evJ2EJk/ppydhyoAotR1C2KaiQfNH7F2kCNAADonHjNU2+3
4tTEbOXdQaZKIXFyTrqZrsmR/GDka0bMEh+ly+XO/h9anMIrSjFoqH/jzucFRSBSyzSSLEi2hv4/
QlSB3oIN70ChSz7lvKTSvjtkEq9CSiglSZxpOLWOQsdNE7wFpDCNkD9nzS0PzTajE2ebW/8lO9+O
ZwWlc57lZOQ9fA/gWIuHrt+2XMUA0auEFSa8Jnegpc1RLn0JIAt39vk5jWXGzjm5qk+KxcoxKl4+
oSQrVJrmUN2fswNiUFFFtBCZ/OClhvo/VHWJivU3EzuIwkeYNWDljOVUGfgcHw4UlUddy474NnxJ
SAANk/YP3dFNhh3HucNJ7AKDdWg89UFl5fybDghlCMPruOHJt2zhFMPNZYqNyM15qG9q83caJAEY
m87kOp6il0PKsiPoUwsvhoG0dOt6CA4WL12aUNIDCznzWulKgEW3mpdFKKNifjrrhq0pdIXI4BqO
ae03Qo9iqfI68Mjy/m442gvG2+tkYNclHNKM5HJ5CXY2TH7bUzM5GZY19u4umXaN2DwYNJk1YULj
dxwmzRcwSZUg4TxxY3ZHUyouVvElSxKESK2c9Mryx2O1tA5yL/hC5oVXFLrDcmXKDhRw+HIvNqL8
upuP4rHwb4ML44b+2yyWfif2gBag7QSg2LMULQqkBrAZWI6zmClYpvzXnov8f/wX7wMM+bFILXTD
TGRw/EuN7zYCNxWUIwxU46stRHPntSpdTvfexAqEIPLV4G35vhRGQVibu2N06MqK1zHRqvxcj/2K
QaKXw/LvsgXM+OyMo/4ehB+xnnHAfAXCfXjPx4TFmSDhWOsIRW6CoKUhAgiZtNmDiH922IpfKsJ7
6WjqI8igD7tYxBGvKxS16FXB21WJn0p2rEJuL/fwWjVvBV6zicx5udr9bpzmrpa4w4A7xvk3qaV3
Y4JaDhryOCOAfYS/RDGsWTMiXlu3dIvFEORjCERetQr1ZooPVh0ePLDZJuYe+5Zv1LZEL8GycuIX
qlEIgnQHhGGz2lqjfy3JaXTwmG/c4mExM+85VKrex8HcV3RU4WXrCw3aoc4xzSnVKpQ6Dv+sa1wY
0qw1aCiMpW7u3T0fk+ZXMISkbcWtlWnyQMzSYKR00sdP7ImBZFUjy56un3hzFkcL1i22ZlqthUMx
1Wkqbtzw/mi+n3FpLC9g1Pql1HcKNFw6MXerddU5Ev8ljPXX6aQTI4Dy/GE0fiXPNRhI8N0sPDq4
zbE0YZiF+EZFsb0ZPkFZYtJDX0gQCDYh9fquW9uE0APAMltroYwovwzxkikOx8YZymuo7TGMYXSN
VDf+2CF5IqhfmOiITUZukMhoax5Jl1yJtC1mbbgHuzfSHDCqvngzfUoZTtZt7EZCS6zjKRKlbuqL
oq/yfwl7maITbTjmsksyPIWGac7LhDt2RrROxzSPZQmDkKQXQxOVk8hVvLln9OlyxH2yDju/xhxP
Op2npuVwHW7AJNXDZL7sAfGgpLft3cGOQTe/fKJuYF9PC1KUylP9fea445J0TC3Jhag/y8tNkccz
ratEGptXAW8lW3jhEhg63/Ny4WBoGatJGwCZ4ikgkVRqgxGwwWXuC3wAJWyje8JznnV5Eb/Qca4z
8UsPxGHlEFjDcPBf0Jig059PFvMwRTHMRWIhjdMrlLqZDsdOJ4u8Za+K5OlrzWPAfJLBARu73CDG
U3gQDpW1/z2+ZXaWk94N3aB0W0AR0peOHvsJzaVIMtOgsRwgfIcKZvUDrcuUVEhrLF1Y1vMnS8QG
FaAMLLHp3uxecc0HT0zmXrQqqZkTD3jPSsYlTXMkI0FABobGvVeeMQWa/dumN478sTpbFE2sIz28
sy1nFDi2AEvPAXbmZBcbNZtMJKartwiP5ktSfa0tRcK2SkBrAtkM1XhxlR/llAvQ0rN7m2mc4bmq
jwSmb8t07iXkIITlW8dG3w+Yj5AccrGd8vM3HVmB4zBDb856BWADESJQbG2Xem6WWn44VTjclRHT
4IN2o7XF+ld/ohOhzL7l/BqrcoKQFIrkZVc1M3iMd2q8wDmL6sioz0SDl3bgc+kbNWkzIviLts59
c1xx7SzulR/0F1/O1G68aKSU9jNmBcB/32Z8YW/+4jmAT3rwvETrcZQ4C09NNmxOKxBuVpQffvAC
dd9B7+rOvspeFL7vXvGK65HSwS/X7OBiMUM/wYkdImwPcS2ksJQZ8xjlWgahr+JPukXdqQt2E+Fy
bjBtVBMm453KmSY4EDQxHQytpJRCNGTokyBLWhKKfX3QZsjBXsiEtQw41sSigT5ockVn/g8g4nJ/
iAIjsD+MM8H16PcncdASU6fGUUu9cEUP+yG1U44RGcRq1MNMzoZ44xJqvPJSuku67nOKym6w7iMV
yO+JwE1lWCdSoR/TCe2RR9JLlO/dTPr//ZipZkgFE5QWsgYcGdAWIFK+GcFicA6xmCh67Cba04oF
ctPWxr8kaZIRbyS4+igVqEc4I++zb7BXi1HTH4EGbE7wRfSRcANChJmbDayzQpUnC5jt3kaS4tBr
AY0cI+6Y7Iw+mBqv3vdRp7YyGHTwSW5B/u3gOAzGUOhDEKpfJCR3cvtR5FqFehlPvJDr1ysDf8ow
c1YFbj6T3B+kOClvVHSyFeDi5eVxuIS6rfriGwxtpVzWF1V7Y58X6DHNbZkoYWeWOQcztE5y777V
0q2zDuIK3rAnMaZCVUf2nbV7U7ZFqTtV2JIhv3GjNUUTTgemXMSfWIl1PGinL7EX/crfzXTivGpm
Cv8iWlPkDKrg3mycFZyhMp7wt52a8VfA5yNr7HvGVmNtCN8IhCZsUdYcalrbKGWicWP5dKZzG0a+
bAe+tlfy0i5tIFHGdcrItjXy1nRC15Ld1Eyye3tCCUVFt7Uf55bKshThck0uoCmuR/8pALovlVDX
F2UtWUsZTYk4vR9daykSh7B8M+Eo8dXheYWeJ2KUnU1U396yi0UcfToSYcz+g5CshAcE1nYmz/Rg
hfDCeSThzlwz94bcE369Ik1s9nQVIrYUKMqfNbvpwll87V1kD6FIThFcu9+ylRQ1h3vmei4Z/6bC
Jto3SzGYLUhjyg3DAP9dfhuITEZcynshL1nx8CWNHdEWWuiPc0ENiZM6/sVaxv3f85Mcf3kZ8NB7
uiVdbWco/kiH3P+BvtGubCXV0mnAZU+A0B02auZC8xfRPAJPAunz5EG3BvtnwjSxcJXJt8tT1sfn
d0EjpTITnNjLsR5vXO9XoUS91KS00dq9uOSGVJydvyaOHwRl5kp21+gtYcOO/ZjDDZw1kGSTTX5T
Tl9b9lF5b7KokNwe7ASl15+pm7+DfqRiINh0g923XkV/IkA3J8doIa+Qlwqr3WcL3nEs9zGr/R5k
x+hwLPsfQ6AP1O3M80HWzVfL17gUNDSitc0iFrTkcoU3kcDV48rEw/an89iQZqu/4yr4ZQvRmhoM
kisKCNeeS04XOApgIAQ8CFDWi3HOSRZyHKogrY2gem5boc/m7Hwz+I5v7HO1PnG/9fF7pRo9Vggr
mhEjgtWv255G4Pv7aQ5CWyq9QcGCJ9PWbtxVphDJthYG6KZvDNAL5jTz9i0SikoCwa9Q0SM4/mrV
XRa3yIqVjHdyJlEAYxiIiMFdJXTNbzMpK6VaDi4v3I91DD7VGOlj3n2g1ko8+7qThhCfcEYrhVjh
iGuNYFrR+exSfh56930edpbhCKficfy14Vp0al4DUGAxOD0laACAm40JC5agwRz1dVShH4QFdfTs
CkA2t2O/cCwCR5FEZ6TT773jBcKbGbInz7tFPi3TL8gGQTPG1QQL5MfoDCmXhylgK3uogX9/nD7R
6nAo2wWsngxQTMsDhLhcjh32yKkk8gc62M/9Hm77NBoWyFrkGSi5siqzrU6c4CD0MmC0JbEYS7tV
5iL+ayYh4aU64c2H+pu6HHgqeSrhOqMPShuMoRCymXAw0DGJb0X7HP9Y5w8dSskfbCECV4xzfP3z
EWpjJcIRKQBcXbQUubZNNavj1sr8cT0Od5BWx6t2fDX7B52n+DagzDHO2p0M695jtRZAEjozoHLl
Cz/IC2opYVSePLOlC26CTOT+FdHPq5JG0G1mIocG7GxmWSH0Gmqa/Dhanumq7ZhItNsFHmhv91RN
knMa7osvB0H53tZiw3wXC4etCUbJ/p1Z2Qymez6o0nyGJaK1zFfY/7Wm29bCF1iLDgxlIdY+3MH6
YaRcR95sQWLtN6WOz5rm8U/Q7iU/yjK2BB23HOAWLYnmxAJNVXgVhfjENIBl+gI4SVhubFrZLB98
0nIqeXuORaqv4stq8muEAE+70hS2QYrIqXflTdCk2QUCbg4s+s3lBSzuy0EbkmyRBF5r+34IMxBT
wrAQXZGqF6ojJ77YoQOr1H3Pw6qCbaN4Mp3GqMGAl8y51XqSb6t4uE/z5kzB1gizxHZKGE8LQ1IZ
W3Tzj4Do0ppJfmHOWKIzxQIS+bS7VgaKJORQFSqKgaSa2fhC7YBt0ElHA5qY+/68ubuZkmlyVCsu
V4rdlZw+IJEEldYgHP/27KK0oH6R/+oxuGP7dupBx+ROQthRD9+5hamRB/+xEdwyCJWG9kFDSDTg
oeVh0ck7LKrAJi0V0LBFXXqJMkHPN4g4uBBByP8RNg+URCvwfcT6FX4EnFaqZka53Z6gruCHMK+7
0R8oi96c96U1xBen5sUcy3bbRY686nGnTHmsJaGECBUjFIogevgfmrLsO1NKIA6aLvDSMl1Htz1V
++BH3Vy2eyhITCbBwedB4IjniQOqLPTUX8OvSWAblzSOre/C0LYQJ3qbNtNJs/BAeN/EBi8uFe0x
mb17GNCmvUyD8vQcHxbGUXQmcD06obM+yC2yfP1ku31kM4AMUhcLYRTt7ch/e/q1UZctOhKp2qlA
ZnCmYK04JBZ3xGkqCl4HcHxaPqN9hSYu7+A4GCsZKC2z/Oof3AptEO8tiD+S90DmCm6rEP559/nW
vDcVG/NLVPIoo0NQvv9Qn/EpH1aDULS5y3HDJ0oRDgd5w9t2fjIyqPcn3IQCx0KypVcJP7qEmBZO
aUT+6qyfgBGsfzE5rVLAqHPw2A88X9WaO9rzZ0VslmYtUIzd3n1XP2IeM2ObFWMnipZoxgtTWWOl
0IxzQnUEvofEbBGYblgFIoi1US3tbh8Xhtt+Gr/7OVqZc0reg56UijOn5GG1lTgR4IUCLtOq/nU5
yEe90RBZ68qiUju7L+jhybopVAe9Lx41I5l6uWnTGYwyAqnjkVRrD56j9Fm6UwAtWHsWiA0MhuFV
G6sudl8pIPMiYeSrb9uL/EDYNxNX22b2/o2NUOXJ+oHM8XNgb0OHziXlA4Mg8ktrpyO4lo9wq6pQ
7wEGMovjyGhMxZML3srnv9hn1QgCbfb/RCjheeXQogkmpw3XVTtCiyq0EJitjyT86loo5O5hgLIE
ImAQQOkUckwXLYTJkXPwZ7zSUjsW7Wq+JiiWtxmyWsuzNQSaZcoLMlA8WBmgrS2k5n0O3DPNCtY2
+RpCStUChuD+MsRTVhpQmQQSrumGMRqzCyuiSXzay5XPq43xISGpngnA+PahqYTruSj2EV/gE/UG
mDP1NS1JY/OC3P7c4XsPZPvsKppZDQp5ocOEFjpl4q+ZlWnmiFDUm6xYv93TlswV/HF4Mrcyk0LD
AjaikzCVEIE+RNDCpnxB3qAlAbIu6Ikfzykp/h7QlewIqN644Llcs4MNdPwCXvlu1WggOUinXthX
5X/4MLlKEgE0EYbkGCSIKYJIFby5nwaPw1hn7JDqdgRpsaHlsPbwbLhcZkQgAe2LmNOAnYNfvBB9
A36/wYyltgrQaN19A3aCMOXSLhTFtAMj8FNJg3Aur6hUePDeyqpIDh7RhRnX2cuD1nPcZQSDoMem
dUEzHHeHAQkV3Wh+Gpjt0ctV9hpO2vseUilEdY87Z5r+kmrWE1NH5auJGHd4+RHAP7DPxP/lf9xC
6Fofg81zWxmn/MZx9v8OujHVYp6Udrx+W6CmAYyYcdiph4SiAM7BhBJjJy6ykwSXPh4U52jqWC/j
tQzp10LmsnOG0C5++Myc/Sz32g/qds0Ew/J0wLo08oUKn2qTUIJ8JF/7jy1Oa4XhNlxXMiv4Tzni
TU4/AX+8PKtxhIIll7luWh8sfPe6DLBNmrFPW8OcpZLanFxhXTcOu1fmONNKSsT7nVsc4ccHd+4l
vlkINVewl+0krh6lmzdWHu8HtAerhI1k6Zepj5Q3FKjHNviC2m2Mre7Op4vk36Z7SPX/K9Iw/zz/
z6v5dAxZ2CgV5xTn9OScAsHMSm0eH38sfJP0s/ynLPgYCG7RRizhSUjXr+G9F0SWyucnLFv4pp1w
CR/QEMk7t4FE3T/BQgYmo2eN7cvxi1OZXOGgYe6foPMR7t6C1mbrxDgxT9UWWikFpiJev7q5/No3
zMaaVSVZa9CXq3ey9NOKBwf8MEi3kYynrAe5PIxvS+w/O7XgkLNLoJWtXtyG9MVAmYzN0KW8FLWP
tFgMfU2ybK+OdCXITJPWyfVqh0fQ0dEH0uYrmAZ0Z/mq/fhYHAomYz7Jwddeo/xwxt0PGyZlHuvn
/cf1VW3QLgzX1hD9vA+MGz7tl9gP+/6+PbgYK6QbN7M0Xp1kobt5verx0BsvBgJTNgwtUMIOdVvL
HCZ3vXecP4AbyqOneKxK+bwRN+GX2ViLPNAP0cuRNe1DH0bwrmyVjDpsNvvzDxVOPTAMo7/3QZac
5UrrUnrn4dn/c6omzkfJR01uBB2Y0WJ0KnVVrhLb4JpqkNcRtwRSdWSI9DcPugK027Etxjn82Rfi
pGnyj6X/tOMTOwWtmCu/OS7FJ6a9xPaIdPGB1zGbhQqbiKdBkmk0YBFZFnCos2XgZ5SvNsOpCuGE
tsp9aOd8fs1hpHdllWdGmjFNVAQZE5l3TUNgkTbP3msECkN345iJhptPbF0TrQPoUnHwvDgO7436
Y+z2KQQT59Hi2uEjLo+G9ay0FmZY14qcA5UvtamtIcT0jtN6cJNNEHGmMtOEuNNVxm2Sk+lrZTHL
H8K4RbBc8ksZFWKx7N+Q64WlJEOTnpJCwHb4IaXO1tmfsjwEJPrXssGMJbmQHeB0thAp9yLf9apg
n2WLoLXp0tHKmthR8kb/uMiYdnT2loH3ZV0//unPfGYDbQv82X6V+3YfvWjmXfA+BbAw2/0J8f1W
EkYwtcTnGtob3JKHqlceO7IrxCs7DegbPS+p8/zfKIDfFPF593+SDh4k9M6/8ze6su4CoEG2kj2h
scXsQAQQnUIPgKPJwo/n+wBJoSsCLUjHR0puzOZw4hLo2trAHsNeXcCYDdGgHA7buwa+hFgOCh5b
5Ri5c3Rpr08FEnZC61fspQyK9sMLWKPKXX12BXqvXGzkmbIfkVqlLvsMPAkdyRK0QMr6we3nppe6
7cF6eAgH4LRUAyygn6EiGvOiNuP9sOFmqfFsl5K6p4Q63yL7+/hrEVPinM79mRfX11r3OiO0mdiS
4/PhYhKvcgfyLJqn6GG381RZWgOpkbOE6HlyGvbpHjm2j3p+xwjtRy17CKi9QcJQw5XBYloYvO2o
aizTBe5vFmKNSpegRF5uCUmIEwn0aJhMIjaJxVc2DP5df8AEUMg6lXctN7JXUYck048T2G9iBMT6
1QWFDQN9Z3UjCt7v0IcVtD1t5ifI4W81ZVGQ4RKQW668an2pqzouInU5N2zMzpuhCXCu7mvm+sK9
jr51kaJBF800Zowiwy84SOEnIN3vxDfmTmrGL4DMWxYt6tBOigOGK+rtChT1XOE7o1NyHo+6bwDV
3seBa6d9bpz+1Qa08Ruhpfnn8xDNY16RW2PTGC6SvSccAYwYy1iyZsYMLtRXAoqvgUWWAQmwH3SN
tBDYykFssPiLk30lzXSSCGHN9nYY7h4ccMJY+ndD1eujTj5w//+VIlHBoGGP0wvm8oRLSzdQDVDH
oWw5/jO/TcjcdV4pj8sJnOaqmWJLMBcpd7Mgzb1lPOvUVJGnVqgRhwLHit4ZI3I3LCFjpEcTL1RG
lW8aKhLXz7HSo1oCEWB8ulD80bUqNS8aYMqsAhP9YHpMfWByeml0nwUvGouuvc6jU4kx/goOclcG
ske64BsFNyrd35P8QrqmNeyjFpi4j8OhZmRdsJqjQ/Wd1eaiOyHfCzcLAKGfd4qtcLDK2vDRWwR/
jzPb70XdX10ONB/4ER9NIsDxYfAwwap43BWhMCmZK1lbV7h0oIHxfSq04HCIrGjYuQyM8+Mq4JGl
844T+2SZ0vdb6AO/dhQ57OWRWc0x0rFTsNnH5TevYIeioJQmBl/8CHVKE0iBA0fo5LaWiV22tdfS
4L/wRJsNP6PW/s64NuSi8KpcwJ3+DWdt2m0ag46+GjRm/rfljRcK510jfbAW6EBNNlN8OF4Q2Fy/
4YEzFr41GF12ITq9ZF6Er18ZzhMiJqIoxIs9gUR/rYz9nGQcF4LCDDfkPa4aKlY91BT9ygKpo2Yw
03KMaSp0+OGedsx1qh5CTbZl21EXRCOjc/4ibkmXJHY/W9KxtRmagDJkKvC0JODTncF16azVl2X2
weraCvD8kE/397EIf6KepMPVc+ncHFyT8QYBcl6Dptv7Va6G8m1DMEO9H3RgvGTSWQ9xYYx5jm1h
0cqm4PSSiVaYxIY/K9w8IqAjDLxSyjaFaKoWQDv1O1zh+Gz+vWk0hJYTAgMUSSVnJPTUprWHNLlS
Q1qc6h9/rqWPUqAmjh3vkGo6lXFCDkr4eXfAaJqYGiaME281WfYsp5gM8idUuAA93oXR2IUYZcDJ
Le7aXElLnLGXyESu95UQ+BtPv1rbo+ZGuFB/lzlaudyvNCghpSLmBVensKFnkmOkZQCfTl0jlzkn
Zr4oi20o+35ZuRRAGk4Cwvst2lPu32iEAEQMvD4qBgc9mElPWew5yoQxo4NrUpSAyEij0EplVd2s
w/1C3XptJfcLXDGG5boEqlZLo8ZPWQyBLqwdAY63G0dTsQp+GCqgCwS+8X9Jm0BtrHrQR+UkvAeX
aPKiNdaY1tnQpzQ3r0+uzynjHa7twO3UnLLBvHTQUddIxLqd5h1cVLz5m5A2U/tYFtq8S67u6uXt
BW9In50CP3B8Jm9RQ9i5J/J2wR/huSKtRBpXt8djw+NXX1UO98LmCLJWsRlyjczmxgpzTRdRxDkZ
m1AstkWjdKr6RZ4kinpwL1uvF9qF4RixGRUJbHiK5SBGOGjNhS3avNz5CQPeC2ox2liJeGjEp/Uz
d7xfzRsWCcYnn4TmESF4QRlwRrCaWiMJLF1UB7Piqu69SC4LrJNUrSy+CdcyNi6LjJRzHHnN7ApY
29X3YHjeaqOgzZDLf9J134zxin9aXvUiRBp4OYhmC9xKdsSHwt2/B317r4udQVXTm7V1EBZSrBAj
WQPZH1cl6rPMFGLfy+7h58HPl3UDxYp+awqJOOwpAxFpEURQeS93yhG0gQq9VJYdim1E39BulU+6
feTAML2Spu9F8sRmoDlJmb3j/gcUlNnLwoZBOkzwokmRozntpfsbcPXZduUahw/rauvnPW7JBu/6
x3wpj+K6+Vwf8hC4J6J++Z8Poz/mhZDXuyKMbSaU2vOMQxZVZggTrEGvdhiA/Z5/c3BY3xy4y/0T
x2i8qY8bwQxcs8hXgN83mPqyj191cm58LLYtKEey/g4HmgOJs9qLOTJHBlnGDoRlGBrWpLpn+6Oe
xm00NqEic6nRw8hMsATux7gjU2gtG20WOYZ/8NLOD3dDiE0vWGT6IUqayg42qJwWL/06IMzOvosP
RZy6N3juuwg8+I1szavavIkh8yHFulT4Z54Zar8gW6TKEYcd4qZXwEmQQ0Sz2eyUh+4XTC6E2SoR
QYb4HvpknUzMIhHfOLJaQmYwjini4C3VoFxQP06hqHyk063Zb5nmGOUzn8Hzrh25GxdvOYyGmgrC
GFwersBYU+tauU+zy2Qx1RYI8Ykwx4dEwV2dkdzVkX3L7B4BboqXEagzao6gnai5ujkeO9W6DOPN
seJevnLrk2INs0UMemDcuClDMA18LAeyl9E6JGW7HTV1iXUHp+X04+DVUKY2pHTieFGvmhFD7YVD
FPsnrJccAnmQE6tiXS0g5P0JgKs5XRw5o91GFlFgHgul20HXeRFh0z7zQo89+4Zzf6PGubrtJbrT
RapWQYJ1BNtNKMjLl0mpN8hntJ85Mi+eyDl2TuHR5q/Icj5a/flTncb+HG36L7PDtRuFQlV7zg0/
KRebSwlhXLrLow5fAek9t2GnlEC2KQD1fb6PjjiCNoj1QCwuWOrIHX4JlyLlJQ1JhDZaOZMHZaXK
84uXZDzWH/86G4RICDyxQg3Osxai5FpF9opXFp1FIldbiHUmnRpZOF3bBMUxozTCo95BL5nd9i+U
iXwIGsQF0fNQDy5630yEMuF7MOsu8g7iUPhAKkNR5QIDuI/0gLKZt15p5GIpo/Mwi0GgW6nWio1b
7vons0VnQS6K8af37i2G1UT4sCAjirqBLDfC+nfAf9XWBYnjvyITNN2EP5XBYcZUp+9mZKRz3USw
epsywHyI9rQnbMLWgM/j7EOTpBqQ1Q4SgC90mtCPLcqc6UoapAG7rVfZWkwZLE5ZRyZJzacwc9zN
nUe5Z0NYsdLr7GATTlJUY2Sx25fvUTf0DdESFhnRGl2HuV//AEv7t3Y8b+9FoQ5MJqDU1UTkvHMZ
q30y+Aylrp5h+5xkkharNOdMQ1SyWVnTuruqsHAFKxADTU2MTAaxDM+bXOqgk8UFr6wtsEjo99D6
LF2QDf2F5muanmeAFvVU/Hf1xkZCsqsRHq4u6NaGwwEf+jFBMJHrhoLBvjCZf5ZSBUDTdeW3xuX3
MHz78Vtet03baRuIz1Me4W0RV28FxHeZfG+1rnAf9RL8L6tb/Eo0N2HyODUbD/F1xyEvoU4xuDuD
rBEbJQz9maEtHen1sVXyQTTApsTqpK+AWZsZseI7weTU8Vpa6iRfE+YHWz+NBrzIYVcHAgThcUPO
esWKE7+uUUJt8G/dDYhlSSiITYrZeroyTE/pte5KSzjaYc/AEKfW5ulC+OqMT7f/gPVr7L1rnvZP
iZr4UynM+dC+z8tgiLk4JlSuyhEW/hBxyaGks5tFDf5/Sd5mOR/CsMGIDeTN0NrvQwdxbMywQ97u
7qUL6qP5fG2Cew33+ifuPA3MBC7ZK86NF5aapxVvhzQ6tbR5cS2lMGQ44QgtqApUlMzf+60gCoWH
ceAm8NETyCrTiF1d7kUrIMNQOfs6g75E6tUK9EO6tTPAm4yjbPc247qJsV/kpMRtnxWC9/A5tGvs
7Mok7uLNqZDKUP4fIWOqKpg0z6yPTOdj2TH5b9RHIybypuWE+2vd96eDth4yLPncJNkV90V3c4JK
rk11RD7ugcrJsBhtTA5AhLFfqEH8ZxhApUqF/sJpjKAyfxtIPSVnmXZJxwp08AMlCVyHFHYkTjZS
4X6dJxuCodjs0sxBfbX1eGqCtQ4m0fuh2xKRNGrUDDWtWsEnn95ir69WgHM2bvAMWFx5oxW5Tn02
3WL/wABZe9rxwN8Oq3i6Qs5lPX8vDmbRCrcK+eiiCloYdBVvMHcEkhFpIa/0zc/Q+GOBdrypXArV
Cn9fs9uSzYtWyuR5A91B8Y11qb7vSkt/HF347yrtmt+eP+Cb7DYDuRQ0czFxpzUVJkVb3nVpmlf5
wVw45M4n0V9Krvpe1OiF8hghMLjo3vpUhIAh95GwO4lxaOKtqjbCjFhaiDuPmw7zmGTDJQSnryZy
9UfdGBRcap0JmIYh+tXavpWGu9dWSsfLnGa7cYP8Zmwfl72F1Rsgxh8UZc9rjxBhg+we4MNQ7Dka
tqeyqtNIwbde3o3JnRYZkUkoR5v3KI7F6RjNALWE8T1K44juAUtMbXV3T6oEHnZpGRez0suKoUM7
/rHvfv6Pa0fTPf0DGdzl1JYkgm8PZSLUycAWjdV+/mGkrQOgmXdz2lwsXXw/wE4w9aYsLykDJvcS
5bScrQINwKEOOOnECYi4AteVyiYQKgHelXZqQ1gSmaGvH5uGr7yUZkjuQ/Tth2N5JCxvqyNhP4xG
S5OBZt9nimK7sSrJifWXrId/86vhtrTBqFuOfUTQBRApiUUzTJ1hVfTOLWw5mCU3D2a/OeRKyctX
rbA26ncg7cSWy2QeV4FSmrWVKlxz8oBiiLopybk8JUYGoebUhmdwazb04Biibf/nQazXqDdqfa2H
+kD44bS15YSWhSEhdOE7b9B4rsl56J/NjvdXrzpwomezjOGGuMQaROUhKbXjCF78IY8r8DnsWC0N
TF+XlWMs+s9nkVCrYvwK1UxDIqcaYxBJ5sgGW3djy8YHD0kGxYfdPZHGXu3J6chzdha5ck8foIPC
n4cUj7A7d4HUhHbSbs74A4DEQyEi6/EWwySY2I+QnaANXFcdSO5XrMbFqAmsdnGh+rXRTnvIuVWo
bkW5TlDayFte8ry38vRxNFfzURjiTxwLgv6rty+VKm6ZXmPz90nEYqAA5YL1C6W/bZkipudBJgZC
JWvJdQvwhj8zT6aIiAOTM+CXgglsLWxUkLdgxSPjtUb0zOrsSWxXbpVxi9MLnDzXdu4CYHF10BHW
juoxg0vd43XUSHFgQRGpDfwyInlnlumTNl7WaaJanW7h2+3vPBuC7F7YL/FmMmok/MhAJnH8X2v2
EWGeRAXCEWz4W4XoJpFN9gTpDXF59/X+SQhuZl58WiPwYv06HshsiWmdvuzd/+drru6F2WFQ4FNF
zrTK/kOem9W6xcN6I2+zTt0PWtrU0/y9Me4xTWs+eYMCPm1IwED5V7DzZaipeF9RGPYHaooSE96A
l32aNHFsktdM9T2+jo/jO2NxZ6U1N7dZbwq0a+bg/4FTZVwjqa4ZWczQBXLtY12IjQydmfmlCbjN
SkNpkIABiTZ3mBLYVCI/l1DPkrOejpleM8twNpNuNu3scRNzBV9TnyY7tAz8cbw77+5ynnSTSz7U
vPo0qbY3hm6ELAyGd8/tYArnejNdWQYc9FqsB1HrScm6aJoW1i1RlZy/2uN84bLt+kpOaYDevto7
ZYwk4GRuCnBUa9rxfK8R2svD//9MvFlKlEvPIbMIodNlc6UJyhlx2cykWSUbI3+JlEnpsHOBZ2w8
rsLxdhI4wIqsqy2QF2t+LVGZT96PfU2f4Xd1Tdln1fVcD9hDLqDyWWctQBEIbfrTK246iZyepi0w
uufbjbZaQsHFRA78Pf2cqxAkNTURyDA0NAwRrRXZsdO+KYpkH2rU95Z94cucMmf7VxTUU81kF6fr
wFD/AM753m4LSygWLwee346xgO+e77zn3v7GR7bHypkwewmyG61Bon4SOL3iY+AMRpZ+i2NRBngA
ym6mPocf8mXcfJUnf2qFS1JX6b9geLBMtwEZJXGtzSYIqfcn6LUnUNC6arhq+LOzUjBrrbpHckV2
JkEJZ7bEV+HTmHN4ygFsHa0lNL3oYPLKAqLpawL4qU6+XHUbJw8YqeYKP7ORYKw7BbhZmnx6KYJv
DSsNZFmn6e829Zeg1FB+4y6ruSC4TznScnN/U6/FGeazMf4oJgi4qv06uXfk1Sm7VsXfNWl1bxl0
/J8psWk1MCUiAi3aUOXGz0Uy+LX/1P/UkGwYCv101IyT3TXELLwenLuUObmOTGzs5K1Rua3UIUG8
MERru0ruXONuwzOHH+CXtaBDvsulO4qo3RJHz7KjMSpceg4qDS0mTFspQLN4i/gHEzIuohJuDFPQ
890bUhk5WuczP3VeJ0vKQ0ZfvBZLPaFJiCQ2cKzdXlRqRzsl5Uxab25yRuPckqUnmDSAf4mgyng6
XwM/c/KrJVCMNgmAHPDpx5NFiQJJk0OlXEIkKCX73Hu7+edZzsogKT3QtuLgmjCEeKxWeQyKcfL7
xdygpcyM5eph771fdClAniSGwti9TyYuu25LzWv7uYCGHos1TjojbGWV0mbVsk4HcSDWB2NqxyIA
O9frhRZGmyn/Q348M55L6XXsoHycbpIDwmu5lTkE7Zs31/oSPkXmfH1kD81exO+BrpCKJfKFZh8h
83Vw8GQDZdGlf4vpQGU7WgtmJwq0Mz5/0UtBN99xhKm33y0H0L4a5k4DBXiOrDJuAMkIuBylVW2F
qyh2xx9fs0WZVxU2fH5czyWykebZ/GFW623QyGy0xOoNLKm7Et2276NXg8I5HXbMGyVYvWxs9Snn
6roVJqNgpP+3oiEOYjESek5eiBN24nrCK31ORp34Z9zupH5S+wfJun7xCqZbkgjVaotKyB5i1zn7
7w7Y4T78+wyh0SpU9I17GG6QttJuJ8FSzQl9bDJYk0VHK68NVDNIrfkkgT3hCiWV8+Fol0eG4BBA
PXsy91n5/0+DSdVMG3LlH3vVCMEneLNq/Yavu1AREz2VYH6YwO40PsQagOEBvxZUpRJl+B4/lPU3
kpA6wUzCkCpqiEhhypbjvpcuv/x7SpsqroOPSu/5YCKcioNkLoSM0wT+OZ9q80iwzhegV2j6E24a
q529It1T+WvA1yRNZlY9uqk1CyY8E4g8QubC+kj9mVrl6omjuKLGD3YgSJZlfQ8gr3FFwsL4xMT1
xav+ZYOL9ubhsw2Toqh5jbInpOjaezIWKcVihqYmHyQQI5KU8DGFojl3x4rNaPA2BZJyT1GI4f/q
fX6tohJOm5X4zOtK9gXVxMzEwLgM0QT8nW/Rac4cErHvqm3kBOxVvvgw9efSbOydktmaPlUmMaj1
a89OeOOcd32MZ4fkkm+/P2TrY08JAkq3i4iP4DhdbHM0/GViGjrB3xiRnmKsJbhEB5aazutI1meS
CMGBjt/pf55bo46PMwzRec0n8YH5jY+YkRhlsN5VBttqxCrWIrhMS/8eS8mpKKllfPK0gO3J4EXs
BUybmNI57Npa7/w1xKxha6V6F9ehAdQqT3u5zZsFHWu6A9x7E6havSb2cKP29W879rVHNK40GfMP
fF8XKvSIqRlFxvQ66yP4HtMdGEDUE6jxVEUkPGugRlh+7f4tMsLin26RWXuJDItFqwBTZW5/YrML
0uGwrq+AnLQFU2Gei2Yth5HQuc1Anu9Fq9FhrtTNkkLvMDcdLIY1JrwudnD4JUksMUh9H0Z0JEFm
hCjSPLUqjDd6ChFnclln41rV4z+022i/vo1IaJqlB5MOCC/bSYbnz5rZ9j/eE4GlZ+9osM22Y1EG
+TrUkVx0tO0At+WvtubzYnqDqPuhXIv6/O2Zo+l2vz030G6jb/7QWiVyVhOsl1fJV6rGaMzeX1dO
HR70SUtPx4tafRvkv6Ej4T+BZAWp4yxqrnqR2PpG3KXSCtajW+EoNdW+uxRhrF2HxeLgs41sR8Dy
TJxdhGUZ9qN86cfn3spm5iC8fOeVKGmrwwfv66+LtS8CfLN6qQhtf+1cVP9XIeshTHvdkqF3zTqj
BYYk25FnddLJTn/shkcUGhrm10cfbhaA3U2CJvhXgWhN8oU52vK62ILUpYklMsApI1vM4ExoF6IA
waXw8Tlszr2BNwPkMjeOYLcRYRVIfXAQguuJfBWOAiQIP2nnmcTUIwqRZ8ZiOSlxYRUtcgT2XCDY
gF5OHhMlzcbajO/z6vUcH4KonWpfUsCpFv1iKDNK0AnVgWo45nFHB1ja+tt0q4hxmwU34PCCGlGz
OROHwEv+3aDItlqTVlD4Z/EgWBMfQ5TJtJlUzdHGRb06QUu167UyGDpnydazUCvnAVC+Zzgo9rdb
9/ju8g1p7xu+VINukgJdUpkIwA0XCAuoN4P3LfVUuodos9ZVM6rF9fGZzgUucWbaUZiNonf2GncH
zCTquQbeT+K/NorEH2XciklYeU+s5h55X78GhM5NLF73KqxvowKWssNtlGxhShvZjuy82oFaYiP4
rmJvOU1UsrX69bx2RkUbAVc/EuvEUrdXzRC9x6Q+0vtKS7YO0QCWUUtTC52R4dmhqaCEUJwK8Ve+
kNkHvCbp4oHYGV631itkOyR1OEKtDst1MxxXN+QIHxbsfyyUaGlO3rkw8IvfVWys/MNzwvSTLgI5
0khf/VK8mzCXtKu9dDJ22OFsM16KdqYDPLxTx9T8TBtPYQAWYvxK24OPLDGB751epfxOd0Bo2I1i
9cqP1VTZGjGpT/KXYWNMohI/ymUorZbUgXe5S7n/eL6lPGCw7mAILstg4xUWSYya4BdgMyT+XK/C
goV1biLR9W5QVdLZKXu9sJDXlHayL7kUlJs04+9X+HhugSd8Mq+5XWteLf8y+3w4DweAwRHMuNqK
VW/l5OHb9/1WSHpgpjRtCRD3Nvmt593iZn8xPN1Ar9mRORZPxSkiyr8BGkBF4110DzLEPqNnCq20
KTr4QEVu3p3ygSrf9htQwRpC3lPLms4Y7lfduyNHZWTBKSoQp2FwiIyeO3srWlV//fEA0S5GO2ke
CsyWE6z1hXdh/NSBvWyx9luWp1YWkIl12PX5BdE6gmXIn1J2sRkxW1DuwDecxKS3opht07alHNd4
0dAHl1NtVgxVS9y8XNRLUcZ0KyzL8i4faO+5Y3IfVBhZ/RGEYIDaEcC25WAqJm2rbiWlok4IMkSn
JS/zTyIyRgJqBmhSl4yeG2mw2mqaPutA6QIY0szsi2V74AlFiWCp+z8JWgd1s2XrPX34Xt+vjYIu
92mjpJ95wA2m5SFRw+2XV1ORpOERh7fqTL6KKK22683/iwsBA4O5ezcdhCPi2x1h2l5PIMeS5nn9
J5AH+PRlUtLbz9a5k2ZiGf9YSkMe+6Jxr0eymzFATuUBnDCXQNS6JFw41WTzrqq7CgqPUJTvnp3z
2Q2LpWPEWL4NUWtxm54g58GnT3nTLX9UPjMY7VV2SjK7NobKVGl0t+YBAFKZCqLdY+/KY6Cthydo
p19+C57lxqzm9RY5cPLiqEAkouJZx1O5cbTPNeRcxzLvyL1QuvxN7VIep/04W5IiA6ayFlx7o+47
/ptnCixXrjJ+JwopgwOj9gH+Y1/adh2FuneS0u70taRpWkllqAILpvovTSvIgW3tVrEw10z1NEWX
5D7544nP6EQLr1IXfXT1niMxptL71BazeUbqaYn39dK0Puq9qKwoFOgwDdZz+WJPilEWbqrKlYFC
oHfGaYN+cw0pDL21x4i6+W6KBS0TcfVmNlfPTW4CA8CNoVBUVVwtjJ5h0XYZzrtXPZHu06SDCC1L
vwbexU6sZPOmY43SVkPL3SMo5doeVOv6CUSb9MdhC+/dJZHtAHDTVpGS1jqKQKT171n3FNyJps4p
pzDYIC6sBM4aazDNR2OAvpQ2AYvMeUBhHM0W9ZXugMPYxfy/CMaYi4KElopIxosK+5Go9s5HZXZF
P1PvnaA9ob4MczMtqLdI6vqdlZfOaEvTUMm3pIAfzCVL0dA6D9xTM3ebb9XVMbfl9Y4fid16rhWU
9NW8afxbSMaL4ANihcVFT7X2FE6YpelvThrKYOnEI72mKA0YGi0FCeJdBSL9C1In91/+ttai5L4N
OV/wVLZENUyhjxIVX9LUEkvoClozmz6iKmgqMnlK9Du5JPcMNLR5H+wJFuK0gtGN0XrDohS2O27P
2TemCsK5KdZXa5MfXwX2wB75yCsUCnW3gDK1jLmTkkzrBRrO0EC3q64l/AuAv9V4FM39WTDKQ9hw
9RTmL7EvPeTlcqgoFiqn1OVVQlvxFmAdlaOYhxZKWJ4V2vvjcYCdtWtCWhREoNxgYZaaUpQlYqPk
2jMEPgc1nU3xFj6yVWzgm6MG7WFH+f+pkJL4/DoNxsOtDeATc+VpHd3kieM8FMdVshgPN/rJN2Xr
m+ca/FExe3UcbxEMBJ5QJi51hmYIyAOg14vLbIPYQbiGbYkEQGmvzLMmH9BGF4daFfOx0z6dE40D
CYxSFdk6/Erk5t0+hEAR/KzicHuitxEN7YiVgUyvyo4hos3Fu+/bEjSxoGY0T5BnIf9cGn+H97ni
CbTGl4MIsUa6a4CA1pkJwKpihYEVfB2WRrKcvj5qCQTsWKYIiMa1ASLtyoigeb78fQSejXAYW+aD
aYurFMp7GqMabCJK8oeEnb5NiRM9n8EmGuzcOW9UuOFt0n1y6wxGR76NtmXkKWtpTNYZe1+IwHCQ
VzgUuBOrPOdKEfkduAXxRJs24K7MLRk7WxtC1UBBxkGzxTRPJidltt5z1/HxIEKzjzQJr3nZfVsj
0fSCW8E2sH+Jvt8/aU3MllICzsjNEEPMOzlWd5lNecSe9YE6flQUBgWGnt763i1MqaxqYkLdpsMu
p9s7mES3xIYOkoi5OQx/7vYIAY6aaqShkSI5h1p/W/YkQLGXHmUHloUt0+qcli7uRhlIeEd7Vaq2
85qTrYTwcwyCMISIJZD5UxN7ZVzb+IS3sjNJsvgol24FSv0jJw7DaD3UBnyawKn9+5fqnT0rIDjD
1huVEvSUZlbO5eeccRKCabi6dquOL+0Js51x3Hhzu43j6uvqCccGNvs7MUiqIgumMav5lyNXfZ8Q
L8k7XCwUsrP+yrJfIl+pdEanOr2+fRA76seoqertozk8YwN7cRXAQlbE/2Lu9mq+CVKSBv+Tp0Tq
hFco0b1OMHTRzNqQ1g7sAdkVil3cSIQ7v+1H6BHapMr7bbG+wYopPR1Bab8uQATOaKeHjOKU54kV
ePp8raOjHyeJYS+VAFSFfCioiNiFV0TUOaZIRWdwhqPVWRH9RHAPrynpVpRqrxSLJMoYDAzmo4mH
9mmWO8bawmdba0fgJaMONEYl1Av0ztkFvAYekNecTrAIizdmpnTvssEp8yXvSWEAivFikId+N6jG
aya5KOUhxyJakrbvOekAKrXz/9viECTm/detX6sDCtGJCsZz1oxxswqdeRSrTd4v28NMkWAJxnuB
wMbuTOWTtMWohXeNvlwYp6kw0C8D+Hq9M3cNnh7o3MUA/ZVYZxBL78SD3cQ4DdwAepD1FYdw7MeB
dDCjY6LrJ9vELtoApToR7O+gwBbRs7oVeeZQpIM2yA25alQa4T1M82UiVxUkTw14p4Xx6sq1fwZg
Agq6A6/cQq2vvpWu0ZkecX5N9S2FarqllGo6HTRI/0GesNF6kjXs8eZr0VXLtQW8OABS/U32lzIl
XXRA7wnqdh3/KQSn5R2vbPRBSna93JsbStzEhEWwTajiDcBwvgpbhk3Sd8pQfqaDgusKyWU91VHc
NJQoKL0TMCPScKzk58ifcs+xclDo1xJqmbXaLz9zXGgtLkAqx51uGq+Do9rvO6lxYriK/kpkeAVt
YLTTT/mmITHpTgydnPjSIzIizhB/KzscnPWgQRZtiWZjV0z7g3GNyZAlRNCO5HgmdZap7omxtN8K
807kmSOeZqYD9y+BiRebOmSJmy2hPV56kk4ogv7yVSo/eFRXVdOPipw0koLxmW/SOQ6ef6SUQjet
Dy+knrNAN0pPgiIwTOrueTzTVkqc/OwA5LYssl7A3iK6qdH6KAHRkMvRaWhNaxPtk9YzTT8aENnz
mHTFDflM6tDJRm7cYJPAKZfv/SD+DqwPYOoIj1aESFywBhBh6ihyKExcwXBOs83XqYO2oIxoEj8p
iMbf/NhJ1JlZwQkb0OXBLJ9Z2yz2JU4QcjdN/KboudpmYi2ofaswYEzcEoHCFiZcnImNDScocEBH
1Y+QqIphlCTAjEw1WhMpa7TkHlS6F8ivAw0Nc1jv/K7HfqpJGRAdNG8jOaMk0RQCTLq1lLgnu9HQ
3RoD+AEX4qnLs65sZ79SD2euihGOwwWfhP6li0s2nKx/hcBwEoJbu11b+ODZJT2thnCUhd/pb1tO
fctprZksovTuEvXexD6Rf6efBgD1jg4Cg9nuNSJHEsEqhrPOjbqJcmUvzhkSPdzSfFpsp5rYB5Vq
+N24HaBx6nS0VWbbCP7ZHG6/h4F4jXB5jA35Hd8PaklKVGMGPgmwdGMJQN3jeOW13/Ds4f+3Wux/
AojAGQI0vHWCxwi9bdZqAPU6tPo8QX2MHE77rCvB7xQhT+l/lphy3E+e+vmzUFTYH12WpPRPzpgs
X0yqiToVNlIlQxXmxf+y8PAsp+l6CZBvCteJdov2+IHWPsbh2ETZ8/P5YR1BHFKPs2ueFaxCO5ju
fmeC8Mt17wW1svnZmxqr1qGIXnFc+RL9WtnbCMq/3Xx6jsoC9XLJkcRur8bR5Y5Qh94+9X4EbfTs
T/4ycmkaSdicvSJSpOJ2IBxJhZJPkpS70G4SHNew/3qsUtSSiVcpvd0d27CrvHGaFqgme5wavm0B
24hTEqUyMZPOwHq0QAkCSknf778lxKJxaM7rWwqdz9RMjAQ4iPAnzjU8aPE8XcxS/bUkrJEwlphZ
SG/iOlmd9L4IXkyff9leCOlLHatUnScadHnW1/0S9epSc7up1Ih3wEAdsX+UnxAJ4CJ1ikee+c/N
WRQfCZ1Q/92Oma6bll2EyplPNZt+L17FdtAgonKy7uiYNNjukPDjVQedZLgdMeAPqAGSAXJrQ4GV
bp8jwC2Y/kCrNZ0QCDUon9cQej5bRDfDH+Bc2JhOtI0tITePodLq4LHS/snEZwCkb8ryT4WHC3ph
Era1vDeBoIwDOB3RvclOfcTxEbl3fG5/oKXmYYg22UeyZjcPTl6nQqzinyC6Iwt8IDraRDcfMlKt
EBLiyGQE6qWGj98PMgA8Gv/5M/rI3uinRF3XEWCDjwcef8IbSh1JvIruqTaQQQ8YFSQiaJUI9sUz
S6pipsbttKUYIzTBbX7tk7oPZ+AMFLAKa2jJbzpSXn8r5J2cDvYNyajzJY0vhtemIYLaJMCxhjOv
Sry5iZJoVZcQy+int6gnsJI2dCFtF33HHxYXVLvl7ag447MtCasWvg+0KDACVwqJqyLgUKsypyme
UWAjfUt1Dojvp3WHZDYhL32SrRxhX0rqLbxdIEIjG/mrkrVXxF+Mj1O8IG22mgxmxW4URasnHK6S
HCm0982IiCheMW+ngc5H/3nenFBcqE0Z38QfX5RyIPon8W5OIE5pceGRtgeYDYy3T+EkvClIt4Ty
5acWrWv/RzI7cB3hFHU5b/WlQuTtDSZPeFnf3y3PPO1Lz7DIBSYjonduzkY/seqyZ3F6dCUK36UC
idcAAxw6nwqpzsxD1cGM1B1535yofdLEnGf8HWYPc/y2M2cpJisgdvLUY1HO9wUvghHkIjAh4fLv
jULqHlT4+/66smRa92KzcJi+gg0ab+7IygoOai6NXCk6XIG3+Yfl1d41lxAGGcYgqRnSQoEwNsxg
KXwNn30aIgnr0vKW/BvSKsaVbo6+CoHZQfraRM4esyVKwpeP0Lvkg75u0t3PJVKpGshsLmq2Sy+g
p/F+l/uDB0L12B/2BuqILEOrhBgUXfKehXtZbcZkYow7DKz5S2sbVMCLxDFiETyx3q7RbSebH9ZO
OwxhxqgSjtJczKouZp02FHBtdx5NDvj4ZDV5RfzVWp7nPgZ0ZgK3A2zLsSeLpllM4dQawQQgxjp1
mYC2y0g4WPGG+ia1lUTEoqBKpEAiJXDfUgnwCTxlq7bMtGkVCoNz36DLLDp/3izS3UNodWjdDr1U
PCmplHzdlT+dR66ilRkPpBy/escnaM9/rd2BCMhe8xyHvU2rVBxJC+UF6Nn3Mot9ZNytwmUKTtvS
FCmqWs77hA5ccW0wYMqX68vrfVtxvZTpuBf3eSIbESdv7jn6T1G2nXoxJzSG0PY0uaD3ycSHvVxJ
iyEkVQYUuxN8VL1zKono5hbQrnk2Mx73UwI+oqmxPHjarkRsZOe5uLSuV9fMmwhQs2jJXcnVuzW9
VzclCd3s12MIMkSLlTDEldsfu2F0amJTP8fPmvJM2v3DER1Lpjp/aqQungGzATaeWfmvUZjKOU89
XYmcC8GDyD/NffwWVWKVDgRrUkYV4ge2bbPyGHbPjtY5gGetSZgpoz3yN5ny84I+H208/0VGZGbl
0/IhWNIEeAB+62eWVowNIIthgVtgbFHlw+lS9EG76igINgXLVUxS0N+XQR3+TpRA4R4KnRFXdS9L
/7PIeI/67zcgml6hLhh6P5QWilYScYaMg9pt6R/x+YN39kLTVLWXv7Ok7PVf+Jmp/6jyslrrbO9b
rlTPCYT6yU2tD2FSgnZgqRXYyeQAtFDaX/+TICfB/Evs7rz/3moa22Vh2w7qrJRvb4X8+TRvpzyZ
94rPXFpOMqNj0eRK4JJijLBdudIa+TcaP9HcC+nG6bvehdzyx1YXkcCxyW8hHK/Nwz3L+EVlCoXB
SGxfcTDsygbD9qd6DHc95PICW8MilsM814Z14svf9lIz6gDHVhOYfD1XRDb30FKTq4owbWXRqsZA
HFieScNl9ctVZ+mj4PErUBk8tFqJ05Yy/aOrVWZgxm0NhTBMQ4RDPE3aboXXFxnqOzU/MKtlRxOX
9yZPC+gnFexoPlYnLsMiw6SP8uc/4UzTWZBSRWr/GIkPf8NtNf75d2epgSjK5+Ior29b3wdeX0A7
4KQfXLfLz8YTIm21A2b6WbaIkTVcB/lU8+BY85D3EN160Qk/bCDk39iHlfJ9A8iW+IxTUStKRPhs
l/BYHWHGlTSuLuwQSWZFMNm1+S0XMoofutbpggAd+YMDdcR57nXboIxmHJgbwP9tCiUNn4U0BuGx
WeijOLmoZmrLddOETf7VH/BHVHDPEFfn5BnPzPohPlpAM9/BIkMa5G7CnOGw0o/ILFaRzfPDqBkb
lVmbCVgfH9LPduLpWSj2TQbaIOsspwvwTckYU6ldm32uDZrD+adLRyQUfUrrcQh/VZhjdtTd0D79
PtOPw7qCPirofhXjcBQUVIZSE+a98sLbdIf+aFjaADShYy1qkIFKepnR2qV+/O4wrhFmySEpaP4X
70pnhZk8KCioyP9PcFMvA+gPWRBoxguB0e1ElT7G1U3S04Qtl7Q23bb39uiFveaGGZ6wCfe1t11S
Pty9wjl/HA5JRTkmkh6KLNpCGhwVf0Aw/EmhkBb52WhR5b+Qw9XdcRz24sRWi3n0JFE6B9WAyjsY
A0DKYfn7jpAq7O33uCSW9VNN5MSx/koQu+FksU+07Gl7OV8TPDi6wZHCbqVHhDU8qiA8249o0D/d
+Bn/1slrfJ6+rjWX6Zl1swcLb+JFKImQCYcK9g0R72pMt55dvrH6WDXJSrDpfzW6cRmuQzAy5v5B
iKXpuzdItTr6wDyPSjGeOVooGlnsKvQFGL6brAHEk4C1/tA5DHe52noHhzR52bmx3SW1CRWygWw8
VlH1iis5YRvfZonZo3xT1M3ERc3Ru3IOcQ7eagoiDfQ+j6tBIhjYR9Qd5VYFA+O2SvfAtIFxqq9A
BIA5/9f/9OZwnHH+brUB86adZa0MoMntMt25ABmqDlxEIbFFJ6rWI/kCoAI3i2efHcSbsAeBMFbQ
nnahy5Y3YkaaWxjYDJUdpeav3dHuboK5VvsFTb6pNoXj8BtoUN3qPtxP8zP1GF4ktsWMA2YU+vCJ
EUxxhNGIgDqSTlCOl4YjO3uWqEFP0OsR89wYsLHgPFPwYPcIhZTfhO4la1UIYA2bDkGbVNuhVttN
1Did1LYvmqRar0pkDOUYqJSdYBqyV5xZVwvEXXlAkhKwx+hojtmUcn5oxhxaj9VxQreWGl1DG0Ex
pAAfiuyzE12PDWkLCES7MFNjxF03SL0bep+CotTXm0+4Dux+/kWuRGj3GSNoAlJHu5jzaoxfQaC9
bHv9ueSQcTiZm2MVwSrx0EyLBbNvcdzwJby4XAcPvZhuMkTXCMXr319NS/mCVwgnnm5Givz0MaKY
MDxbrKTar2mnDsDj0B/P3wygHOELZA05fUtcM2UEfopfQANbZuArXVCJwd16IwFD23PXsh14etEf
x6lkwKabhBViV/Ejv6tO0xWjiccCdgW64kndPnbxc0EQ546n97Zs6Q149MsndGdWAA5grIt6K53S
tw7Lh1wb2SIeSgUh069F8OwkEmXvFQ7raywKYaq90JPIFwYuioS1UmmcuNENecVbeSuU++evxfmA
8wBL2TSULZG8rg+LazwBpzTDLoIeBjtHCzeQQRgRg/uRjMaXRphnwqnIfn73ByM8V+Hbh2xMxWJ3
DJG44QN2OvbGEZMtehrJykQADPZ85XrQc5My8FgNsYbmyAVhAJO9SGs45p5Lf4U55Q5+jQE5g012
SptGxjjEjEdbG6sJDmwhD4NGXsUFTEUkvVr+tWUCv++jwKQCmCjfZISagpCsWHQm12zWzT7AMw3E
b3XwJpKs+SKahrDIqBeC00b6cEJblEjbDJhQF+DMZSvP9loVCGtTZ7sns3QYM/tKeowuBY8MA+yb
ccf1k0KBlThDyiAnqPK4RZkf9es3M+pf/in6SXSrCNtTfpmUyuRzEu/iLkmLOjOuYK+J6YSf1Kqe
yYgtux7I9fqTQwp3AX0xOjXhyMNVZQV8cB3bPEHdqj7KfIc/aSL5LCRgkcjPUlEAG9tF4LT7dy5N
2i4vIzGGf0pWh9gYNwXpBkl3fdsKbedbfwvxB8FxWq/dyF7GNFJobXbOI0tbsxMjc9FkJGyV4iAE
3qbJfoS/iXzbcAkhHaivwxhC49ZX0XX7JVNodGkO/dNNtePQCVbRFivA3e6UaWn+9mHTeedTdxs/
FQsIZdHxkPpfcPXF3dkELklPIc7SJ3nLfIFhsGmyxR3wbkabMwggHIx8K9D4i8QSBApNsov4jBt3
dpje/s2c8yPT2RhZMhL+0tm6gOQIM4JSSoyZhs417TgbAPNufgT/slsXiW5CUMNjaW97DrYFhp4Y
XWTZvGyuK3mGqEZraLecVXBDmdOapgh7/KTVugi2c3C8gIb5/+AzcvlBkLZKt5I1Wv7FmxWfbbhg
M1N37j+tUzzpqm18I1AMdTktVgfM7NTEfHKK9XhZmnkbEQqxSWH43D3Pq8pCLmOaau6EP6PuaEFT
eW5CHRBzlp3gDe1+lmCHQz3yyEt6Lr1OenBwCofIW/wv8tMeI5VoJNbMCbBG7K2/7H1FnkDGnJ7F
72lEHDnKTLtn+SFHpMRnFjzmcah39WgsJLO0ALv6R5gU3QozHXfqDXB/UfW2cDQyMIESWE1vBVPC
WWyhvV21N6c/jKeFALL7XhI85X6Uvn9ISZ11B2kn59zQwi4O4E7z4TtLG/V4/7Wr/3kt2DK/a/2V
0vhVYz/DXmVcttnFNePgglkfp09M0OVaWQZB8TqSz4hUwaj0iSdL7rlq6OQdvlUr8gzcj8r1/mVB
aXcse9IcxRfiCu3NuHdTsf7rHWNGIDrpPhMYV2zwkZbFIuwmBah1qsdf5uSWQQFLA7gIPfMbY7dn
l6VIQB8/Cg+7HBhR7hX/sslJ1KhjU9WbsronH2xY2K6zFD6igwJuXnO9rewhBll13Y+5gVTO1Rti
10t9sAwTYt+jOyZf0NWcVdc/gL4UXn1XMFRTM5mkgbjonqyqJRooINQSGfNVQOI7QvzgswUadlCI
L/d6N6K8mhIcyBHOOnBO6fdq0E86WqViQoH9G0RYinxH7VKptNiNJleEOgEURRQlIaOWR+axZikq
mTFZnvyNkb6N4PT0G6eX/NU0Qi/QyC4HrBuRUbLbyJK9KPR46m53EEbeBAooHa5+I7wI9shd/MxU
J92/MGqM7xs1GuY6vO0Bj/KxboqzWC8gD67rt4SLE0wvqKIhzj35Ek3ujMzOIMY20A/FGOMtXc1R
6UVkYqNKXYdpgoNTEx8DX1QzCAL/SMXtI73ml0N+qli6hqNjWZs9+nkSPxWOOTACzYD7ndwD+2QV
GfxdhjA1T/VKFjM3igzMsbaAfLOZKLKxMBcytjMx+l81OVTN/MGpCKNLXbA/4XF1+7lFSZ/lV+ii
kvWKQazDTIwb4v+AtdDUCb6qk3MXYeWIRFEvp69JuowLe6/h3zyYIQ1U03Jtn/iaQlShaYXbnaIX
0QmBz+sd0w8dXAFjFGT/h9coKa5N/gtgcEICc1axsx3uh061NSknJnyqJqWFRpgbz7+bYOtb6wfi
ovuKElQED8aRU5CNACZdcPaetb5/lNhH2IbVDpc829vz5Lz6kZDDvRG9tFTLDZkTiS6WfBGbNbV6
58imJXBx2Bfm2eE/w1Zh4aRhcEnXiOU8bfO6KZqv29VkSVQGNDKFsPGAezeX9+mxhJdx/JXndgRA
2EjINSSqiyYg20xOP8x7lqEWkvHNNokUHTqnKTm43pGcIegStPiU7XhFnMvaOWyHOFks9grdeKaG
ZB7tLgnr/7s/zLEPKHBkR+XCxFuy+zTzqk15+yutqyHsNSSMbRpew3QgsH/H+sUvV0g5i9Nc3xqn
J3kD/hpbIUEILQ7/BDEkruECviZscfhOoCW2ZYrzZI6DSTFfDQbCCYo9nuIKKmQb+xZ436+OSlIp
4vEiVoOewao1F4Mwf8hIcs7UEMj13B/DpLbZ9SDgKQS7eN1R2EEioH1BXgpyggk+8R7yptARqOha
RiVBha7nvvUdzrzmN4cddwzgvXmLE6Fq/mb079Qxnuv5o2g39Nw1G2tm68qoIFX1F4Ides1yI+Ah
W492JL6BlXv1W8w6MTnkmAIWCZD4x8E1N3eEhE4WbqJGamTZ59epeEWKemSvVgvKDfNKKVfAQZN9
d+D+lBXVScLV5TxeaA68p9QSAlBDFwdyXrAfD6DVYUT6XGlE+ooYgenV+RNrC+BbDa0DgH8JLAdG
eo+md6+bMpuv3DXRR55Qe/ZEUnKbU1W3aroLewgF1jsFVdtG94F79GufhUcnV7Fonu63A1NJLecm
M57+UfYM9mXJEp+yaV9j9y/zQ+4Hdcq+tzoHbsmVhphbhf8PQ/uESb7GJ+x5WjKhwHfEt2uHikxg
bOh3WMSW9JQ41VewJnYnJY11K1VEU46Xj59Tne8yOALZwEjTbw4ERN0vZB4VAlznRL+fb+ad7xjw
hc/rfbGHLtYsTRaeDI0fgFe6/nwfeJ7zWPrzUDRk7TV2Edjs0YVUkoKH5YzzGYpJ19iQDbPEm7Q6
Z3Wg9fjpW4BOLq8aORTrBG9JC2t5reHo3XWmWRHwHQLqzx1nRGauAYJ6Cs1i+KK3e3Qsux+odhxQ
yU6Yn1wk6G+XLgDXp6v29J4GxNdHrrJRYeWTWE6kzOvhZhzZzR+QOb9dkH/cCFsMZpypKSF1EQLz
GiWU7VvAkFpDAAqjgOU1Mh5O+XQVvjTXJk66HrXDX1arFBKKrD3KTlHrZL69WCAGHAQpjv5mEAOf
gnlWstrrwsgcRYr1OEgVWIA2DqE1oLQOgjJfprEFTJtBYHo/Dq3/xD0sI2yCRKPGDd0oFNbYKgnr
eS0t08P8rfgZbk9BL3FP63pD/gGFrpFkPBwBje7HhpeBm7l6HZRbvQO7v74RLMo3YwdlFaU/nxA5
ZbKnEhhl/GvZs3VJ+h+SWGyKWIfszeZNckZKOTo52LtUQJAwpDU/nwSNNjBD3sJ9pKjo39GDxync
rKNLDN/DGMFrasSte3iN5+L6/hMtG2ojlpxGlbJaBCslKGdxb1dX3Nug2PsRBI8MaFo2km1gnzpG
ZmKWfgsfctjNNxTqvGvRnWGcrbNvZ3gjhL+EHrPM3meR0FLK/BIM5EFgFuhTJwypc3RbJy3CMznk
gat+zhCRdW5iWJIXEBpQ5Q+ttu4F5xN0/yW6FWDxg0Q8IheTEDBka+45WPCuUBZ0GIaVH8xpZPxC
GIP1jxnDAmS/oCyxd931yy7bLFWuvLHVwOOnMdm81h/FliZI4bJYV62FNcuSbT3wnJl5BscL8aVL
38ztxNK+R+SBK04sVFKYIM1lZrWqO5qmBccMdsWJ58miUNxYRs9cB5Opdfy6lDbtP7CI+F6/XhH5
MLcoKKz7qCvPGU5CafspaEE4fpvJQcwqmsIk/uRhVZdnqfTCdO0pe/E9jHMYaDHeVcbUEOEdCVh6
AWaiOqLfpbPXNjs0lHQwROL3v4MIaFjZsLJTmd4HdtvwIuOdvLS7aHxzCJ1cAGOgEpY8wPmQrdtO
FqLhNQ7/MAxgfLU3b9pZlMLXsS/4oD24uPcq3cPSbdZ30yZ/kn1PIr/JN4nIKr5gwzkK2pBD4Pnu
tt4/6T/HKJ2GV3FKYNCtOt4To7VPp6kXXfmgYjH1KdJpxaq9pBpHdq7cV8dJBiWUJfAJzyZ6Y0mo
rRlU57I8Q+vRzfnaEr8qDvtfL8mTwb83thZKr3VFIbyVYiSg6yxjIeE1QCUbTQzL2FT4gszC7Oux
fbmsWx97h4z7k6A0DbNcqk/KrT/Gr5/+R9ivi6pp9dRb1k9ur6oJqe1n7oz49b8finJ3+5IUjguv
fQam7zEBpSzfOdyxA1+zEK35OYJP7FxnrzHR6neXpwmEyR14WzBB9F4zpJcAZtRQbbSrb83uE+wG
Q7D+rUM5Q+bA0uBdJpLLCaGj9MTGxNIkdR+73f9iBNqJtlEvpxEt7jrAXb2N8JZ4ssPg4jM/Ur2S
EekQ4wr2fNq/BJ96tCoXOiEQbg9u1qVck73qvxT71qhnWajI7AwLtqxJ/qcFabgiwpGMe5pAjyD/
Dk6v+uMKcWvGGTT945pTt0fCxOELp2K2YfjHGf6wG2OdTbVuXSW4i4j3FJOQLaGY6yZf/lvnT8fv
Z8rP3Fo8Zc1XvOJHAV+40CtUWX5ug4/QctkVkVFcTnZz3OjJTuxWUvkAm64OpaPAE900J7Wkm80J
mK/nfCJ0JmOiyb4Ff4mWU+9ADqyJljUAcS/5/i2yfquOC5wy0OB1jcvlZ4Ur404Boq+PpXrIwXDS
weoxOs6Q5NaD9nLu0dB1wkWYyE8ZGdg7MXZ8weEURMSe4S41vTomHd0faoqYDOWMP0ajX+G7GKEQ
LneZpSTTkmN+adk+EO68LlvfqkR/oCW5yyZ7vPr1hQcnuIxyfLcTctt3sX33f9DP2E2HCiP0Lpwn
v/uo5OuuHYWFPq70GUZSk418vkCtcJnk8o/o/dkHRDWAc+l1esFWI9NNcBkW8mHAGAslfF7L4dQe
7PXgahH6JgLmRMvnb4LS5Q+eOmncSUj0bn++FD+a6mWJkOn/i2vcahJPmii0jlwyvxRGH9MCvo/8
x9hqwrmS+FSCmTetKkGj7dFvJ8BEZsN8s6GDZ7e8tBkBZtd3p0xUJ3rJJ1c5azV9r2vJtmJurADg
TTn7JvFZf8sK0UyUtwLxQQuWAbcVegCXAk7cT3mObHNh8IWkryFF2LWkjKS82oqvR2HizkJAHxsz
3fE8BQ/vYe4gRa1+cgpuulbwgazLI8oziCvvT5WRyxG7D9XMmpqtkQ34WrXufzGwpK0S0FvCFWbY
PyJ8GPa95td8AhB/tfheELOYcfRcNnmXjLPuo5O0UVPy6YGPOu6/+3y+XMNQNHGsfTUEFvGmunrl
Hc07fY2/KpgQTC7yYlRosLR+zNkg9NOaFAHUsr9g/sgm3s6+yMb81UMtXQuPCjRryhGAxfswLWbM
19XesUiSwNpWCabFcIh85h30ftFve1s040FpHCOPR+DbCFNgNKyUa5VpTAfmo2d1R+0L5QkDCHb9
R4licCOG53BWOOr6gigwWrJaSQG2pZuIyGShBMShhFgFodPRePIkRVDrTGPmpql7Z2UdS9cRelH+
rs59Ox1GbXrkMYNhY5IcxIOHSLulvHYf6AFMt/JFOSsVqrjRAAA85ZoUtKREuvieYxxY7mtRg9CB
LKa+eiZEkrB7lo2smifXKnYd9jr+0y5LzNY6HwLRSK/oDkPC+AQinRxy0HyRh9DSHZbldIS6kaLR
GPezMfcW3bQ0u42L2lg/oEdo6C1bRtu0O+DjDNqM6d9bUdyeg9FAyf+xhv+vnbbh4ohrJWomPlp/
2pjWMGTq8fcxO8r/KcZxfEWZ3oMUisTvggUtl8b7IDMHO6LK8k8kOP+XVka+dFF7Vb47JAnEAI1q
NmA+6qXR9mq4ZBBt/SdRdKwbDe+Q85M6axtJcz7vf93fqWI+UueWq6rXnUnf7j8DHN8wmpENnVY0
jnmbqtfd4PpYW2uH8m+pOf+gBIwjPN/T3tZj/kyUpCFdPKse/+3MNq2NfHYtOXdKI3Nvx0OypHZt
XGIzZfJZKLSph8ZkJqrUm1uZQeV96nxHLYtk639ziKmI3HaJqPijBxq/VOmeCx/X8VSP2B+2wjxX
OI+R2lN9F2fk0xXMXAHWh8sfvSBku9M48lMyHWGJG0pmO9cezCkPBYMh62mKlZTdS/y41/A+BcOZ
yeRqgHyR6JDsHqlaanO39CVYohIjqpxmMfJ/5P1diQgAr+zuWmxQiFh0WG/U3pgB+K+I7UHifzFP
I6kCr4RLpSMpRIwir+2gakyySEFZEZVZQvIfw6nyezcqkRPAk9nI0zo9ElAS+6x3OVERsz/oIxXB
BMvOuXM5c5alekl53BogFzQL9dTLopPRxLauAMs/nRZ5RY3eN2m4vUY0to1dNFOU13gruyA74J+9
S4vgNoD+w4HZVNLUQTrBj0vFgchjalg1gX4c9UzBtaqtsWV+blYPYm+U7t3ki3SNn63QhVwiAC1o
h9FwYQkG2NIw3hyjtBFhX/W2QRWo5+EjKJ1KDBBaFkfC/6hNKsXxrH+BDF8mlVWam+rFdik5Z7Et
jTzGeVJNtm5OJZHtEfcT+5VrHhO5Unw3/ibHJndAuh+TNOU5z3dVXwtRbwR4KOgKk2OJ9NRLfBBI
s/WXL+hBPUKEcEMt0XhS1SBNrHYeAPALz/ks7OnoXxlslKCUAzVrVR4jdf5l4JPutK5AZmxzK10+
nTbGJHEKRr2QlIrY3x6Ec9RbD22CxvixwQPRHTthl0a7dr8eBhh5jYVaPWZTLhLEvpqjFLph/s6y
mrqi17iViZlnMiyozS23sP1jP39q+PO3LnYCWPoE68jYlBlxZguvRzEham6R9CFVeHmaRai29iFp
INL7NCgWdDy22ztlF9Hu5/BlhndvZmKm6d5f/uGxSyM/Zz7Ztv71i5kttWn1GzCYLx1m+8TtXUUx
1YI/ajmmAG3TeicX+c553gegHdb+jwF80tiVWA6Lt6hYKdtgxDTO4NWMUqAru7ax6zDo7jglimBn
guAvHixhLQtcfyI+P9t18LX/3xqj2lbasn3WbxEG+4+j9XoVXl0SMvBK+FmUPFjZYTavDi4XjjRl
aRdEfEcU+M9C+mOghgfJNcCjZguVBOo4W6FMlYlfoaSdjlgqoMLi79nGyjwheIjxStOsyADjNrjC
C05wh05fgK/ZIt1Z4cFBSNm00q41EVVZyo/bUGudclFCunzA177LkrPmlLYQxgSZ1QOzkPGX/h1H
gZ4EWVwtJz1r0gmuKvGwC3y4AtuATdpzgjFyzUraC9c8zC0LZpsXr7h6pmGiIztqnin/uVfGRw7Z
QsKGvD2n9UAMZiCdSshjnISywyxrGDdzo+SE/Yv+PuH7wk8K1HuIq2hUjegdoNFTodxFXSV8cWHL
gaSjAoYEPNhTjjww9/bepuKwz8Q/QCFVPJrnKKtvRM36DOIhTg1bOVNZnpE6OQX9D7Z1qRmtMyPO
1stpmMdfVjcHcqKljWemR2VFB+aS1dMO+8Abja8bCCiriv5dXLNz0Rz3s2GZv/gL9dYjjQrbwm5M
sJMnMwmw0/fTi/PNbkti26bNxBjDXkNEIFgzQof+HgipAUveOD7noG/6/oVkRGeN3NG+IXzUUu7P
j9cNdmgvyqtdDLvBsQvfHHnWQcmKx5pXqGNmOHXilRg1PMFzkmbIZAfL6+UQU/XxVVD5DbRxXeZJ
7binTDZC/99hbDNXrPsfn0bNTKRnrac26Jbd0Aje3q+lrHwO160igTKjniV3I9MmNIoERvtqimVb
hll8I0/MrnjkHmUIeBPFzi9GqNbf+LRlCEH59gko45ZCY83K3dHTcD8Y1kuOvE9UOrIbsqfuHgHI
YDHKH1UfrwFXXWgHc6J9fK7kV4Acu84hgC6OIhhUoHrIVUGZynbjunRRQ3sb28ZX4iMMvDgR5+u1
jGp3XxCxmvonGB2EPcsctNJyCV+/QydifD/UZHQa7ntmmFxh3w71P1Jbcz+DJhSFPDunS1/AJr1u
OevfVh3meApl9lRx0L3ixy4Us/NSsbHDup7tnHdZIHJBQx5jb3t+LK+6wlVqAIUlkHWX6sI4L8eL
utR/Q98aN3SGyRFuegDghyyEUUd3hd+OJLOAaoyEPOZHPqsKuPY+kZfCwTkS4X12PfrySMVkbKyp
Ie7dTjX8ewVBcjuYZc22GMxris+RqFyIgg2mwWawVJkDmQ9ftK1GhhnAj0RosAVey7BJh6f2eAHO
Acz8AXljeNCHmK7pt5jmuIky9n6Y0L7BEKlFqxhOh0RlOlzCfDhOdeRPSqJ2dCU+O3kvj8MWXtqO
PAtBFtnVySxVgbkmt7dBQwevgO8OmSAVwfmvoiWWV7H8VJKt7tE+H1gsf1pMCafntbHpj65Pn0bt
VDe5yPeOblFs9+IZzblCbTHfpBkZ/KBSd63GaiDZhDnEvG/9FjiFF1FEHl27/PBzBvNn9sckKtrD
8izehXEiSmmd39uVGZSIJdTaRpJQNkzuBQFmm5pefFoxr96PfynWXA3qQOdP2matHCm+LjMFzroV
tmdbVixewGkyeedV9hv7C2NRP+bxpvM1TjulF1gcqh32dKeWAcgX6Ts1rGrwOEUr6mR6Yy3yFw2D
PlbLBenuAlxTOX69KMkYxnYlqL7aPquSPGVGU8axmzy6VfjZDOsfmVWv6vPbz5qtb5CQgT0/Czjz
hCiJgiWBi+X0epaChy4qYtcacPRhxouP0GB8r4agm7J/RYcDfmKUERtzBAGq0Ycx2cRucS8uNIZj
+LSsJUtYNeKke2NJOrVJ8gYSJgBGfK7oVQJ5fo3zt2gpEyjr9hHHcQTKXIYprARCDWa/TylTxgNw
zKPwIOXG+Eh5tNCyV/ZsnGbw8UMPsFn3hy7R4Rjeh+S0OcuDgCBXQ35ndAdvLVSc8sj7b5WJSxJg
HnEXlCeNSXQZWqzldG/TKBkwzomcqm8GEKcRhWIp6P/Bvv2VeElZ4HaPV5EC76xsL1NuiXTH0ZQK
hNjsfe2TuSWHViLDsD2aa2tJX+1OYxAnVsMXVseCdgTYyjbzlseESQjLqw/8ns1NMAlPas+I8kkP
O3mEoOuoCF1wAucqJ7W0AWoPi3qkiiPp+y5KvlV76LSySuNVY/MhbiOoXurtKWbAg0lJGssjXOuX
6WUFys0X6rmMm8rleQ/t+HSKRUKTep0V1VNcdnHDOnsSlXGKpSuKUHgU7rTqck3LPCGBtH/FJtNs
2nZbmpZaI1KxCx6joIqWY9fdnWqBTsbG0nLm0CWfvwNeBYbZ+G4q0zmvxrwCqBvVP9UlH/iCjT+p
dY+3NzzbEoiHKVqC/z35VkbcZHQW73SsmBgBMBInINVkyN1s5g1ZkpNzuDRspd4OWvaC/1JzYSAs
uOSYhTjFhe2cQ95ttt12eJqGZPLcV81R/IVAaMTdhCYR2HwllTkL8NByChPzd6JKaYUrQRZPoyF6
xC7KFdJBpsuTds+0kWG5mUQiUVNbOq+1j78/NU0Qn9KU1pyAeggxRHi/KTj0QJh8nE0L/HCFD2hy
B6o0NTJLIIG0qbfDLKdfrXKZqN6MbkPWw+24z5ILexJcIam4AusiSGusy+Zmawvukt7OWuC8LRJQ
ts0WfAinq9GZKktkb4msHlJqh67Oae3zS5BbCnQXMrs7X5CpnKFau4yYUfRrUU2lRfkMwM4sNNM5
xr/1CUkqQULz9MSw7V2cXBUQXH13QJUAb+kOlS72RCrC5ySE/BC6VXRMKDx0ncXKqNVTELd6Ucjr
OEPIdMNIbR42yi8FtYuQw1naI1ZxTRnK34t+5EW6VeAOehv9wBi5Hyxhg2p7pPNwzZiCOsT8i3kt
Jmg2w8TroLVLK8ETg6FDZhrrSFx8GsyWzx5WiA89f6ATIUfYwsVN2WmbN+7y8SuEtKNk7WXpKijy
/qnSbq8Phgr8Y9Rw00Oh6jm0HRoxSNR2ZcESJ+IGNqSFkj/oIykzBRA4RDOveRV5Z6jW0JKDL5gu
2KJKCi6CXgcZtcaGFz3jRUIMEPr9XyI02Y8ezMfd8HPhAj6SSzSchhC9RAdCphDy2P7u/o+LlUF5
nB5Kdnf6U0UFw4jHoYqllnYkCTSNGKfFKS8JlGwEEeXlszINSH3eCbUo3hLMiiBxYY4WLa9zvBYT
/mnduhNv8JXKppfv5vMHMpcdSmNadE6GsZSZYBmlOe3c/rV4H9+YaPq3sX6/+yxlieiryaA0nVLL
6T9oZPUOBuoFSnQbsApkwyh5s9HzuqRHuJPJV5fGL2owKjBiQ4krqOj/5i7M5zCTk3Qa8/meJ7Mi
WP86DYXpj8pJMWzo/qA13C0hUA/qcovAmJnB8AkjrMhSk1ygQ3u/p7vLvSK7s3apAcpVWYXxbY5s
Pb8XtiF5GzPvhN6qjtlE7LUWAcC4TMF+OsPInY7KVdlyDbzinHsv2NP/on1D12vQctJIW2MNdupl
NjpNgTqY3f5edjbOLpuxxMKWZs21Jaqe0rxsOtqT1Ul7r2bikApCeO9xpTry9eLJcC+JBZMJa/MY
yUuGe9YqaD3jOBmqweLyCF75JKHPB7ZR8qP5ULW8tFuiV6c38Sm41OLXgAxOXg4wR1g0KJhiFKsg
udpCKBObbx8UXFso8qH7eYC/ZSbPJQLkWn2f7RYrw1i0xMmTWAsjtzKMtiTizcQutWzm+msZAsW4
VJqxRhrZ6SbKhLsDwsWSfhU+k8FAHoiOfkxphBjjI4RFjjRJk/Fxu3aANHnSCIDGIwmIvKCW+6Je
HKyUKoQ/FZ64qDDoEwElRBI4cMSxBT7idahFoakfxYCg+cFD6a6myLCfFwIElIXqz6IjheQEYnza
3XKwUfHSorLyJsQHIZQ3IzD+vxjBzE3AgQZKO3mWVyLWvSIU2hjR4rJLpo0y/vNm9ZpUMTUNkVQz
T5Qy1TgVktmIzQGwsnTE/MckefiCxLi/oTm6ah7HFYNY1bZ8WluCPpEcPzMG2GsyQUL3wfVihHsY
gEb3J06Ex2HSvzHqTJOlmbKPW7M214sAJ16RHL/ODOk+AmXzqBkGJFiMQFuinqjqopAQ1qOJAlNL
SxD7iVwFhONmhF9jRaMJyXWu6jf/x+Z37pcUquvKwnbXkNBjwesz/3wK5hrDoGpk99sv1f1AGAGs
0YmOXnUnrw4lmGZFNQVEb3PSmiSiFMHEqh6LvDjkdBreNsMvYqCv9HCDGoj/N8nXZls1SCSH7awx
GKDjAZT5aLuww/6hxaTKKQLci7i+vKtM1ThHKjGztQpBCUYPYPjVw2GX6gCbyetQ3y7qnZpc1z1K
6J6PtGzF+xduJ3ZB//Qq08OAsFSnSIIjd8NqwTd7xLbvJC62OjHxsppdkL50rNnDEgbQtgGDIW3n
jpMvdbTRxJnbiYj1wEf2tgq1oPaWM7qbotr2b/rmtC75+G61PmP7FdKPftS/YomWjzoD3VhzEVci
b+VYG9Adsc5ohgE5lqWp4RsnKO/NkbzwLW+8q/qut9DbwQjIUU2B6u2XD4HlavcsDhDhPALuhMxf
X0s7cmn3FX6B24eQBv3wq7ubBw9OLbZyj/enxGjIHn/QWR72s0MojI2SngVysxuij9Y6KZYa7uVG
Hfhp+P6HROzjDKXEVDPftp+dZu3f8TH6nJD1/VP7fpJMrtmX5jY5vMqv8mHvIqhXbsOBnCEkBiiy
2MtcQ97G2Qdx0QMCMefaqYHBvnawddQDZERmzZAxMJqevkRidTi+uARuYUDi4cutCSuydxCtdleq
xjGgO+c3wZFiqV8bldZ3Bi/C0WSYTTZiITdf/OQDh2dg3XcmaROeximaSAyWrr223Ooq/uvg1mbB
RYayfhvda2dvlvwVrhmQEqotfn+GcgZgWX7yaDf2HSwRw442sMUnmLD9zE35d0V+ptNcAPPlph2/
MyFjEqsLhnGmjuyJC911iOfbU2BWrNiGnvFko4/yUSg29XGgRuQl21U1ZUrbUMSHhEWWIlMSIhWu
etLXosA3+kRS5Lk+U6Y6wqTpg2IvAT3WTsfxsG5eC1O6nszrjy9843tBgsofirRUD3s89mGDk7vU
hFaoVQQ2Swl0wFhDPzKQwYTgcvVm4QTHDMwdwWpu56D+p9u7DVVNZeaAiLig+FfVRgiIQq6WKRhC
3Irc+n4E5Ggys0lkFM9RVKXZoKR6Ul05RWTBj/mBmyrgcnw8BD/n7TDZ8G9CuCvs+HqWtuy2Yz7m
/sHYh+mf/q4Uz03aYtecIVIOX+IV8OXZ+f04jRJ+WtmymppBk1ygzo/GQifzyNM7cvzOf0Q6HNOL
IlNYQ8LFW4CEyqNkq75D3CkBwIjmhcqH76FMHMnyeAhmDsDqrpUkiH5nP819h2Z22tsbDIHW0TjA
BLWXzXtRAfrzcoHs7PZH+eg7UWv0ZBXia4tgNF3zLuyHVobeMEIjiUcdOEFwF/ROw4mF26fL2IH5
+5pLDuQqBj8z8OV6OcmjEyPGeTUOdgW34hgHR5nK+xXMtRd2sjsAPKhY+PFaR50wYUUwrHygyXWV
fUl+mbxVYBZgdlvLiSSrr76ua9oVnkDKOuk54xHH0t70xXyn9tun8jVjwsHrqge7kfQx+jPHt/uL
3h80Zx78nvml/Jey8bu4CGjVSU4n1NYFnydgve32CWYrVZRkQOT+h4dhnmPCN53uEO5811BKrb7T
4hPY3FQfdpZJGfoBPnvypUTwWqYtP6Fzo1GawX9HAqu105Wvqyf/JogGmP5smFmkVljO0zMUlV2Y
01/Tb1nRX5kmVZHZdY77KbRw9vbRyYsIEpCSV8PKZ0AeXY26gnAe4aUUVFtGK3SNkwVJ4YnHorYp
lZqdIMV1S209Of/uP/CnwhIsVJXjuw8InKSHXqdWBCDogl3ykeLSZrKAwA7CuWs6qNhUwA9GC1d3
LS6ejZ56jvqJKMCtsDb1Zw6I0tUUhpbeCd1Xkcdiz78vRt8NuwefEk1+dvBjrozxYtKf5HOtXM2g
VPbpMGdSvtfviAcmnSAK4aWbh4EgEWjuMWB1WXa1PLI7wTE6Dd5EwwOJPVzBGYoJ16fvkFV8+m78
VMWpfdp/SdYfPXBWGnOzbh/SEtY6jyhGT93NSRCEsbpmKaHKFMTvzyaGFUCYNonBbvRVmMDNn3Dp
v4u+cpl1utBYg6VDiT2HQr8UtNRJl3pZSxkJaArXGX7Vv9oNgn77kWtXXjrrmSXajfSfpkTZpTWn
/5Gz2FpMLHZhjP8uZbOKcBkUsRM8Bamd0SEJvWn2CYRgqaXizhORNX/r/r8eqxRi4Dm2n8J8LdrH
rga4lMwl3T2387WDLBG86jrAj6cw5OMVqbR1DV/SkmfP34+WofoHfkUa0wOJZwYHiMuh87uFQG2q
Z9hZngZP/9EbtIgfXFE9hes+9ymtfDzvjSN9oN7yI5efguj+y1O4Dk9flhZbGj3W8IZV7UDVWARM
r25bXgB3/4mIc0w1ePMoSYY0PJClMd2gUlYBy4GzPqxaHGsBOp6gC84849+vVr6BvQzjVQK1mAS7
QFaeGw8rH8rDMfHiv2dRhEEviUrwx9wE3SDbElcF2mwgTv+QwoXWAEK/vMfrd2Tb9ik03DiSCt4h
lg5Vs0YrK69sDD/etdH5PGjEorch9fHwCSEpEuNqy/txMLrzej6SnrEgrnesfM5qXHP2eH5E1dzf
tISRoGZzGOJa349CKweAM+SHW9vOXx6JTmHwASlQVmQJJOsvFDV+B/bbGxUH6O2/oCuycHvW6C72
OgPbayoqb494z/JI3B8BXaOlvBqOnwZsP0FE0PUDRAXgPqAb7kG7+l2foVWED5zWi2BfxrQz3pxY
3Y/4+IOwdYADSeB8YNb9Tly+wTybQFfiALzb+YySnoHfm5TLK4uxcLMj7D42aLFTnAkC3x7IhVLE
FfnQAGnV2pbEU4BntPdX1Dw3oYD3Lcm70uTCzMx3ZMchkm0kEaQ0iBLYoYTUKGmJam0pnjWfCDHO
pjmswmczqs+JaYjhiVDpeNG3Sb5aQNiUPvN09AdpQjkHKkaCfuUWyKqm7OWpKVE668LvJf6u6pop
V+/AA6/tWkkVg6RNeKSNwteD6Htjghi+Ke9kcZYBH2FnDXlwPapTivrqtp9cfRT2a/fHzWvlGK7/
sZPjD6+FsUTeM2BHBYWqCFMhPSR9KU7bucwsL+lNrmX9E8IbY8kXPkfiquXZkm4ffVeEiF/w0Z7T
pfUY8jlKTRdiMv5W+qY5lLkT6X33dkd8afTfeah4XyDFedPLpxw0AeOyo2yM24STbXJ1HLy9/IAh
66XIw4Jy2dWaHC9ID1Tky+PtDpLqGUkbg5k0j+8sNsmGYYfmJZKxR54ULw+cbeT9RremLdJWk7af
qHGbx6DG7bLLcKZSWXH4Atsx4AslP88BtK5/DapuFlgZUa7XZtlOLouExQQ2bzXdILjwPF/He5rX
hbZShtkl9wZjNs8aiOTKMdft0SQ+fBqlkqNuRTdRH6po66R4so33nYWInfPbbuu/Lk1Xn1cJiNWB
6onGNG9kIcxuG1e245LnumWadBW3V5SRNDnxhvs+LYlsv12KTWsUl/mJC26G/QwXYbumLt2ooKbs
9/sFBpS3fG08kB4Yamahi4L/TSSfG0Gsi2Tlz7UanEY6JLMSbC7gJRBLNIAdlQxqLwon8GELf3RT
tN5YEDvRC7b4hAiIisiLsXrgHBCmgBchG96AAIeEVpy8aC3ONXAyNfmomyvP0ExD26pad2+BIkiD
ewGH7wkmzNSWaOCqNUokQadZu07x1CDqWUpqLgBYF5qTMyu44eM/vZtfMs4QsQZCbq2vanEklCrF
Hb0fpBIzLCP9PZJFmbUHHViirU1ttq0DebOxYWiolBHyB7/Rc4KhXdCTozbuV36k/9PoMMxkIiZI
ymvsO0COr6/2q38PT+JAbTFI64fG187r3gBSu64RPU9NYJacI1X/kq7QXX4tMlTE40z2/Tt8DJyI
TAwn45fL+cDPC96OEU2UJTB+e7M7xvMUBn+7uLWcKXkqSNYGGVS2D5D85dlHsG+mCYPQUzFJykFh
yOm5++2fS8/2w98f3V3L0m01AlSpCoQ0GgHeyWbUtK6n0Nrgwkl2/9zh6j6hUmV2SG2n/rRpAr9S
RlB+B/Q0/h8KtD38IWbxBydNLe7tHN2F0+GkuRVqmeAXprYFJn7rks2lw3MtdDcmEafvq/QV8259
pch1RWH/zZJBXfRuDseGrFCKUBuOuzOM3ueFc6sJ+NAZHZf0vAHMi8gZ6kaR/v9crab+tbdolAbs
LmJwOGxgltz9R8Kn3wMjoaqt4uK9FM4HjTQudtzDYwuIEl1+cIacBcOtq1icPI0lrmd8IjqUbEWg
DHVM6gL9mj0PQuPnT1D2ni1nKJ00T6IiVR8ik2Z1AQGh9A5odFCIwTKBQsZbaNoeDxJb+TZXjPZm
kK6VsYSi2/Lfj7wOUpqPHckDIxBKTT7Kaz4KL3sy4aTRV/v54Di6NdfRDzXNj8syiZ1YJ7Noj6CV
9Ma+VSD7tmCSsWbOPdNIfmpU+/CFS2BW4rfhqO5EvljaNC2IRWdeLpD6Sq3aCY51h7F10Knd5TCM
g3s9AQ79nzVij3lziRrWc5QULrN9Mx8GCgKsYl0T+OqT9ZhWerX9LgWMEvi00feKk7WohUHN0tIT
paBbEYePwqd1GTcGc0iH1flghpYhGqqlgvdHGJ/Bhy8QakMtK4zv/vNU/gfyeXy4DOWsuhJUoKgo
Ld2xpWGP7i0D7bBMuuHWcivw+oL7HviZR+ore+OrtaiSsXw8GKY+nhnExPP0TMJ3tbx/DNU5EASl
W0eXsfSTn2C+1/wD4G7Ei/xsXTHW/aoplDainGuToaUKDXHGGWnlf5Cx3QzU4d2OrZoE/hwg2Bhu
Ph7HaQ5mgnY4J7YAxxFhJIpkWwNeA9uvxNYexugTFVMbDEcsJoNgkBYgaBoIYX3VArEHNcZcDqyc
25pTG5GaNfL1uoz3X37zbL2D+/9bvuBhLQ8YPb9xMdQvxV3USYf2lxBFScV51BFeOUeKVRT+rojt
UWXPnHR6tgXh8vVqiM0p29nkde3Oro4koha4S5MShTsgLJv9iG9htF7pt1oylKXpDTXwL0SBLoAk
d0fm/bYgVhNQ7b0JOm5PERTH8sV/l0ZHWq7PMgivGdHLIocMdr1zkXu5grDpd4OycvxrJERMzdF2
w8hnLbjDKaNc+PzDnIrztiH0/tDjpRVsj5vXeN7fAVNDjFpgCoxRNdc6fQ6oaA/Wx1sYuxdfcL5n
0H8Pi6sywdkNkf02r7H9DkRksesxO/2A1x4Ton7rmzH0r5yfeMdumhbDzgOURFF73lAw8liVImnX
G6Ys1XwYVUxKj4V27byGyVbtW62lRB82OYJmX4OZHwj2k2Heh82Sxxm5WuvmsAwbKMv5PgJ61ktK
tENlPLyZxOJnCU+6Bqka4RBxASLrn98tmF+AU5PnAJnVI+rBc04jz/xK5htLFpGc2VzxQB+wWeit
x+yv1FxuRbFtbecWx+aJby15PKU10tF4Jf+c+BuGoAnpuEtoLptmtLkyyVQlD2YXrpl8G6LeGV0G
60rJ5JOUBh/deDGpZi8VT32TSbfIftj6Qt5UJ0A4zm5cQZflB7x1MkZxiBADvuPZhYhth7ezZegX
+s52bsNOwVm1l3cBfP+jfzsoLujGtL4m77sRW+4lVdA8OWO7Y27sdwUwHkeyMbG6wFTUks4xggbr
NTaNR/s6SxtajbGd5VIiDgQOhfxQ5x6UFKydS5moywmF6I+Cz/ag7uV8nkCpdMw+3JK4OuQyuCNe
KF4bFke/2LgcbVFFTzBDVOpwPISyxThPyLxKExvUDiXmHb8JaLgVX06xKp1rZkBdhOhddIEf+ibK
51/o6MF+ka9GWtA8l3gR+TceD4vyfSdYLup1r+cB0DyQKD0qOwdDnCZkCD4hyUWvpnFGFpIhyeDd
AthkxGuhj4Qr5lRSE/TY5tD9dLDMCBlzTJvnrMX+lCj/StvsJ2aohTFhzJGfWPmmM4gG0SS+Utf1
c7WUSIJzIoqep6sVmmz05k4kBrPVCOE9N8lrwF5IcRDFJa1sFJkcDrmjndhGQJawDE6Dg9OLMGlO
fLGq8hwJ2OV7kUFywJBKomVU6qobDwBhu5kDHq6Ov/xostlfi/SiSCTwoTUjaZBnoJFxSbt5oIUA
fRSfWSDFtG/9QGmSOKlJQ28JTdy9SPTrShtMLMjsSPb7l7vicLlfOzgEnthELOUWyX1KbTWA9Bp8
kwFZYfFSocBGFsz/eSVLrvctsXvTuo4zKQ8V3k601Y7FQneoiLZXsf68kZmlyN+aPNnEFc5cTUQZ
YA1imTownAA3u35mVGd0vFRDuCHKjFwSY9KWpts33zqjbn8Vpsdk9gxX/0bOFzuCXx47RJzbNDKD
we1BEfIvCEg/Ap4tvZMQtbo7dPut84oUNWdZtlX/oN3u10j06SvKTz9l/GegTeIfqFbQNFuD4Ppz
mnATM7TwPktOqSd8akZJ0PSt1R5Yf7NWqYlwN98K/UzKm9rln5RET4OFAlYkW8BE98re3Z+ntYA7
ZKhDTiIvp9wbt6ei4ICZsJBgenwhLSkQ/lV/76wFGSTagoTjZnkm8VqH0VFjAlHky2TNagPVMCCn
dMFBpxT7AxANVP0RzxR4LiOY81cMRXKcfYrBSgyFpifZB1C/Rfw5nALTYl13NqtEJVts8SbKTmaj
5x4twI/SNg35S9/RVyhnpKFFOGfbFtfTeR4qTzKkoONJrq7pMMPFg/dwwsW9Ee0oubI5grzL8ll0
qFPXLK1IgmMsFOfttSdxUNxBJV/iIquUZCFv9Wa1o/xxfRy6F1CJ/4It0tGqQ2rf/UVf8Idaf/yR
0cjgrbD/JWC9PlKVowgZxtjs+XYHOtxbIVhvePUXVVtygM/2OprIHWj4UB+m+bY/mzlSju2oL4GX
tyAZMMYZl4fbeLLq8TKIqKxH2r5zQVcLWwfIDqo6A6+iuf0uqo4qP3zviDfawZQarC9eir3LTdKP
kv4e+iosSD+RzfcevER/i3CS8sy/znRnTWeGucBsWlrHgACYU7ur0qj21ru4k4B8b4oyAbnOAWIr
VZkZkU81QaLW6G0ZHodD808V6DGQa+t4CICx5FflqRS3IIP3mxZ/ehE975c0e5/GtEdyrvo5Z7Ig
r0vNFTJPEVZVtDNyoukF+ibOo4pvlJ6RAezsZy16So2ic7PXC+U5DYmggpm+3/NdexuCsUgoMVAJ
xVhKSqEmBbecg8fr3f6dNpIVbTDrHxrXZy8Me1trEfeq39KaUIv3Qqery4s3a03qSKeSTZzsHT/m
rb9Scf1SbuSzgM/cJVYrWRyzciRiKjtLvRg0EhIdHmj+Yg9HQyrRsIt/yqJM7XJO9C0LKlUPElpl
7/W6YmICAmXvycF+NSjXlv46enlBSNjukUUcU9076GdHtSAtCF5BDVb6bE8WSUWnVwJ5WW3VLd3B
AUyYiUPUoqXQx98Tctuq5BiLgDsKfZ4Yvs6MYTlx84NFCyiPvFNmQ+ikRiYl1qZ5EYjhogcwiPQr
5lkwQ0nG0P8MYim16krtn0FuID62OsCzc6nnKXM+deh6a7ShvglGHy1xfZjDotXI7SSehAFce57i
l//CKx/EDme/0xc4nklRpkG3hUsrFLhkR+75+WKWVZzuxmyX06P/j67B4ujBtHLACuBgQXT+7OZP
iCMJdJnJVK42eBJOUi1J1DfPp+1mnqGOAkR8mUpBY7G2B/bjGbCUVM8OorUoFiqHDIprXhdaPqiM
cUzHLSChwnBd96znvtpCULKdkN0b2KxAAlzebAqLBRn/leFScfXPkQfYiOjParXlCc+SAM3vD5E9
KyUtViovQ0TMosy0+YtyUSVcufzhv9Wd/10v0Zk+k8xAEMX18pfi/I9AxHEFes0PG7wPaP9Nq9i8
A3F0ftF9Bq97zao81AcbJYEhsyvngaejmZTs3Z7UFTUkWyMIohrgrAq97B61/MT7qFiVrcm8FxxK
oXU0W+/bQxj4J5QT7bKicCv/MYeVMuF4TAOLYQAYXqdRCCxH6/8b5IAxbMvndWlplAyWe2ET9Siq
rVpPYtDfk4XYZ9VxwFWj0rmp5sZ2y9/r16FNwwaOSWa7J791gyHvMh+aZsn2+sBZ2S9DHfnqyue+
bm4QoQ2WuaFryGQRL/FG/84m1JCbg2sIJHEUN8XAqYAPHUlbvzyOKhIZnOZzWbCLuD5hApWsQA0k
mIGZ+YTstflvM4wgFVeZtp4h0T1uKSAIDEhTXUliI9t8LIMPhzkV/4DIBNCwFWirrA3GGb/7DW/v
0AzaiNJnW81R6VLarlgUfslLG+Vua4BV/Cfoza7VVLpHA+Mhn0ZxBWsLnME4PU6ilaTikZJGbYim
vRZVytwj6AxeyfxT5L7tGH7idnjKGIYecABQBnoAM4S9ybxWzeKnBpSaRmVUOU6a5YR5uUQ45k//
5Dpntc6QjRKrh6ldO+bixiAM7fljff8reO0KPOzAWP5XCvuyTlammQMsAozIpRJ5bAM0PEdsckKB
07UOw7Xidq9ozPH3bl0mLRP0CeBvbDpnIySiSR0KazXQC7CQ4dbglPczogQ6G5tSX7Z5+OCKfxn/
6KITHUIPuHI8ghddsNI/C6r4M8E9A2iTk14ELPRxzHCherRcILrQTtZBffF8dpLXylWXXA1xUT4O
CAh8RLrmydP0g4QVRTuCJSuBxFcNCzh40vPLB9bpVU0DA+k3i0+/DvBysUeJdBwNime6FORUC0ah
evDzmfzTg0NbDyVP+L4S8b86q4ojo5/QTjKQesEte7wHHfwi/hsf/VTYjKV06aXu823mu4Z2MKpw
QWtroaYeUMM6eoYXuQMEs2C5q4NhQNxObNhiCNWunjDj0CuS5+iDDFm1X3f2XjNdFgMiHWJdvesR
6GOZ8tidvACZ1MLeiyPbEJcPH34NGN5cjLWb3SH9CZ0I/VfVBoJt+UmsiPNJc3EhHjJFp3F6XQRR
ujkvbPt2pKpRGW7m63MPBtP04cPGS0KFgzZK+GWK2NetsVPsNfwApIBK24EDdAP2OCf8RIPWCwBc
obHIjJzBBsdmauOnXER9FhIZ5AD9KE94ngNm9bkL/MVWlnfTIpUKXv3h6euFmM/d6LV36URAAucs
o7btheffk4WAqrFkg9ebOHda6qp4hK4ahYXMFtC4CMD6vHYAIQpCVYALZzRvdafXIMo6FDntEee2
YBZ5UhFUhBiV1kYLxwcBQ72bpL8C/lagqi1K+QXYqgjBLE/EBHzpvDbYwkgnZmy5iq7Wbwnnh6Jo
4r+awWfFLioCu3aLXFxKk4O/DzdEzTuAstXXR5ColOD8gcTNz1ZGTg9O3FZSeoc4MD0oR5iEHjwi
ijBBDRmW/oemqJsxvDKBvrYbkrZGlq9124UdLZEDgNJWu6zdU3y7FuGeAu/qOcNBI5MwlxiR1168
kDivgfYgD+N52Ur8Zj7Yn7eMUassTpYjsWjHaSRPA7CDK8Rnxh/6uJ8C7Lv8ZlpTBcxdt3EsVCVZ
8HBv5rMX8nXkMjkBzTIYkUuA+0sfVtevBBNB6nbJ8PFTbQ0gDu9GPwELTOt6k6W+wpmINkzFZsYI
HDhAdoYB3+NvOxM+sxsT3NE7qll90m7uy5eYaG4tCEg445Kh8xlUViX/tyRDhHEcpx4UFXe3EVWL
4flfkzhsmI9YlBV8Uf6Wfp+0ek5p4xcz/dvqkAQ/2eaQfSLv3hnKTGwv3zp6luJFizdd0qIgmXFb
FvqTFFtWYne9yBvZn+U5bZUB+Dk+X+ZkTs+Wfr0Shs43I+L0G7uMfzSaX8rmgtZXe+HGGaQfGx0i
gyyunH4MM9Pee1YGL6WRtTZlKzZfMvlYUetDqi8q66aOnvuogHlIuavqVuEFxXjX7Mb0CqLhddjv
kRtj3Qky1VQSHwzeq9P3/ErYbZ8QOXJ/VdbtkzwY1b2ZfsamFW0yohdxVbZL92gRTYXkJtGfhR0I
u8DU5sNnu9ehnl0FEtUNqEtebiZTUFISiJxGIfjmxM9T+QaEmoInArGS+u2T8LHrVByqecoKTmm4
yg13t7rlTjrmoJSCcjwQoI16afOF8iMF0WC4KPVkxvWx+JAb5v6CJOUahBV9DL0ersfBtBrlr1fp
n7fUk/6n7Kf893uDMaTnkMGFs6O4BIFhfdH2i/NAy7z7meysPUzSV7DFVX+It2UYJs+MHoESnRuw
9MSw0rXphWdyXb96gKM20WkpgyFBNokrU2AYpkzdB0Ze9Zyc/xflQGkqYOXHmTJjm08xgMcNZtP2
ToFXlJMnIZClg3DFe+sReQQxew+dwmm4hKeOBdmHgWwv8MXDQfSi4wA32S9EDwnZM75s+58IaAv4
pWIkyTv5cDLwxoAzIdCjL5c27X0mnob7JtX689bzvBVudKbCW7n1JDnOdfGc86ByaTo7GBbJa+gS
OlNmHvkWYLyKX2SxLcDPtwaphhV7JQk09sPHX/D3M4FTWZZmzLoPpZp+WRMClKVSTInq+PVU++iV
wkpfONQlDuNFZ8QxLAI3XC9o+StgCQBZhCmVEyCyoqrNoZToWuUCspTITZcKxpd76haPp4tKVAOo
iJfAvN+9AVMCPw2nuRYw+p2roQE/7Yyg1InKVJBG9mDw+/BuuxFyD5zLAirQUcIffXqcRss7ivNB
IkfQuDoipqyLurk9vA27y1UXkDRVAnzNhwGsCnfZ7QoBtB/9ZTxHcW0JFrMWx5JuvOseRDlOUb5r
QPQiaeNIBcZISPWPzxBiq+PX0b7BvQr3zTojp5Bo1k0IradCrytdtNaEL/OAyaOYp3krsrrZbPCg
EQRADxbFMhu2NyB0teLyYk+bn+2JVR7pPvJfSgGwokEeCF67k6QgIrobs7Aa9dtDZvpgDvGduTzf
7O3QvxrXwT2vrI+Uefc7P/zB2DB6O2c9x47FW3UiNqrKzOwqckDVYkQAkY9ageeeL4F+3vxOlYLN
LZM/MaauPF/6dW8GMxj3sm8p5/1Nqaw7w+YMsEQ5Z0pWqNvCMj5zy1gNo3V0haUSe4pEuMuPbkzy
e/yXt29VfV2ZQJgf1LUvzRWzYgf/y6u7GBXlde9phrjMQjs+31CKpbTJrjdw/KAqGRbcnbyAYmUH
Ez4vB4MlJnvNYuQiICxQe/kdcmyH4pHHXNFcG2RmOOcoAWF3KepUx8j5LmM8z62ZALLGpJ8hYUqr
nIUnB3IYNVmsjxcCyZ8GbzPbrNTKZTZiPFujonU1ol0zIfuqevc5yOdXpccQkdhh28/3FGfOo5IF
V1AAVD4CTuiZl03qJSEVpi68NuTegW7bBI7z4MPr9ZlXNHL+RYv9Fi80ZXEvQpdwHrhnhW/GBnVL
Cjzxde6fb+LvJubKDU9SrmtF7ztSo8Wx/XuIgSv8lJHjMXSD+mjsn/qwBN/ip9B8y+ylFX8u1UzK
gowVafK/4nu/jae3DDLX1PIRmlvtyZHTdS/dv3ObT2ag8pCQRdgbDY5FaeY0+ReU+5M6jovn4sx6
qXJEKche+w4ppdoWGKewr1yPuRWw1tSe9I1ZXJKhoa96GfpHPQkBiQVLMDrM/nNVlGH0FuY8bQty
KhLL5g/0qcs7kk2p8cGP6san8ftFmip+wZUvoo7altw0S6X7yam6jSCEYuKwCco+fF78r1fXhV8J
H0jKxkGeCUAuGfqqczKDYKqHwVFDsalgY5wPfeCcQ6Qzvj2+rW8gXcaQHOlyo8duS1beB0PZBoE7
Lyv8ZioypRy4ThNT1k3HdAhTjo6Ywc9KDprpvlL2VHY6isdK9XC+VlQ5zZbM+Fbn82T1n4W/hAJq
13N5yF1xKazlQumAXAOOvmrxe/LqYF65mXE2klw0Cv8mpDYH6KmznN/+ZTAx+Mk2M65Ulxf0Y5fP
YCZBufAKvRsi+C7l1rsCImpahzP7G9WAcSejHpC2gKJRk/dSudiP4Dzid4BENs53CY059hdl07d1
PGKM+Bai5SvdxeUOPkpnX+KlIv4uJhg6dB15B1rbfyXVRp8d6cP+FTKl7qfIgQd9FjctYxHtQFTs
c1w7HFMu38i4X81xVZSpq5eZw84BLrix/3orWQUf47ZH9fdnwKdF6dr4XThNtoJCxnm0CxIkFzGF
KmdUMO96q8qgz8wlQx2fNgzDUDxWRWqldFWsEdObtH9XOFJX7NsDu5uuBvvQnzYakxuh5mKNZDvb
+Kz7Suq6ybMwauP4zo/EOM5pGbaGXprtkrBMkID4mjOyIpunjnD7ahcRhdoB8cFjHtnPirvUv0NL
CCvc6h2Km/UBOlXdMaMO/WR9mV8Gov8cBJSB3hhwM2Q4eK9nstqnr0T8AGAZjOdi1I7F5LQsZvkj
KyovHh1RLGFZHWzhxaDQLxsUT0QSnQOqW7jfQ/XoJ/m2rva5nuIDWxxF0DrlG7E+2MRZYaA9j5Vg
sfquhp7txbOX8VBmN7gvzcjKW4+tcXYtT8+QOfFAUIjEukAejbOIsUzPAYqAIx3Z5wiQFy8QRZ/K
EHNspqo2flln0AyOnrpQwGCaEqG1ibVqs6J7/hNEuIh8LHMSPyQcVxjWa6KdebQc3ioWF0bHxwvq
CfTXpO7hjUGZlFctjtLfarw8E4jua5xaSsdlkUW3SFdpjKY63wfKWJuu2mA8JwTS1I69NhVAhahl
QHiTiSe0bhYE/hewulClOKl4IJVBbvI+TvD7FIeohZ4wxpK7m/9C33w2JisYyNNT2o9PFXNVHV8k
8+OGiNQ8QoF4lQuYzIfjgyrUXvFxsCmvK5OjhOOqFjMvZtF1CblrU4d/d2CJQPrtvU2vTxOY4t6N
UP5+GlaB/ME+2/CrVMMBnsO5265xf1NBzlnvKpC2Pzw1rU1PKaNBiS2POjdNzqQX4Nim4bNq07WD
ci10an606qx2iq5+MdFW5plgQfn67tVvQwHCCDx8M6OQ63LbTha8dMhkU086DJOYT3HKnsWG/9fK
vaFGUv43H6p9F1a0Xh4QfC3+9TEGOVZT5CinD007GdOuFo1QHA7hYcf5ep4DwvcVmSG3lc7SzUQm
9qyzVvv28RnalQYedzF+GDGO76B7XzpPugBaN0UXae53kFR5/6rxJeID5My9/cdNfTdWMs0WpZD4
3ZUM+6/MZlUKSEtsDYTtn+5m4NqvTkzIGlfGH8imBIOyrRXuW2ZVUtxfwAR/DcMGOLUOyINZkbOf
x/GrbhQAHspgcoxauTi2V2kQePyD+mN7znKAdPyPGS6cjy1F25y37QI8NaASV0wOv+4sjbpbujAa
K4tTBG4HRy181mNDKJ3yoRRWZCI125j1oFY74hp9rKnyyWXllWJweOBMm0t8slXJm+7ZrTrmkAi6
iOmAKxaWx6LDBpUoot3UaLfQ/gu4Pg20jVUSoEirh5uHPhd/8fhetKfkr7UbZoRShcIp8OdN7yAN
QzOwsn3aVnr0GUmLskYZt/INf6I6tWutMw8uTUTgsSWOrlZHcUCgnFvNkqWeM4jaQEiP+3fhM8Oi
1YTTi8YJPYhdjgmbRh9PouYywljJMZ13jw/yY9OG2tmTC0kSF3V0OLFFqodQX+NkDR6SGpBHj3iW
scFIJjKLpKxApDFDdCdnllP52FwuGs6x91DFKkowoGEV1fYvpgHwS6HMyiR2XvyV4YdPJvE/EyVR
GUuftJ1H2b+Uc3+noJLGeD5iArpJhRh4THh7OsG4EtShcqKU5TVAy3yn4qWVOclTkyz4y/YFtzGL
wNyuy8b3mubKY6H/EUiFma0oc1uQmCQ9r/0DWigHgZiZlM7jUTzWZH60Jwj/HBCKB2iv2aypzVF0
5SdND12Uz5iO4FeeB1D0D/Gfjq7jf9yOwtQYF3lpU/xmFqGfurMPOrcPwlGajXDI+1gPBv6QBXvM
0D6WQECvp1dcqIPdNmKxY50QSx0g4joRJL1w3n1OOk6XlC9dyjHeL0wLAxxH2ZMnl4EupLD34zqi
lw7VxfvDVbGBPjxpq+esAq2yCqbtTM1CA64ldTRs5WEOOB0JkFahdc1Az66qpM3wCB4gVz6wpOJW
4HQhRgtK8eUqjM/GTiTDPk3hoWVYFrzwco7Z03snWjGKbbQ/5/Ro1eZGSyRLrbBJUduiBQM3DezD
uuz9/Yl0JuEQcOi68cFXOXp65+Ilfy8h34PWq2QV1WYB6Ghvz+LGCN8qMGRXxQXFawnDtmEKjH1Q
PB7a2pcBlHLs6CSKRIG+YBEdUSb/dKkAJr5PDQYzsji2/agC6bn6BiT0LfKIsulAGIC2HHPGT+eC
23iye1UgJDuIzrZ2pxsCvQLQrUc6HTnLbwjC9fv4kSdOjbpFWm5qmiV0jS56DknSPrwoE8HQaATG
5/YSyuJ7Kq5r6jooUhgKCS7WUcyF7mUhnGn4J9Pck3rZ/86pFt/Ftf+mVsTxY42C4k3sM671ZN6u
8cYiAfXM+Bi/84Y1qiOxK9LVnJRktmjhfs38+5se4OMOiLZ+mEX2jMT/ztF4WOy0Mu7Yl2TWydBq
j6syWzR1zNXH9CLb3HIUZ1EOLcDSlq4ktMLPab8vqMuhj4d9Lo6rkfKbXYasiL55VqNPchEkUt/j
N+XeVkXBumwIliDy+1r/oKqTAh6YoK+PU1Ha++naNKrHVqZl4Ubx+xWpR8DH6s35CKbhMJcwpcpn
DhwxFvsDu618VIWKP1W7S/CJcVZA28qER4XfdKBxFLx+x5rKt2nLKP/28O42fja2vk+yvWkPaFwZ
ErarDwV0H379HigdS99eNnKLcqPNabbq6YC80xMzOCH/FNzURf4tO0hlmp3ou7b1vejIabceQv+o
jUyOoKEajauZARFU67HlzfB0xCuoMmb0blXEKsivlLcBLY9LKKTtBS+eyaQgxMsaTBoP427TnsJh
Bi+KG91i0FuWqXZI59RbbqiVz4AkFq+F5l/Qfdg7eqQlwk1ljnf+A4k2zDonpa/f75WQSa7Jt6OU
gQm/LQiyqDqvZOuDnzSfLEH5C9vAdcS4WQfOhpVz7n9Cr/+Hf/qFmFDzgOGCI78Dvb12VBlUsWyV
Et4PeJ+nD2TWethrqCrNWYC/eZscjaFqyC76hIGCLffmvpEPJbZEVFlIaDol+axb6l4AguXdtRS1
y7aRPdco0O3Bjhl3oWyHXWGXuu04uW3RvCqnOHEp5f6iR68E4ulIsGfHnQnjfTXznHG27h17mthU
6/FGGm5iIVT1u6rYHiyA5OLL4+SuMrriE1lZt12XN1EwKMbgr6gBGOMCWVhT5GvmLr2KOTYG0iBB
6EvjX3rtlOKPw/mozuRmbDG05HX8QMiajxm64Oe+oW6Ky4C/whJCJcJmnCDcygpZA6JR8WOL1Gsm
7zJ+S6L0L8QTt5RLy0G9e6/Hxr4PjTqYlWKboxkLVxEJ1kJfdGoPXwVO93A5RIgC9UtVTV3FKyyG
fXxcAKIdstE8tWmppjqE26wC9ohGmkptZ4q7r6MLDg8hMtwtNV3R5qpPu3WG/GlJjQ7Z8o4S/XnZ
NwRvdtPVMGCPH4NK9lN4muz6B7BUp6wZTbBdB9jjme6szELyWTOGWa+qHKGLfI8Gl6RQhfs+5p2k
c4x34zjt58625YnVXYWpfKdrcNNwt+KUnow8yNnV7wE4b5q2OPNE2eGjlEU7MzkgzfWMVsUpiTMs
P3lxeOGtQt7FhepGwOpOJkwcgFgscJxR9BO02xEM5YSXNtOd02f++nzHjSqKzxBxRpCqO9qe5O3d
vp70kBOAUowO5PL8pn/xNx9lyOKUb5m2DasdGvrpvr+Q8lUg+x31R6Wf/wMtldXydLM/alhpryQ9
m6L+w4etTA0JouiUk7a+0g0JBwJM2vEkysg+V+ammqeTxzCA/S26sq5jbHaNKv9ZuKI64D1M3SzT
UosxthOWm9daATiN/DGcEezDzppIz6I2OUbEG4kDA4vFZCTg/UB875NrbOEnz0E/AIjpDTRSqLn1
KNf+VmgMpasNER7ZENzYJyqWT/4TUwt2qdg+igjiKdIrM6YwMorzHVfgavUorTbUNj/pW4dE38hj
To3mlOlwHPrGRiZKr7zPZOdPOnMqdVSeuiCg2IIVZFc4Qefpg5aElJIf8AKU6r2rLECKBkuvewJu
zrfunWRitqZunwj8fS17l6ISUri4UObESmhkS75/rve2hiBmQZRGvyq9KyC1Du61HDzuvXvvVsCX
5SvZ2ij28av1KURBmkslWk+84P7JjPJSEdO0rPOAGu5H9f4vMMJaQrwq0VQLSvlSmNtdwUQRskWO
oBuYx7uj9pYoq6y7ZUJ1VH6SfOzpZRvEKkZ/41f0d2/v4ItMn/HrKOdy+sToD76V6DvbUY7t5pwe
UFQs+xhXzZaSXXSRMKAUh8MBKqzQlPHGLOVjnilDxQ2xriovtNgT5nbB79ZJhsnyx1uUYGO+aBXD
Q7h5FKWpRVXSwajv0WzcNk32bitfpE9Wk5GvBCW+tediQuzRQnQJiiTo4zHlHRowu//p+yn97mL0
9wxdAampldXIsL+F9WOZ4nVy2i72QmKp2uUukaB7so41yaceuzIONS+CQKK8IpUSzC0t4X3OP76L
vky+7mFi5fcqcRxMlDfM71xpG55NMwMG0D6VBaHX29DRvysc7sF9XRwb3Hrb6obybAvV+7jNpbO9
F40psnjmPDOHiuTIqr55fqvCy+rMHVyGdt+MxqmpkeA+ZJ5Tu5LITw6dOVXUEva72bFpGSDuB2Mp
Ec0FN3AeJGLe78VzX2AHn/wpLNdVliCM/l8vFX9sdBpUnOQ28t2O6YbYi/kkpyPi7nuPAR9KdzcW
uaAoI9UMrqER8y0ZGpJFXCC7RwtolYpTld4A4PqAupCVFtA4Zq25PJPMJW+dUVQnH9vjiEqzCZDa
uAF+ZGbVelxczOBEyN32UzbN4/YkLSs7Eq6Y/OJYoTDqyaSCJPzagwANw5osXHDkAJ1IB/HpOGeB
R9JjYQlaa9dV9W+/3Zcla7kf2Nb5vD8pIo+Y0/GkaUvWy0BP9R0pcrECFWLmn/PScLWbrHnEtkPg
hfP7305nJrt25FQPaMQd4J+sgcXEZDQkUH+HoRvGOjIfOj+87S0ifqusDcRBT6ROFIrEcc7O6T7s
zSN4Hny6DikSU4r/CPFm4pLsazM4BEkOSTpwQ5z9xeHaYkM7HfISuf82jmVx1sSTQU8oGuGENco0
/WRaaRnqD0BvMFZDNfKODaQR6yo6+xHHll6UHLlC3GIHLNWayeVTYfxd6tOkG9FhxJkKwVyjap4n
8OhIraoh35cdO4zj6Rlyh8di2P1bX0++yJ9EdiJjr3IQj+e2p5ngG3KQ0rwUTBbjgspedw4+XUFc
hO8G4EHVnWxS6ZS5g+pyNuhl2qrH4iGrOJPiE2HoRswUttmYi4CrB51itAgWmo1MHH7IMxhPwykK
c1dx8eAicYggWd08n6UgFiYGRMlxCNuTGwXlTjQJCYi1eE+A2v3rhSIciHLEx+1MpK1+oCRQYFcN
7sRc6Rxq2fK1mWkEKZBGjwW/NbPzy1EH3Qot+IYhXEsGJnIcn+s2VJ3FiBEqhBrEp2yOLCt/4FRv
2YonsRoKOLOJ5uHba5RM4sFnJWruTntO0knb/z/ugMHxw0wV9IQKzwI60Bn7SS+H8ROuf36Ffhjr
iUExtKe3uf+LrrTnGMfJjkpKzseXfQRnaTIsNUjokZTaR8wDL4K1g0kZsyDqQ6Y6LY0atgLz6hbY
Ru1q4hWMVHKQncTos/CFG/C00w5dqAO9AtX0OspBczdrn9pWFS+SAN4bDp10BSbjBgtSwu+fwoF3
qCuQYftg1AlQY3NbJblh/8cuqUMeZD1+7kQNMRjwyrho+8l1Z+QFMDazQuPt2Oojvmw1knqczfcw
RpFnt6nisDNt3rY3QT2nSC5SWNB3D/anfJd4m2J/6Eo4hygcG5NnVB/Wuy0kmcsqNgS22YAJZkcT
VcB3PvTWVIvGyarWcmBLzNlQaAyxCGIIVsd2Ap4v9dIrmMXX9YezX9R1p52poXxLsjTpZq8LqC3j
yE0TPXjJ/YKnfzozQgixDhezxArnT8aSypkMrbEmAh9nGlIMm6fNHBm8yq/5p7Ss3rEndiorDDFl
cXaAtfSQdqK+Wo0anFqdCuBDVlRKn4Yr0bITwcilYgxG+Z4BNPwNiqVt0K356Kgolgne32ukqohX
jfky/gPvwq4raAETNExAUVCI9JW4NOM0+RXBWEAJMQKrSMCJKE00RU8YvXENM0HjUdmJfe4J8+LA
G3ScL9y3FjBwWtmqWB9hNxJ2VTq5NlVTV2q1UpEQkQjBQbqzjfBkn5Su8VwNmDwPAg/JhnG158fc
+GByzvdbb7AdJetWI9j0VyW58psyed1hQowam8THjLvxPKyPsYTIeHsivLTWjRGVTV0/MZnwHkXO
va5Bcxz3dN6vc8aI0LoIp90iYnzJWlHj2qB4AeriAd7dk+r4kZy0IpfzvJ4CLdHTuxORwROv9+LE
2VoJy1/+Ye6WHLZLAaBDu1wzQl4GYm9ewfWQ4gaD66z/spHTLAsxQAh6Gu9eHt9ku+isJx0NbMvS
5sf/Mit9Q/4agLf31P0k9hoCVAl3EhwGyrQRoDt+5bbInXOOMADfqrBWkgWt6Bou5/zIaFyh0JCS
rHNanBRs69xbD78CdUu5wrVTsm+IYMF43givgnwjMnWWfETKoXLjl0lNpf+MP2w8RAxj6hDchFbf
v8EMrM9IzOFJsrbnhq1BroKyVJ2K4jwJFYBwmSm2quX8FBxak99u5m5Qi5g5WwNdngjvuTC5zHJ4
3l7j+9ijIUPvDc6tk+WhCZTkCpF6iiUOwt4fkUC5qusIbRXaxYkWHXBCQX7wyGgpFkD85nOMKBtx
58Z/jKDNa2Ut/wjmCG/wPktaEBC+tCoR02juoTllYkE1wR0kTGfXeylQJ1ww8vjWx8bWXfKmT/Bn
B8sImFPhZbK7ug69PJYtWJzHVsWJLcirQ3PFcoFaoZfqbmyESH73+Cia6gxjvlzsaxBBD3AeFd9F
29t0w5+M1GdZBb9Patr2uHlQ2uTxkhVc3nNr3OrHSFVDnmrVg9+ZI56x7JfhRIGRG6yE8FSFKQJk
V/nbF76ysUe4YNwxKUldCo1ZNaarVjm/swOsuSuBiOqB/0BtIZaNoZ96g6ApF2aCgrGhl9NV9aUk
ix2g6nofGrsMCc0g7zP2X0Ia1GQdqslvMi9sb7RvVXBP9D6cX91Zm4Q6kJrF4YZkOtmLPJzKWkF+
rXgkmvYdkfVAsc4/jBSjB47gIeSfUmsb7ccyr1kEZaRYlY5srI7JZJ21H4m0L/tNvzgThZZitbSF
qYMvm5jUW3k15d+rKZrDMa4w6MwqToJOyqGgpjcrMeW1O80VQmZBBpz5Zj7aQUSvmTGULyhxbibu
IM77vpLKGHikjX8okY3/vnC60wfjYeDrp7mD+QbxcINeUfqntvhBE70irBgp7ng/SZNbXtkgvAU6
aFBzTBMBo1gWN6FgzyHPzEDLlfYzdZxjrmkbNWF1hsZDateApnQxAlAIk98EP2qoiSWjlCNEY388
ll7envGsl5MkNmwfkzotduDcxsi/H6fh4PhjaBVK2NUWtwrWNM6WaYhbc4BtsK4GZN+9IgfhoSm0
K+yUgsdfjv8cW02t0cQ4bfh5OJGFobIHLHC27DscwdoGCXX+mdmboPub2LPBE35ttn5YEiJFTT6v
Ryf90AZ5mGUDchLy30k37cxb2IhJLKuPq947/C5v8pue3+HaOHN2vUukW8jjgjpXWCmirUzKHmNX
w3pSM2b6l5Z9PY5OVldmV3uYp2ntkk6m4/pXo4uYBJhEH5CKYrwDHUccDsMD7EN+FPz3Dtta2x/3
9e8RA9lNDk25ng6wMcqx4g6uRaJOgcxXyq6cfVRs1JXwN05Ra0ORypv0hiRD4DdJSxiTcRCxxdPW
ItcLCiscvd+Bv/J0585N/PoJCPqqIz6JJxd2SXl2T8Fw8nvZ8m6tkXJmWm60g+AaVnfY1TMpEdre
3KqKXHgwgM+9FNgHdyPim0C+d+ACYCS/7XfEfI4eL3JHwUYesf/IkGFMblv8oOZ02UgHlEa8xMYS
I+D1gd4M4KAUzQMwZNFML19G9WgSjbD9CKgBM4EdbC9+1HOwSPmIwRE6yBkLh+2Fpsi53XreU1Rm
asN/bSHYZ4kTkFnSxsfF+IX+a+lVnDKppEeRn4B96A2ysJFAnVFRsNG7Qow8seWm5UCazsG5frxx
r6TZd3JGCBWFyVoCAg7776L+b/VnOrrC319+xJZltcFdlUpXuI1HSXm/KmpG8raracWv1OPIL2uF
j80vmu9nXQXYcaknpy+N2uqLWul/7COLZiaJXbXLroaEjZ0AMiiu+O2ryFIw2CJcctrIyYxuyfCo
pK0oDA2HlTzrCdZ0QVH/9tY7C2h4d1HQMGbzLkuF+vrQeG8kGSYT0zrLt3BTzoXmc5K6IVcmXpHn
XG5JKg0JOuBlQjXjUfxPB+dlscGd7WtdD4dJ8dOBbvg6vLWw/Y8lyWzN7oc7WT7olb+dFeAuRhCq
h9DmIKGL2xr/Pb5daZ0Iu3c4gdaRgvQS8yZevWywJEEStXm0y3RMAvrIamDfd0eHQD2C9k86ylz6
7qgybYsLLxwdUbiLynkDHKI1J6RfCk0uf122O9thg4Ca6Dv2Xdt/Q88OC6VUioKslfn0EuYVeLL8
cZpV/G6j61TlzeMIYgoo9dCEDPl+6vE8JRTnT7Ubq3CLnm7p7UgJAwLN1PAvQV0XfP0BlmUYEC6t
X5Yhr/HAi7xHsvDGYTVAJfFGisw6rz+UijyzAFE+mq+mid5O+OCH9+AEXbfmubEOw0BNANBWiLpQ
j/M9btknPoxAcqVzxTcaItBKCaWaukjgASJCSUzIUljILQTuNLFZeNY0JxXqiTOswmlXsuYFNqb5
WKfOKkHWMGKeoOkl5nqILlB0ExvAi7ETnTl1TW9329MH9/YVCkHNriytZCcH+bQDONnzTJHSsiSA
zSx7xA3t8PD5t8xfAlHewCyvSqm8qxljDeaM7Vp6cgLYEMW+K3HvUyiFDdtz+Be9LVQzFeOEq+Qi
fVTmJQp6Gk4KQZsO+qpoaxR224ezXOSD87QcJ1NuapfPPfHzP55SKt9s5Y34y2RCegHvuJHiuKHg
t7Q2YH9+GZvAHH0F7MFSO/qoyvpWCB3slxYy68wuaS2IL0q5ZytL9Ci+f4u+8qoj2rVe4y8ogoAh
MI1plaJiiSvHrm/hq+5nH/X6HXOKWpRsLf6JGt2e0q5Fe7GAj5gz4MlvOoxpQsQOZGOUT68ihtn7
VqgKSd0TNHYBeZLQgJdBZtLvK0t7l+5ngER+8rZi/70s1Ad27p54lawuuMgiKePYseFaWanbt1HM
BRqv5VlpVU4VIqV202lJcmb5ylgnhn9cyf1kb69jJyrmc9pzks0aNw+63SqCT4MUs80DWFbDOe4F
dOHnTOoXIq2lT9PpllqzJLzw6CrC+dhbW4VlwNqe8AqQcqa5VRIeiO/ckMpL8ui2RrWacUwQseEa
NsvwM3VX8U8A8zfWsnIpTZWbcenByoH4g3+2nN4zr6aruklhrvMpMiW+PofYWfaAOFcpYOtuwqBU
i0Tp3TXWMbHk36rV/X0LFkP4zIKkouqSCOuSvTTPFj19P66H3jHN6c9K6jWketO6fAiR7kY0fv+c
R+QeYB0LP9+zPITQ/i5gzytYNl8nOOesRDVmdYGE5gaYeUHdwHdUHWBRRAlTmDnKKBtLiq8R1KDA
8tDro0EdTS4Oq+1m04iIpQ/aRX1STgwuiqYygoOlWhsAw4zCYFfoOtUFIhpti6H+vCyimQnwxETc
h+BEIiN8yCbJRHTaSuRWmpfHnaG3AHB/xsR8uSWiX12wsCIUILIycpeiYdNbWUyq/5cPEjKrR+12
+fSg5CkUHVml2sf1sPeGZYYX87cbKpq1FK7IwAVHFaP9onkK9rSjB4ByEtSw8sVTqElU24OBf/4X
Mmfb4oDuXrxj/5deHMyz851fdQlUt0nue6WYxpDVaJVmnpxLi3yDYuSdwlUbN0AKJjkUPOgNhKhr
3yKCRasHcr8MAFo5vbOV7+jdnUQeStHX1OrCpS2AGiGhkbL4xwVqHdvgRreRql2VjicDJpjUPkoz
5rsqDd2+DEMff/6hyVzc69XtpiG9KE+XR1Rn3r5n5u5aktGbvGM2j5n+89SBSqK9ufFpKONH3sFe
cSkGpyg4Xkrl6Qg6Qw8xElwXig0KYEjfUVCwF77sfBjNk/HUIurXRPp6qMxANM6VKop9n2J/YEXx
TmJMARVEB7otNOmROhazeGY0DADXxFZVBZkdAYrA3E3jztnXV61YkHFzcNFZIzH2FuG4U8gVLhYW
fwEIOHnseO4GhDXn3Dql9128P8Eo3h4wQl/e5Up24o+UvqtU0p63QzZ825YOOa9VPdW3fYj2/4HE
yCXjucyFaeBZDP/5L+6juKUFegwkMDqFFPVmEiHBg7yg0RUafvzm+C07miVHW2uNKmTH985IbnCa
QZBuI+r2Y8C0RBHKqQDz4uPktf+yJHaLU1JEZ0Af3Gr/gE2LHDq790+QoP3V0PrvYJOKVMVf9RCN
C/qBSb0+usJcN81tmWc6G13az7T/WiTbLev6bj4kdiuivVatuI4HhOKnr2O/d/G++PDBb8uL7DIP
XAxbQVJqwrJ1uuJAEYiPhWJhWZuCnJYkIM6YvSvQ9uRq1ZrsyKvbtziAi1ubUKRbO4umA6mQTYta
ndoQmP3El4YJHfpoOcMZsl4+QfWcSsU1NC+m2BJlBo6WERTZByWRv1jMAOef4g31TcouracnZ7Km
1hQQIoeATACAHeojR4UVwg+CuFCqIsHEpGEck79N4DKo7MyZBWiiwIRjlpPaCmDx13QM34GsipeV
QIR0zRlq7IwTFiMPprlTz7pUvKKQNuLWgQV9eRpcCbF9KrRt2hAFXERrfinpx5CaYXPDW17N1dhB
KkejEV818ZG2+Gt7fsqD/fviV9N81HHa5jR9Yyo+Fe2A248+uS74HzZa3dPugarkoJH7HK9pww9M
hCivN+r38BUsW5mjlRqjQgpoFgY9B3CyYRrC2Ga4rjzHQaknpE/bNMLU0a2E5KuaEtFBgpCtVKp9
Dh/JCQoW22PPZ2zG1A+2tI2R31nNbIkKO7DdJMh/Iq8uh9sm0cLsUZbq72lehZUGnYuOQOFEwR7X
ahqOmU0jVz2g2ljiHwTcedhC4ne1HwF6kaEV5OWhxVvko5AKQs1BqdjPd9FRedEclelD51RiIwJQ
ZuuVpK4eiQbQWFDEho046LYENSgK3BoAXuIJ4VkIpGmZYkx59eyGFQ3Q5t6DGFdSGwI2C9qYoGGc
ae8jKnhbqnr/156/69WA1468fsLwC+5VFGw+RuCQleyA6os0rxVa6K5/XhN77aQExX6bSMO2khk3
T7anoM7alNzw/UO6JPVvCZS9+a0bjO11k/8V/Sj+HVgUr3CXNs6Iyx3/gqBtLsTeITWKOsDgk3ii
mQuwn31FZ0pZ5X5Kpi2VFGwtJRlMVKSUGeA4i9vKKsqTKzBaolCtjCq4ziyFMIwiRpM1YzqtbqCD
mseg+JuBkuE7LCcV5DC8H8JxDE52IwU7do7GVUg+bVGGkBNaM9rH0cSm5U1YGVkj0zoDBUgeyalR
NlHxIHybvbLioqtxAREBgatv4EKyPSTFv9zoRzARrWrcwR6MUKllk5yhlRoPglUZzS3PHYBuyinm
UQEJ84tfr1qc6d+Kl4vP9XLkYoZqUoD4lykrYphULkGjHjs6cECaqJEbk8GfvtOi/8gEm3czmnm2
yybV2q/CkuHQPZCwzssxAHtl8bu31Y//vCM8VvjcQ0zqfxULzdXQom5Yei+nILYQUkzMLrbTSsl3
+a1CdCpJJrbWxyRIISnZ1MPIdXSgUbrizzkVi/826KPd9icY/2W0h9PsUoh5srlOsiwn1l1h5m+U
1JJuaDOXl1J28hLQjDw2A8j5yRtWJULYNkn4mrXKxguPeXA5FhPmNI23bQ2e2Dzg+JGqRLzl13NV
hRkR5uwLyAlUOap15P9D4ILR0fhJI07N+qVocxiAS++Hcuez4wlidSkQn63wE2xKF7hcx8t1NZWr
tt12Xa+wsH0sMfnK3K1WMsYJVqoqE4uvF9qI/EoGIj/zgJqm+4bt9VRBR+ffyh6/yKaFUYNCmkXu
QhV36Tk3yY+eYxcN2XalqZHoxhbw3jNa8MfhJ3rd1TRjvUo59NpLqFykNXWYbPe6inSnsXzpSJep
GA4C3rVe5Z16p12rEvPhKkFD9mkXcWT8VXn+qqT/RaWn0Dyol/1xvZfcuSyxgF+M/huHYXxd2sNR
ApTPBgNOPLSutnsc3FgSXHdxQv2e18iAcrPbXzUX43rPXlTOXXzdMu2Q3MEbrDyBpFXQ+46TCOBY
sXzKRGunN/9hzDUjNexhIqh3pdlX+H0xmZBYGguPxsO1JiqJLmtOw8FOs9rihiPD+NBhlxRwyXoe
bUXlFOngMfFZXYRK/2oV1mBAeLUpFPW4nPosEWZzJ2WtAAa3h6NCJr6pJKSxidtYFn4V4SRqHrhI
4u7Xq0vzmjfoCplV4HM42IvQM92SVcFBtxuJgC9GFnMtoOPJ59sGQAurG6DSHnKEhSP7/uucQ806
zWuUB6YWtBoPZ/nrue8tEiORGH2MAYjgDuCbF5Wy+zeXHyHSu69KNLEDkv49mVjn7HZFtfQLhT8x
GzkhgkyLmBCyi3Jm5gOmyz9T8J3/FJDuYQJs2Oyx1s/kbMrWOC1uQzOQqPi4yG2iX3tuLHUwmZVV
nK9UaulfeXUlabbdS+otmdCjtnBInBlld6v4+1/0DhUdCE7DrVAbCDsCLqc25KTqKzgCs4hZgdId
6hsTONYHVun4XEEQyqPObhFWqePsMLgHnJjOdNAorp5v616n8lS4qLZAPDdZz4MR888pGAW9e8o0
JuH1huGs/CNvd5vZAR1E1x1PhXTQqwRO/pSyoDKvW2dRQifK56m4hlNgE56PNcreA43ZPsFUANWJ
Era4LBPszGcX8yEZEYpcYmjLc+SiXJlqyXDoSIh1iw806pIEURhlFwigxNEsgv3z/Hyp8V8pcwEu
HLWSvIlR3VBFeipzjOShX6uMh2HYrhjIpw2TNbbQw9/NJfy2tr7c5Xzfv9qsy+ZGaAcU5ZzvuwQl
VnHLj9uW9XatOsA+nhCgcXDX0cu/JGMtDEghSkSmbgjoiP/1C0QcSEmIYQsU9dgav5YdjjokjgpK
kl7kC0UK6nrtticyHWduDei2BsbVCjIDG1sN5FbMEamfItSI3bWezuqmRD6LPUPxX0g5KQjMjqKw
nSqV4ePdH9QUiuODskOBwvi+e5k5QbNgTLYWULzNZwGUOa/Eb6Gty8aYGNrQto1udVzDC7oaRxDN
hKU1wHroBKyWGEszem5gJTqS7jV5fyR/RHKAklDVB2sB4jCfHxL9b+7cDYVMW6Gmfp5FEkrMWqgx
T3nlSP/KXpq/oGPWeUv8lQRrdJ/s0mPgK4ysue+GVGRr5hJroPu9Lf056EFNUrTogSndVATgXl48
fRIxoM1HazCihdUW0lhbxF6CRpORL2ran4WOkll/+JZfCKiWPbPIBBIhVFpEr72WTgAggVz4boYw
AbJLyhn3zyj8h7on9HkapRaRcch4XNbt2a4weHcAze9CsW2VfGrkXsV/9RdpNFiHWHoPc1B0PfZE
zSSGqOGxgozqaA+PSwyDGOqzjfKVmf1ixjO03W0qrrga6WZG/rQoy09D3vs5F2xJYd1Ki9F3QfxI
b2dBo8ik0aLBYm37sobXW2pZf0jT6DnT8RIbi3yZOPbLEMTwNHJKeIXpaSOipzTd4WSLIbGq6Jx9
A33pcZUIrWqd1Xo3uNekqjyiERPJxD2eDf0ZV9q5XaqFZGyFgzpKlit0X2JDD0jKQ8K/rq+Q8GKA
Nqqi5RBjNZLIe3yMnQszF9HhUHvtB4qbtctw7vXgP7U840ZMrw/s2kKTTBdHg/cy5Fb/6JtAbJlR
jhkTZh76wR4JlSg4fkmruoIfhOkplxx3Jwq2lBBJ/SgtH0LEE9BachB3oesAhT749t1bfqg9qzfM
035Z6mWJfmwgBAiLGUKKck/xsWAFxtFikmF3oS1U4AsEjQXkeXAamzXVWklHEfb0aIWH4ZKByJl9
Hcu68wOvf2XRG7nVfVODFnUGn5INLHC3M3Lo2DAFIP6fpTa+pyoO2LfMn0dNwa7l2jIiKugTWKFZ
NkW3lUOOq8zdMhbLYzCPHppmEttW2384imk2KWxRA/mIYV6kyzBL2+nF/0eyA/WSK+Ekx7gZST+p
mPmd4KI/BWvPkrCneYTV27M9ZXU+L/1mZf6zwZCTSqm68CmJga9AUlfuwolnBAmtc+ZXcA7xgZA6
zzJypYMdUu3ufDckebPRQtp0C7e1OjyBGO9Wz8BfRvkx+S6mBlI5W1I+ODC0kPCW2E5qOGMuorpX
wwbXPf0wxTnjsjKlSXi75P8lEZj55vtT2nA12H9YCEtfdwo+rKTGav5dU846X80OWJywG6S9klaL
MyfzQHITKmQcNV/z/TpsT4N02Ctd3BWxskOEhCVQ75ysJ9CpqyFFBH4Stqno/0Al8BmihxS8cMkz
k8JTVfd3vggNHbi1ANadu9/qWfPd2/J9iGaxYUQevKD58/OsLlyKNTrWVcMEYMpvnRmt8+a6QMvu
aL4L0gdHOoBKVwK0ipA3JRla1hkTOlYkdn+udLa0Ogteud9cy0hcRVZpNqAX7/l01EmMOWuqMn2D
wUNSucgwZjdjmopSv0X3xbcdP84t+c2L4fEOBoZp4FsgqAbzC4tYJOTIT21NfmA7E+LgaXpwuQaf
bhosE6UyWV38rLWxSkCuUO2CfTQ8bX/U0J8BeKdYDYFE/sNrUVOE4UcqSebXS0h7n3N1xtdBkTIy
x67eeup2o7gKS5CmoPhId3tq55Fj64q+R80JvHVJxoRPmyT4lmXcH8URzFRVIN6Y4I6CFbbiWIjd
BPrEIVwlX3IA/N4N0C/z/JhQ1Cn6JwDhEw4eEG5tn1cY4Q9pz0hg9voIMt2ZxRc9WM09p52DO37j
vUaQWLqvO/e9UIaB2xxC8vicsaWRcXrb6hYiR41k14Y/PLLigffs18Dtjb3bXMm8Hx7pmUPqgv02
AyEOAdDFXbPrjjv4zf0FCcQhYxJyuNTcCIZOXSEuQ1hDClGV3Qah1xpjfC2E5cBjxgh7IBR0rgaZ
8GEc47MeIGtBWsaNKhIge9Zmx+z8HWKJfsEQ0QfDgt9JBsb1XJEp+PwRiwU4Axjftdt110xrSbt+
qS517nddOgcp/npD06cAb1C2OLdLHPUpgZrnnEASkkv2yESxTHlgGR7LF6SzmvW6u5HXJFn/o9W/
uiW0+P2WwhB0pQrqB42dLA7nceCBUMErBCZzknedNrKUE7vOF0VGdLz5NMB6OLQaPrQxwUMpCd9F
I29tQxKDRsYRrXeMIx9uKo4VCoFshe2Q6nAFNRgo3P71fcZ+/x/FgMNM1e1qGDYwQ4D3Bn1j9MAF
MYz4y8HOF3EmrNv1PZwymrMl5tynTPMN/ch/JyYjwq5MRVZiA0AjNfCsUjeZbc+zcY8KhyhSqyeW
m+3rV8lw/gQhT2EHyxA2yYImCGinD7qM2UXFzekTMjNAl5Dd5EY26S/My+hiAFWzGFNRY0yWECfV
fBzx48hDqFBayzka3mpDuzb6+ZRlTPc1bgB4E4k+LXt2QC5SdpKjbZHcb4t+Yj64YzS5bpQxUr1q
DvxRl5Eirc9zqwU2babwC8blnToXa456erSLDM1jyCu1R9pJr/RnWQduEMQGCgc19S3pJhfLYoHD
ySdyuszYpz41Ert89UCLbTTPXFfPF/KzFtodVpO9MzezY0Z21WTUfKhsE4EexGJxqlU4C0v+J3lK
qeoFGtt6cqqTPuBcSZBFbGUYjtOrfnN46W2s8MT2JTaDo0GhjuKXTEV1gD5UY5bNgmjXwyjUHWou
aTyhxY63lYPnb3WSEF/mSfKH335zr4KZBqgDJt7hNLjZrqO1xkNqZYCugzlPc3bTkdyUvtV1QY7K
EOK7uuOSQXNLPhyAciycAm6P2qFxv9xM/HEDdvudcfH3U1OgBSf+vXFadezj56TYonucxbqsMtUL
GL4y2xNmBdxpK6CIvgkexE4KxSVFqOhwouRImiC4nB/5A6mgRkEEa3C9Bj0pYrG9LqQ8KWBnmmxo
1ucmNoXYLpoOK+EiVw6B8wD0J9D2SkgEk4CMGpuaGObFj+GGiqRTkA5cuDv6tMT2XwX79qSsmjPw
tyuivtFwko+2p08mi+VYbyYpmfeeccHEmF9qchi4rQjbamlAM9zPgDF4iqww3rwL2WS2EOkW4cEL
d/90/37TYa2ze59aXyypgjPPnv00ndQNZT3OgYdcYRwS2HQhHg67FiAjhkEuwW1ANr7QIF5PlAgc
CdBZ07Pbf2ExNPHw9Qzmx0xwULVvnx+NxLWPYoZ7Qh3wW3Fnd9BtpX1chiUdftRcMm5AW0jIrgGL
n1QxT+dG+9/mBRZkZ0rpXXhizv50V5abUWo34c5ZqM4UCk7ttKbqaOHOWWwZDApwo+3NzNfFbb6j
4JNGvk7VsAMmKHeCxKvvjB1v8o5TiLqzbZEIWCsqDq3LAAwUsHtPdYsM5KL7vjXjnwK28vp2jJPq
9NK+nPLZBWkH0KH62Ajbl4PePiXTE3R8x8kJbDIAlTXmfjtXPXjkJZ8bgOx8HNug4DR70xkF93yi
NSHkByEVJ52HctvRgPeXbmzgAanN9RNqrK8C6DYMeMq2JfND05DExU+HNrL3QowxqdkcyjziHm9q
7PbTtVHqf0x8ZK91hjHDRG/uPouw2Ynf9zbDQoA16sCTIwxtPE4jsifFtRKGqIQ8Y1SrthY/WWSh
BGHm09hlYZe9m/YcPC/V4I0pA/frAiq0BKNbfWfJCrL54vTI24CTyL5dVaPcImiHJW9YzENzZy9P
Lt7rS4HIgNG3zD8AYCEnBsa5aLrcvqaR3j2Cau5jJi9eHa0PvQq4tvxP9eQihRyiYCqkqMrU0duL
VW9AG0MpBcGssUMIJK2UK7RtM9suEAf9P8QMgxtc5uOhfDD7jUfrmzQhWNxcF+a6RH8LYTqwwBOT
HSwfPEDupZz0iAWopSJhGRDQ9mBHA1ztWD69RvAf1WVc6CV0Cbmow2leH/RRRqrN223PaqLBM3Lb
DjvdZN6xj2fkLibiS/6QBSBqy7OZKHlvV4X+Q/Kg7VzY9ONIt4LcJiIEXxg/8YQ4aLZGWSWNp0uE
Xq3aRoJx616F/rw7QtSMWFcWGqX5064kzsUMnqehJnXS6sLkma4NvjqZbOcvbTg88N50YDyGq0hm
HKbGQhLYfbaJJy/JNlFZ4R+FX0ZgjW4ylqsyP6hubU36mquwhNBJY8jf9qxtRkJ2Hv6FKcTpaVtW
W1ItQFDgslFDEOSd3xMpqYrfllXkg68Fg8+eY1f8t/bnStVby/MSY0RBUjbYM1NtPLelbyQlrEaF
mifRkzTk051h/xxCroWRNzaRbxF6CjPGta27RxlZlVnStjEDdxfsU5eY2QwS/VYbaxOdOAEdoYYr
wpuxIcggDNj2EmRK0+18ZWkRj7UKlNKEOON6iKTRo3sBxd1BRV+iQ9GEfOgzTbyAAt+ufsSLbDj+
97U+7d+/xGpHyvURXhtZsoJ3I8SItTBVxMftp9IA44kGsxxa3vK12T5NWf5ETSggXBTFm9gBRrT/
V82tKs+F/D9Nys/CgUAheetkgEUtwE59vXF5fcd5F9j1ntqMklAcYIpf2lwGgoUPeTY9KRh8Ywex
/Ueg5LSfB8afk43DPJWx3V94UqFowK100TNLYWlvTRZwbo5Bypd1GGBztqau4Xu9AcLy1NVGJFcX
BmZieDlu/zhuEJxNod4KXydWLzprrlEOq8RO/naczi7eH90Bsf9YH5PYMQ5626Ng9IwcV+JcXERn
Zo5jj08HxMdnAXkeSKe5zW1f0T8rtPKlazGbCIlSwMjzFg6AjWHEhshFKvPkrTB4VTzmYsYuWk2C
N3OizVpe2O83OyfmweSU1wqKKebu4AAmM4hyC1Qxiult8tw5U39T7CvW/7tPrFjk939nc3L9PXIq
jmZ985QDhUS++mM6oFY6COGF56v+Me0jLoaC5b4WT/EG/smSf/maIXZ8eZ9vKA3vHcInILnUHCGP
o1bqYAjtD+eJZ8L8MWmE1ANikJli7ZV55hlGNnlvx2N+0xqQoub19s5Bpn8x6Lrxb0W3HWMXJGlE
ZjDtpVU/ZlDsjIhdMJkqjP0VTPI+pkFxgpjdr8zu3pAhWRRkTvXOxdFrIteLNPYZu/VGriEUNt9x
Le2MKzLeHJNOdPWrWTIwQOMLmKCexiwVQZDnfvI8V96tyK8lsdl0BHgVee2580tbR/VC/ikYbZuy
qO5wrxdnKfUpMGluuQzqKkhcINu7kqCR5Fj1UWz+On4DFCecYL3Bv1iEiuc5qP/8f/9j5NGGa0/W
CKrd1Ab9Oq/FsO9AfDBoSXWN5teIWy0VclEawGdp53EoAzgPEUvgBEehfRCEvxDLTak6GWT5FsAV
iqSlTeLQT7VM5er2YWc1VMV+PjL+7saJAXXjUUIAEJno/Ck2B9CTXJWoYqKNBzAKtlDR7pB7VfQA
v/7lGW0XrEqb9h0qv0kTFt8vR9XTMbgj2rX7VDeknXxzkB4Uth6RhYphQTHJVkxWLwK6cSqZP5ph
rmT7bp6mZxn+wyZDovNgVvXfYISl6yiIn4kvePwvbDonht9DfSeNCMrAaftyNTLmoue70bYHPOwd
FkcAt2BYvLv0sa7vz5yMcfwdPLti+f6hZJGhzE5g1jHJ4eTvuGz3r1QJu99LMDgZNdqgODRo+3WB
86P0s5zimTScgV96QyrEpLo1s6C+pq7wRLxc4qUVHYlUzSbQqRHMM3b8Uh7Cj9aMlQKdrrMwe/xg
irpJyxNJzFyku8rXb0nl3vqznTXfWipDFl8YY7q/0N+SZbjzsUPViHGNHFiZ/VdU5d65AeOaBA16
6sjGJboUoeNO9aOpthbTsTmOgCwBDrrQxk0mhcMwELLt3YRfTk3dKFlbk+2VtOC9iz9QUqsrVoRj
DTiYRf54zt+csVLeCAZtGCrh8W/RSPNyl8YYsuvcecqWS1mYQTaI7cugfFimqbxsFqUEH8I+FTtX
Y8Tx3xkrKgDZfFc7iboXlnB4K0dta407iQpZnZc3vezaYleg2Mx1eeuB7b+SMY3KtShEZPT/Eq3i
bmj9f35MRwcX7FlaxY0++IR/H1OVh3QiByTl7CnszF8TDFhU0qphkSuMHiYeeeMcfELcsj4BLnlp
iEj5FqaA20scpP5CsOhHY9lMtD1X4ZEdJMLEwNmJGb+uRr9ZlHoqwh4/oAL92ttV4bztRP60GXYA
YV/WNgORQsKmZjfp1XT9YNHgKXgE6gb1M4yzmIv1W/N2M+Q+Xh6tVVxqUB59NOR7tRsBqVRMAoe1
vv7tuPhJvwxtUn2uKjYo9CfOxzAs6QpQveQcH2UQGeypjkJbABpgHWp49vCQwh3DwVHrIC2AbdJZ
TQDffsWRScgX+Y2b8tZYDW81dZc3LK22ZV1DanBCJy98iEzYQMXrgTMiYDBKwLDAZLmSXanmVfIV
tTVTyUgvzdhF46lVsBjvMYPTQWPqJFkIK85/KQKwsYfP+B7IAMZ6yyyFY4O/lsvEBnwFQU0zvK0+
ubNigN6v8BBUGy5hBSJmjVuryaSB0ziW39B6TSGxbSXbpDMkHA70pFAhqLb7DoYgc4OqciUtPejS
p6HLcOlf89Nh8KNieC7bDPXkd9xiwWwH9PE7oMWN7SqD8zVfDVLlrADz/Hdy+8g8fjkR33ufg8fE
Zg7qnlRxZm/ySVMI2ykpqyHX1+aIwRNcbe91nUAjuBnORLUv+4X8F9DIrl7v9rvZVOhJTQiRMpgz
OZMK6dHIH6kEHmMQN15OMIcOndGz0Fn3S6/xAhUUTPH7szPEdmY101Z6GMVP5FROfy6ui1Eew1hD
hrHkbbsJGu4d/oqb8GWgzg503Gc5xqEK9cr5Yn8TlZkKqBQRdpP+ZvKBb9cHw2TUNahEAkTDQWYJ
Im8JFHozFAwHkoTiSpe8ZHG5yW0LBHPJ2Jf902Tx/HpCj9wUyfg1R+RZOeftYPESiNZOuzsbVRpz
55/zf8/QDUtlx3qq8o4Nn+Fo8DajRUvG96zY34+Bc9iE+vsUySjAaNpieZMgIbYDfEtTjEB3ZWr6
SluOqP5MWbm5v9CAiSvJXKgxdc9n8eGLrAGQfnDtxLZlUdu8RgeB+z+ylYPlObe6dj3XJw9BwA1B
dCvCLcsGbMhNBx/73XxfYYPLK0RjIdlzShgHOr7psrzNTP6Eoy4ylfLt82wQsEFHXIRzfshqBIsh
UcgUYc5uizinDDlmXpHTNp4CVrT7nynl/5gta74P3zrYb6PIp5a8Mjd6kHN/eAZhMOlpCdO46Dbp
kdYiaxNrPjOJrmA8U7wPaaOxzE4e8m8FTlf3MbhK5/yzpVOde4PBUkoO6n3C20526H9PhsgDD29E
UHjbjqHA2RCEZ/YGYO1e0h5/o3GGaq5CA5tNDSmiyg5KULv7fgmJO/9IESUaeYKFT1KghCRb9AQ5
J3E+Yd07svHffgxTdZtgHOv/Y5lhXBhjCWjjhU5Xgrp3brCJOhwpoTrMPzbMEFICzMQ81FndQ4rn
YxEcSd61AQNth5aTV0Wwp78vc6115yXFVr+hK8xsPcQIQYqfQuC8wg9oX+TZO5wfIMH2tQZV1+vA
hslVowFtXqvXyAW9Z6lBRM4nD2J6W2WEuUu5EQnaSXwJlEZXQ3pOoZWB4JIZ4GXZZxt46/bONlYi
SHGfr4MmrccvmI/USXW8hpvZ0tLA/d5OPwdj482kHUfQQoqRk6aBSEAIHBWUrsrVLqTNPD+K2obS
AlRPgmtu3MFPb/uycnm/YOkaXwZ13Ifh5ug2K9ZPBh+g2nmVdwghRlTRYl8ITBpyWW3IzHth0jGV
SuMHFs6dYUZxSVsBnes3WQbkEEdkIAwhajWHCy2g1DknkfSh/kKufNfgmX7byEbZYzUnI0XL7ajr
Z+OuBXL6SUccoo4wqASN0XnHp+O961t/nn5D5bLtoKoYZJpY2S0H0WuDuHnd5tT7zqdyiwjd532u
Y+mE+y2wAcTmfLJ7v6YXdiSJ5r5UrYU5BtMpynAOwYg8M/+OAQLpAZ+NSg+VMCzebs9ISCy+oEYU
zAGsRBXdTKiGS/4AuDATjLVFgieWxKYB7SHfKwrS6Vbb69ihHhLst87XMZFrzIGPb61/KRTtbVNM
XZ0F7Mm2KU7Ns5k+9wnQm+gYUstZd82QPnQpBqldS0zLXo+xcuQFA9hVo45Ps/6lzYRcbtELQPL+
EfPZQ6tFYvwjieRFLYvuyOIlM4ie3BuZBP178hO5JL8tpbr+juRBbDYYUSB0KYYoYVu6CCIpdW5O
LOFiIBMH/sBpxy0+hMwk9D64M41P/Z8JW1CHxStRNSc2BLN1+eRAp6LVnFvBvW9gr7M4RMkK6O/P
E4u41OXpxFQZKD0USat3U+hZctJx9ksqHj0j0EC1FUDHp0w8zQt42Yc37HzeDExGd266LnIyJ+vJ
isY3SU+pzY25uU9IhQbdLJPxweGiXh1Mw1EIHzE8i/7SNrIObSDt8b4fo7BSnea8IsPR5gR0bPr9
RSwP24OqYsAQIM8FdhbXXX7o9n/pQG6+l9oOE2i0OybAx0WVhKh91bue8PJNxBKff5aPAtqcj4Jw
tMXM3P4MAYJxXyi51APCunpmdbB3kh2NFNWdK+GQe0aDdN25i0LTXwTaLDkCHlYbIeH3yyiZI7L2
7YLg+mPJ6z/gWGIysPBMgno21J2dp9Qb71EFeFf7FU4JgKcHG9PdSj3nXRO/I2SE8fnbYRU9beDQ
vqc+algwE0P+TsbsXj3sxNP8S0ToyB1srvpvcT94jd1+GkAez585ds6aI1T/q3rhlfX8RFKWHVya
sKn/UVdj9PliQ6Mzv89qjRJ7NdWuCP0v6Ic6ACwHROKdbQobC0dugZEAh/XIbxc/m/dWvDLfTuiA
0AeQEsSM8LFWye2o9vCK3XBTEWOcFFtNN4fevyWEafkj//sVbEeOvytR+HFFNstM10nu5iJfAXqh
Maz3JeF1x/J98QfGJkIAT+OqbICzlWwcXte46oerkYzFk6aMr+63FOOCdGxedh4U7k/vCmiU+hDP
DIqd9LEfvWhO2Vx78KBHFaVYRF0+keUanQsD2tYDDRVMhAkFF1cbNEYfyhpWfH9ZsGHNow50H0Zv
uhpE1dTirHiisdqveSdXt31XSalKnoxsnL5qASkcdbgpNztSmKzt/opbgo0MuCIWtBhvgU57xudY
qphLWaETUnooqpGw6stldMCLtr8ql1/z80V3wSiMwUjcXCXfoFq96CbzaGgUkn9ZP9L26Gri8ten
4c+t63qpxi5VQErk7wS32E8dyTLdb6D6TMauuhA68vaxPhXZ4dlwvymYsfaHJquF2gXeFQHVUUfW
qViFcCcfum86ZTDcyTb0u1d/xxa3VuCm5nTsqDhbs+cKBUrwtSovdohbtgSB75d+IB/O6u+QWrQ5
FSxcxF/nIFj0Nkntk+mAgqkEJNptK7DHxOyw2zXrxGxOwNT5kkqfVpKJbzxcDqhJPbi1q1JjZ6Ev
rr/3pEfsLa2BrMK269Bfy3BIQT+sWlOD9LOHHM91Uj4XfHaYTU0QsHpRG/zn1KPn022z0jI+lmUt
2xVjiL//xsz6e9V2bVDbygZCBwM5M+1+/n7IzDo/rsD5JDjXJIjV68oueueNgjoy97cY3Dm/TaFl
kOvbDhrC/0hagwMb5TJ0lrC74jTmzqrHMmEp7xSOcQZ7gh6dQbDcSAZsuwLkayCp86LeIdH2Se6C
BXjMnXzsfBNqlsbBWEFX7xpQt+SIN2G7hm4fQq77e9GE5wnKF8YQzMcECG2fh7aVk2G9kbJlcSMF
03NgIdwB6aXG+OQdIeOLjO8c+KzcjWz+p3j0soecs8LRn63OSZv+eR1AjAOSB7WQsRpYWCKLGmzs
n32Os79mQkTP+i0RONQoUbKSaY4jf1lnYYwyT+GLJ/woMG+9xbk7W4AZZIcIEiOCDQIafOIMahBh
cVkRU/NGqXAybQQaq6Z+TkI4+rZ2gp1oesu2ad0jyzvlniaWUalw02oQdom3rqGEgVvV5PRTtkCY
v2YJdyJJUy0CoIn0p3PVAoyc0nDiPa+8u3OcL4U7lcGpWAYNDsoXMs+wsBwG+utXVyjd5v1BBObH
37JzIS5FU8YJ/ZINE+ufXm+JljLqIs3HnEC+vWJhf2ScUL+SyRZ50gXi3ImOGfZbcxGaA9vKN82Y
TBDAw+wmQD6WQme8MhZeUdSBG/bWXup2gj2sMr7enjkPQDZF4/2Vs0jsVzM6mLf5snsWspXhosT1
MdVTh3YHu0PF+cnnrsiOsYZm0RDgYZjY4RTs+Hv2vELfi/3i7NTJIjpCDbZ/teIc/K9wV11A9qg5
V41Iu6bmYpXbLq30/xQk9xJpDF1WbK3RT2fgX/BOZbml4OcfyHeHQDnVfD3T19cUfYqooE8d8fCF
akAvbq/qHuAlpg2HjH4uTTwNNGMgcNfndOkcorrFFA0gglILVh6YPWEuBmkEln7oRkMDXAcemT7t
DB44apxlLQeHYzcrpl0RE4GijeFdzEfmoQF/Kp1oqOIEEGDjYOZlKhf8L7NlM74ziFPvbgseVUkg
XT6w173of7zyIaEPovOZngmh32YI366X5/pb1v41SY53IQc8vEkClke2wRUhmIktW4Du4Ulat02P
a8frKyODE/XCpL8b1zDmJAf5F+5dD9SyrcQSX1gRAk8lEQcNyRoYQ24DTCmChFliY0L+fvqb/dL5
o0Fcp/+b8ElhH0/geZaTT9fECKzwsYKPULFrzgMIVDxnHqUTr0D3BZPymruIZRPcHa4V4cNLnBhp
dDartjGggYlgYahh1ak3ayxm3w3iqDAsiqmU6/PN5OrZMPz50BgNeww+qJ4PUmXUTiTxGoEqZIFg
9B0vfWl9aGHO8BBGlP5vp2bfYfwDpKq8xi7t66H2tYNtv5/r9qfj0+sZuVct9ktlR96Gj9nR5H5I
2207HA9t6nesEgW0CKFxcr/yPElxquUReis6xCo400qWf+2/hOnjwDobe1XCHTEgVZHa8dgbCgPo
N8hanPjDvbcLL6QL1PYJji/yFhUMabBetldpgMfgzs96ATURYXf/OoZhjEPUz83TTxD8gBj4x+gB
8qrvWWdPnQX+cpxzN9CiVRjoFBdO8GnT6OizZwunZWQzRIHe7CFegquN+YuEAEGzr+ydCuGiWve+
oSVNS60ToF0zunsMhJHKtKuORDbZBVCixwS3G2PAGK/2nQzeiiaCymPuMmz+nCmu8JFyJiTpbBne
cOH9IJ6is0KU9MV4DrywukRd0gNYXJ+LI7+gGlY10t314boCweX6RyW+vNoW+asKLtj8eoEAEQlS
5b6wdgKGDGJutB9ejTrp/J55ctLXxaTb++UMVuQOyAGNhmPNUHRFhKL/Dz/nk7rf5NJbSMLCCDBI
cl1eFhDC3PWOrL79MpKQQJW12ZH75nCKXZ6dkNcDpLEPXo/qADXkj7EMv65ZXqLALA50Tr58CHKr
CEa75MiX5Iuo/OtCOiDntSrwhxa+zDAQzLpPS7iUNkRwnCsgA6yw+/dXGgqOFdS8Ql9/FWwQML4E
TMoMpq1aT9/2QpVH2Hfy9VOd8breFRgq9Pf5wzblf3EAJlshHYs+auHue+YyFGwVCmJtiEEwIWXb
qphlnEYFobAaZ8muVYeNBMcax1nFUAEq86P4fWALBKI6BNeukDQELBmWT8ub0wk+4+7DYlpGzkCJ
Y4K77GJvJQPWqi8orX5W61pOKD2TsrSfeVDSPo7CGZFzyZgpbKyVpNcqnG9vz6CwyP/fE6s7KZh1
WYn/NLQm7nZeaDlKQrCVdDQQIhxRxaSD4nnig9fO9iDKLzqEp89FBPC+gy0xAMhwgtkVdAdvcM1J
wGFxyV5E0BX2T6aYS7uVzTcBcuRHt7or4llIu7UGyYcanJJ74lkwtjdKX+ldlLUQzLreZKou+xpz
aIDq0bdMDrtwdqiJt3Hd6KVLtDcZTGoEk5BPZ4D33X46BA5jE+t7jzpV9lnWGxOjXoAhPY7TQbi5
zF2gRzfcIBrxwOsThXfbgM+Fxo2IqQXqqzGusU1xrZ5tvuR9ley69vL2lZXTG+Gi6Bps8zHSoIek
1QscsT3FQC0NLhU9BTTkcMwENoml4KpizW7+AqrtqPxBkKs01wG7jN8v0nGIsWfWe4VoHqhiGZWb
EZt058ApS/VK4gZcjBf3+uDiEl5+6tZ/9H8KNtWTeEMiwZvmgW1rbeqAmDJwFyIAt1azh7zBRJWB
Q+h/MVdNBzly08kaPo7m3+EyvBhKSWLSna/Uss2fmhZ2dA89G9TqGOTZU5J7+sH8jQOHZ9n4RYhi
nWNvGPvF306gUOVG/Ywdd+860HfMb2SVTstxa9RX6l2NSwYkTXB/gNvxw54tn5gCQ/uSeZsLLnJg
p3sBiz/W6UEweH2eRvyu6wzXACG9BD1LVize3+tHRVk3uR4rkRo49B7l2yz0z//+Vb92BSweg//k
8JEUK+1t9yOsFzRK9NhdH8RME/MLtnf7eZmhOFO6rfVHGAKtFo9x5VwwXP48q1JjID/LkPtjDfto
+KLyar754GQzEeOmTBXUfnz0Bb8p2tGWw6Et5UhbGeg0XdIbFvrPmqKzkbYg7oCZLY67PMc2KVP/
rcMoOH057//lz7NHWVuTpQtzt3H5Oj2hmfBrBY6o7oayIERE1e6ZDzB+o69YGVALvgLM2A2ddqTa
msJi7bmj9qFqYehzL7hoOGHVoxs6kF+ITTGPVXoFOstPYIwLZp0WgRwYA18Te+ybZRA+waF9ARPe
ekGVW23kYWSZixYzCDnIn5egSlsznuciKP4hxrT8AT9K7aghLXk91TmaJh82msJ8nTvy7EZam2gA
GPtUmN5fSEoUYca3X0h4hJy3g70dxuXgR4anKpAoXbCJVo/uOoOJLA4KMXJkHCrukckGFt4RCGw+
ubcsFdkC+uC9t0f+s7bxY+DgtIO1Xks7plOL4TApmTruzZhA35Xz5vVLPo+PaXANlmZbrl6veThA
Pm1xaMjyFBZBqpe+1sRkcLevQdAXpL6i9yIOisoY97tA5+EyYl1ulY00zJ6l8GtOQv6mSiVrQ8uX
7lezd1igPU3QDOQ9Y9VbI9MnLgNCrtjaYSBumvcyNtdbPcdVsvqJde1D6XV20zycP8NTW4Yhbru+
qf0pYqt6UfIW2MpiH2/Sg1O3SyUPxJFZSyT5Mw6ZrXEkfe7BtKpnzA7fVtdhgY46UvFIlMFwcW3C
CDSP4F9v4xCWGsRIDRQwP9UQwE6m1nlIfQqKfKBc4Dw1FZc7gIGE4Lai3wwPwVZeMOOoyq4W2urs
zxdHGR5joha62nZMD07UpmzANkL6kALdxYpH18M120rb5nzh5c02HggQ3YcUyAXM+IFi+kIgK9zU
9GNPklp8mGQe7OkNVNe7in/c5HF6YC1SFtRohLIco4bXIWfDH/T73Q+YYiSaG7aevZJOxhAKJgMi
kc8AMoIKOwuNFSsGcllSbRvjCiXCoSgrC4feMXgLP6HIUFdXGxmznUO5xQK1le3dn4b07m2CmBy+
ZBVdVkWjiI2ZjpTnHaUliPfLW9YvFwu4lrK1HL5iALqfNz0G9uBATYqxw3/6TV/tTRPtgApB1T8m
RyYQI9hjwqIkfZYZO3b3OQO97c/wHvzXBBmpdM4WSTCuPp3+rvvoMISrItoXE0Hiu5eJ33iexIc/
4wDu0y7V88kuMl4lCQDhYOVs+j93m/WEOxUAk9VFw1420VreWFaKMh4HUCty7JnQST6kGjZWpJjR
XDm/ETUBABWc6GinZkEFKoMf40hbwt4ShQpApVVJyZWJ6yxilA3rl7I6S3cLWw8jIpIvB4B2uasu
+yfs8SJMuQsgxBu26FC/Ck5z+CZEHtQcQ6E/SendlNtatyTfet4O3tx5d2/6HdfWHFO2UqJ9WalH
uCB7nxht/MuDPyRnGraY9/VykU4SLQGeFuNKa09f7AKNVZblL5oo+b0+ktNZEf7B/aO5zSV9S62D
UrFetLDq9Zrrb0w/mVvgfQ50s97JuzHS/0YGugzX57vnTQvkcEVXqZTzGIo98/kzDqzyY+UY9ypr
z6P7mtyQtX7ed+SSiLJURS1I2jYvopIpnNhfXFlJUjwWdaZkQ/0GY9Vm5q4YLfLMeqnhZiRc5ibo
J9gH66V6sO2zKIox/Ue7DYv9oX5OpTWdVpkqOTojmnKxDCJddkGjl5qo13Mu7z3FfKZ3fh0TPdRZ
6klUd1MCvvGGXhz1nUAqIXdu2k2f2I/3Te50Gu1xTkosZlKf0+ubczQtv5Pk0L1aS5OHQFDvnpsI
s5ZX04YNhj3skKPNuHMmo5rMnOTU8yRPx9bD//FOBDRke89KEr0qAW5JjF+7r3QuGvERDsLZoMXt
4ATwz4A3BYb25yDYcer5ThhUdtHcNBos5K/+m/4Wc/pLUciZb886xFlUSP1/NdOD7eXGgYkpHboy
NuS/HFIdg4dIp6H3bRXZ0AqvgXl0sKYzPkUDmCeCiRN29/O9T86SsrYx94EzqDwDtjjNd7n/bWix
2EksbLuTWits6SZkG6Vs91ND9cwVC0HsBe9e4WgZkYciEco3WmO+e+lnBe4Z55/hjxxcRPKfhL+p
2INyONKBXjZ8ipawCHCZhDnV4ySfotb1mOGvtjGMhbTreNOvDt5kL+i+arl7oJF3/UeEBnPJv6Wo
RqipC3z90DRZAmlb/6OSYYIw6yaU/jNc1G71AS2wobq+OcOtpW7IZuLbJNv1+XjwnU3832lU5bdI
6ux+nUvJmGOz8re60kWPQI5ryv/vmMnlEbLhHtXAlEWvPN7jwkb2BSR8/52akiTg+hw89eD4w/qa
gz+RVsMoVFPST6E1qJvWsjxkCvLrzmI4/kWt32ESTAWrpoo/rs2lY4A1Tvk+OhNvEXGtiMNnXp0a
FT6VuQvE6HT2lzi2KYPRItkHAPZH5qUp7+a5OPp2+YNJrYjNggiB/TiIpGBhpLDXdojddLh/AoIx
jE2yD29OXmPpmWzHk+DEBRUB3nUNIDagS6gecLdyqjcxsb6qkzc1yvP4rPyAQcmmPX7mjaAuvOD3
fgHN0M+Y8UbMlEffvM0C3K7zj6zF5vsSRvQHPBQBEb8p3on29uKzoKpoP8SBOL1XDSO9hjNgrYQm
yyqYQHiiYdpXcNebivjSE4QfpqyzQvPJZyfy0EX4FxVW08KcThsNUcfZcsQzhqYXBTjUiocEPviK
eppOK6wbPJsTN+j8J+mpzXPYRcx9dQdcvOo8PvGp2WOk6ltSNHj0HuM8JLco2xYVNDhA2P5VDspm
+fWAze2ct8DAqPVMQyit5sDx61fKKuUq6o2A0H7WO+9VbafbKbWbfeNsKuRm4HX0uQmw19R8PQze
4SL68zEDNCDBzePA0dHHhDJKPLoPLJfBaPCQA/OvO3HTaTvPqr7LQSWsxksVs6Hfe8jq6HrS9802
mcAp+yoFcwdSr/HvLw9KMStTIfMP1WPaq4b94+SvQV+Smbc81pOgPH2rgtCGWX7adwS0r3NhWrHe
8wMEWRNKSCFdtL/vPOiXwWGcYXw+9JeEpH+OG/WRE3QgmiPQaSPgCyy+YtpNuBIFXjluoZNH7vVW
zk5gvle7Q/CQ2DKL0QPOtTCfGPu1AKNgss3eTKwLeKJL4aUZnxwZcUVguoFOLBjxk6glffAAqv1l
Ik6kn04WT16/XxPEfJDV7DaoH9VyjR85IhCk6ePolXNd8e9fnpB7PutruRnS4wA2yy7XZ2bqR0GS
i7hEbgyAe0Qemt78+s8hgpKVM36iAXQD833jjXSq5l+EspzFQRN+H4mmTS4UmzLNIQp8qUD9mdzs
5Z9CZXO8ayW/diFBIMuRuHC9SIoW4nfImpXJW1/LAarnbZND3vvECVZ5qeaHhyr1Q2Ig2bkrMZka
5uAMfPkOw7T6Aqi3e/JmEMScIe9ft4EdsjKQ/et1TfLbwz/GI7iSq6kaI66KPKVTBaF4VjKSTtpe
He7/NsQq6zSjh0TsCC1tGQLBvag4cR5V7jzE7ilaMqqmDrR8Gzb6x6hArLxQh1Xo5/eeWI2tk7cf
0PJbeQl7nxZV7pE4JIEAKuZ/sBZh/wqjnSCsSGcx/fCCsE7aiwXuPRPBsjC049u1TOJo0Kue/L5h
sTWLsvY5UlgmFTll7h7Ejx/D4CcgvK5BQ49AehphocPgjTYMpgVKIKrlc3gGekqOHCfO7WW43K05
Jc4QzVclESYKFbUgnJMP2za4tMVLgd/7/ShBc8UcKB7LDoELlhgA5TknE7oQa9u1xuq05PB+gmj3
EUYESY+3fhszC1fQSuB8K+JT2muE18brklPNBs6v7/8JkPxSjg1Q/MPYicfeBrMhm6c9/jqMYA0N
Wyk2ES04xnviCKn+VS3GRsBpJTIabAXjpPGqVPjPfOIFnTnITbCilWX3hmGw/vvrmv0IIwkJzBrX
6rye2bHvQvfFNKVR9+FxCedEe+KjH9g8SM6bHmtpVpE0/s+ND5mcyvUAZfBf82WGuK4kxoNVkcUK
E3cDtfXzjIQ7lH4F3WcOjaiCwpi8OOvLxMbNd3dENGQ0CVtfwKr5t59BFaWkb0CFI1LltSRbM/bd
3PsPHLR8ctMyVz5TFTwI4Tfxzd3ZBbvK8XIKyIWlqWyRYIBwTkyjRPXv4ktNBopIwB68j1G0sD+s
KXiODtU7Z7xcgjG0B7bDTplbsBI4sdLkfg/nMf5wcJkWDPZwd5TxnpkowqTEnIPq40n8qPzbN8ND
wdixk44MC8lrq1fpNHHKOlwSMBzy2X7Yak14J1UjAJVH5x0loO/yXzpP2JtNB+aPoZuN7t6SwTu4
O96Q0Gcyv/TvB0XxhfDiVk8W2k5mj/8XidMRcYmVm3biLSVXimszgxKCrzL+8r3HrsLzIliIbbSS
Q1F/K53GtVT0pxwKr2yPjcVS2slkBakbLyepGj8lh6FMgO3zUssWVpcCfHRUEJhS1G4lVsEP3vSn
hTvyBUPF/R9yciJGIyZNPkkWqGYlBoHJIZqUfMBq0gMpoN8RqKLfI/gg/6FZom3ScS9o3CIhG2Af
34EcYSylGNIOm5B7knkln16zfjr8Iu3c2PW/FzQyvxSPaYk+UqTAJ3tpTbpqbDQC6Ae1Lpyr137f
nAL+fjCMxOgMavUr0Q25WnH1cwcv7Dh1AlrwRzx+k8ZNJC/834xxbqrj9UAIBU5L9/RLi7emUsJM
flzteTxHwZKbPiSW5TynDNlrV3GUtO5SYnekJRKa/v2l+Ns+XI1sj7QuNJK4uKua+9ppKlyn0yk8
FzstPXcVav0qBqMTzAMIRDpaFi70kW9vzkiMDghPrQn1d+P4hrKwLTRIQ5D2bx1qUtBZsghfAf6S
Q7H3rI6zzYxQvOafDngqQcupqSNmP5bUCvYkJQeXqV9E9RR3LZ59QHZw+K2TejdwWatL8O6/WpvP
wHjiE3hgfua+r/hWUfxlZYwaNA8S/SnThTTPh0zW+YXKQAf6N0F1HD3jrskgN8fJ4T2etotnsv8H
sztddpsdywRr0Zcpu2iiRQaREdug1R2/Yiy5HUJHwALSPgdw0VnEsMUxPIYiEeLgEP9gE+8QFnH3
VOyAVR+pud1QFvMGxnXtxgK2B3W9nSCVWMfxzgI5xzwDFWuQHum9H9/MTEaNsBjH8fRTj+aGlMcP
MFC/iJgEPmFwNhSPHP+ycY7Gi33Epq+RTB6ZWyNvgckv52zBkytEvmuoMa+F+CmEP+kPl4SR3I9P
GTFhptn/n7zUjfD4DVkJFMKdg/JOBKSj4hsZXkCfd4TPiPL7gDGR7X7TAz7tVXMvjdz7hnk4eVki
G0DB9LXfbR4LO/+CjMaLAKztOzxxLQSZj+mn/mE9kQ3OmMoDasaQwmTVc6M4FmWvRUJhXndMYF6t
OD+RUfusMmMXCw/MG8qx2Y1l8oascCzbvYZPubfAd1tzQc3iL7pkggPjazP4rB2ru5P/pssgwhvx
Se4sj/Qo+AtbMVbquyfoaGddrXOGUhSjiOR8JpbwmS1T5jHuX1IrcjKaM3CfZ9f3IJ/sUw9Xp7Hc
pC67/LyOGxFH6dsk5W2fgF4r3pRCaL1mAZCZx0i+RCbqnSv3/WWhPy/3usUp84oxBYCLWm+68GgS
rGRmtRNqusEPj7MamfNMy93vcsn6JNYL05hjWXgQO8XRQMpzRMSHpGU8D9edKoflKfuHyDSIx0/F
NbxY6d2pYkEQqn2sunYB6TRhP4ZooZftlyyk4nQiaBV3u+Yn1izOOR2BTf/qjeHP+cf1YKvcE7Fq
cSsssIk5B4YusPaB/hovHqLbuWFB1HV052+aw/xz8N91s5ppcTJ261dr78m2x0SAbdAXu8JxNC+u
dpgZX1BZilTDvbca8duZParIOyryyvp8hGX8ya9eZbbNeGTE7OatDWbOcv8lZhULrKcGhNx9/Wfh
9Vd+OQMVI3E4FXgBt1+isjylaV9wX6mWVCfTOjoybZMswJDj3AeL+64HBn/rzeKmLng58wok2EU1
cSjnBd2qB8Guz1sTuguzTfcHbZ8NODWDfekC+qQ4QGZz97D8W6Qgs++YZi1lSUZnfIiEYIq6RzDB
m2jtUh7W1fUVQr/g15P15wLV35WYZDF6D99Sx/4FvI7mWDUqjfTOJSl93FzCi9E6kJU5d8FdIgRN
/9xyBHL7hS/bj4Hbj4Vdbe4inwfObAc1MzsxGuGEsuAR3q3iZfvqfoDyQF58yRsxx+tFqWe45YWV
fqfYsRppERp91I/zvw0dOAsOzUWrAAJCNnDUlqLNkjhpqurGvsayneFr8T6SvybvXUm/i6BsytI/
7USFPtPeagFnJqlUzJ6VJrtFEScQzSVV9QwkfYtlCQJtyYZIQzNfESBuoBx+TvFo+I+zkGh11So2
6v9j+uSWhGk7CFMJ38Q5bgUTp136X7mixcfYKhp4FYoWsksg8lROu7QcOujongrI4riBOMlIvsih
BX6N/06FrZnQWqjTIZIpE33yu23P/ZlQ1Gq4UMnfqygJ4XUQMcmoxLAnMBFXkR0omQMosgqLzOkc
FCErCH7ctTrioLijQb4Ikf/E9S63kpmvEeG3etCq3LLS2Iv9ERX0UIzWGhNJ1nfsIbWqL4/O6WE0
tsJ3RQPhn8zyjNU828X/Cm2RlcOq2mqLA/Xxlp6DA2ElM+4w8B8vy/6hCN+CKgavMVsynCBtqU/V
J99gBVP6GfmB2TeEN41joU4smSaw6P5v3yuiJqGbbfQt/Oujxh0m2BDEs2dErSTlEZIo2qD81VlA
zYNILucoBigNhKUEQYWe1abcRYu6Rz+mRTaYc1XGogXtE5YLcqWoqpKhg6pVepGBD5bi0Igbtkz6
agomrxhCE0No9+PSZK0V7reauziamBezBxg1jJo9aoBxsJxKH8Z+m89EbPYAJs+/6AZ33wL6WFuF
F5wvpnJvunTJtkfe4/P5neatL2D0syVbkDa1jOknoqr8bhbuvRMhLEWS4aSbF28g/lkR0tBVn/74
pZcTfwu5cYcFNaKVeJYREdCtFMye0+YPA/1YFHo7w2MGYijYGvnbzyHqkXOgsl/EHVyPc0SNPH2i
EvfvLaqxn4JNnEGFBaN+kVahUtr5nDLjkqFsGPKqCC66XivzibIPraaOmV5SoEu8tPVVF+nYXAXA
NWsnz4ds4D9BQ+vP4rUi2lAJwVmNw+JCLtjV+UE2/6bSHlua+2vfLyqIZ/Xn903Ru8xm6Ol0KdyA
Tg/l+kTElhkv4Vb50fBb9ptO9HMjYBruKUymgDWhzXS5YP9h93k7ZEqZbCG5wcg0vP7WQ4/HM7Qc
t15xbybBX+BS4ityyFUzjJObQB2ebAIQW0xfTOBDgJA8l/k8WMo7R2vqdg90TOfM2DuXpS21rIxu
cUJv4ugQmSgP7LH2754iOG5WEgrJJIjBSBcvocPkVEqKrGmvoobSmnGa5jsPSibxzXlWlf9t4KS0
NmvaMq8aI0+ZnCk+hSNVf6t4WcricuGPCfipOhW1slN7mfjaqwihlFHZ/NCHMZBVL24fslehNyG6
w3Gd9k9HatM0GDSvBI8bPUhfU/bjL+l0Q5Jnz37DaNhHj5T0aDu+Nt8xH0Cw16E/hDykCQ17spKf
oxbNVRLW1Cak26oneQ5i2NctDgJyThJXUt97FdBB0DURIe74W+baYJfnENpd/Xm5pGmDVy66lvat
BvW1RmtGP8kYJeSF938XD5+7vooCrmrkz106ZAS+NVdOd44v5zxYl2u73er6W0K3oKq6EMBzgcwx
e0dyRaDr3BwkIsOOsAIJq2km0mKvHD4TTme4Kye0QLpsircOSk7ISFo6gFfA/ZM8xX7g6QPN7yIL
KHctv5y7f2Prg7X5nVtTBsWb9Z8GGMvzrlt9WpZ8rNSSrjiF6LgcKw8VX80hZKqoGX/MLdK58818
lahY/+SbWlOi5wUDPU/k8Qj330MystTkuqeTfocsSCO4GXW3dKQ4hMvX8ZhGUsCINMo1bZTl7qh5
Re3/SiPijUVFo0OcE+ivntaq1d3/qSQujAnhLIK/neMZMhdCxt202GTrRQ/f2N2EQXWe0QmF7nJV
qYdY7RPGmPR3W0B8jnfKQXy3Po2nYEURJbtYW4V2lwmxYPB5I2Q73yDqydCeJnN3WKYacjVMGcLv
B6zr9Ccahwu2o/8cYawZAE6ICLsq4JGXrC4JrBwbdaoGofZlWcfaj3s9BzOg4RuFK+Ql+f55bYKY
n8lsYcjyjQmi8UcxXkLa+wvZu7eG3BPupgiu4WJ/vjIbP6l+iOuO/XhHyvvDJ3hUB6sjPTyYoYyr
2jBEuQUQFsXEOqkje21IfIv/HqQSOx/koUQqtzjslv562Tik5xwwVlZ0XX+IVHSpWOYmeS5XP80s
gbtmafek5tWaPs4N5KpyMBuqlwQPJdcVzTBr3OpIQemYRXZ3P/0Dj9bi39jrQLk7vSlZcZrpMWPx
Cm9UmdDYcAgx07PpetjXbQIOpfUenPoeLN7gDkQskFppscDFHZ7k5JCT5E7STD42lu/fgmueNQ1N
iDY6p6LjgHDPhgJ8jlkKk8FoUXMgOOOKa0/5ZRYswz3SmRCRvlfY47oiqfSIRrwDxYkkRn7V/SvA
bf+PK+nKeuCu99vkCqMbQaZCdD8Go3CZarAfM/lPEtG5Gq/czkBJ48tW5t+e1DbFBB5BcWr2rygO
cvZe+sABgmqYOFDX11iGfivXXGFYbRKf8zGbnz7cDnD2YKCWwaRBFd2Y4m+6RlB2mZgTlFv75tOA
mHjFHQrlNLiNqlrmKlMZhvS89QZq6kcHFfk1jc3nbe9kF+kr2QHA0SDOgiwvH+hHtEVrSvtzY+Vu
+z8KXvs1vARkIMW6evfDVOEMNVjkp7ydtcXGRVf5vOrSS89vBbAzLJ9NQJj2CCD7+A4efvw85myv
VR5z3p8XEQt0jiHRzs9pvk+259vtFm/yEHXiWE9DhkpQwKLKoTdEKECsVtY0LJZyq4T+tyOMlWtn
VN7UnHYe4loBzaUl2CRkk6nuoz/YhgH9EzzM9t6cOVuDa1SYr88MQOQ9xtG8mR/EgIeg3S6/Y+OS
+jyplynaBLQ3bb7OyP+wLiiPgA/8D2G7sBbVGQ0XX3rN6Bek+eYa7VNTT53NqXEGIey4g3Lei3oR
ZrNiLrm6qq5Myvlyz5YnKm93VdL0NLRd0/+SvZwIa1DIG3sARytydTdU7H6u2jv8oA27/Qsl9Gaq
GEZdd/QoqLVDWyRHgEbia8XHpyhad4h7nF7DBbLhtfo9QRQwH+Kp1iPlhmdnprCAw5ki+2+YxbUd
9gRDuFa6QuOvAemeRRzemCpLfmPCCCCQewxmFrjO4r4QYBHPvrU1Oz+hXqlSoVoojmVIg4CINeWq
6kDeUt5nx36acCA4yx9RYr8Sgz+F+43ZQWyBI87S35q0CE++sEiWX3oDU3ufYtINb+ZHiFh2Ag4S
CbxqEgRrrLklZgMEf+7HZziJ88FnUsPGPNQVjuqxzsvHWD6TJ/FV8UdGdBmTDd97ohYFl10lluYb
ABlWnWYXNm019di6Cu+x8SG04mBSCk5gyLbSjMrAFMOG5qYsZwpr/1V77LRMXqXK8HvogjjAAqLS
+0weJPAPlSjL7lubtqXILTXL3HnDvoi5tA0pqlwuSZMwygsYxlYC4BLt/1Wmqw/cdyww1ujwIY1F
9RWGLQe7apa7676tii2glKWBC4Nbvw9Oj41AJvgJQeDnNvSBBnr0WZTDolupe5x291qSwxWkmbL1
JHUHGxF4NmFgDHxyWUmqB2P7vvDk+SDcTOQVy512FpRj+esKbA91yohmq937WdeUZJV3nf0pLpB3
6xa3jWJwZetMVTKOhUQy5vuEG/e4uiuTVGVou08DZ+Uc0J3tH11kY6InGLLMX7tuQWSX5a5Up2pw
QB6VoDEx+BwGzZdJ0auaQ2ulRW41pDkLA+OERXz3ddnjJRSQ/9lJYWLEuf/ZpFA2ds9l3Rps0x5S
xYcUVnXRFsvvyH1wSX8sv9+G0DkxbV4J/pahCm/Nr3MoIdHgkQf1H1H7fVX9xi3NMzowwvPej/Ri
dA/6Cwhig71zzfag0HQ4a7Dp8gy/yGT7Ggr61w/Pox3bwg8jRa78V2AavekK5+wbxbH0jrwb18Qy
eapDrQ18KGpnKBv/mvGPc7puCyayDlM/rAd1O2mkhwphxCtgNDqo08HlPbmNOZywZhVUT/MW59Gg
O9xetPqAv7EnhnoAnWHb5CCH4zpRVjKFLy3hf7GEnxaBV4UlJDsD8a0H2PrmcImCzDKxl5i3oHu+
07OwFDbeie1EWrG5rxtqSgYf7iRtsrtKCMFtlk392vDhiH51NE0++1RAF0r8+FR7amK/nGz/671V
Z+PSKylYsYBuUcsyYTYR1RYW/X/tf1FydxYQ7fZNduwydlfdJa2i93blxglXbH1EImDJAU2aktp+
ZPuWY2TwXRuTalbgeHUR7Wefe5Zm88rfMusyXIIZ/Q68Y8eVwEpsCJW4Q/6flOVvbjjnHdxLenKM
izAMwVq4IWoCXIJn/Jyqmt61kVHGSCTWpMNohYL3TIR+021RWWLI5KT+Du9EtP+bGgwuJIoxvm7Y
at1lSeSHDlFilHV6jfTd0NeYvyzM3defuwgCgL992REvrtCjp2cxvA5DEaP9bdS46g2FUzzMJb9K
jypjjk2MogDO/SDjxSQz26fbdfRwdYwWm4WKx9OJc8TLQpv6sbz/+Fw7QPaPjjcn+O4AbgAelCKF
Njse8XC9jdebBDXKULpOtwyObw+2mqo7Wy7V93TSvu+T/c/hUlGQhCP/PupRyAG7AoN0G3M61w8N
uIGIbFVEZHSiF9voZ6c0bFajJ7y0Q0ch/izHUzHAwQvU9gxeIvRIX8YU/4vH0BS2pJaVEjNa0dPO
60Ke+a77kjwbp1DI1LdFZwcqCtOQlwFT4R1S+jwxw6HxfZS66fFoNIxxiQYhhYcWhqdIsymEYS1k
EZ7KZBTnf//2EZWY4z+/BKixd5DoxYaZzE/ZatGGYhZEDO49eZxLgnRsGnmdSJbujSws/3gJG4+j
6hfIzEOfbTeMeAHV8U7A55EEvZcE5mk6jZ17irSEgejM0oSdSEwMfeVNRAEEYwZvYeGW2v9EJ+NG
uGNxYrsRendFYn13Ir/c0hbqziuvG9oz9EvXgh43Sk/etNgA2oVfq0Ap3rSE/LSm5qfmMHkK7Q2T
tso3ODu4V7Tj2pKsN5+OjRbl/GQaiEYqg8UBjQVN6+Pxw9C+UOU5193VCeI+RjKpAs/Q8PZJBj1t
jvPUXkCap7bnhoygOeXfLaRIkpbaqMVC0w3kCiM2E/qBNoDOQj55rzVaBIqTSrNdplcJNT5Qjql1
sf5dpQ4mHgoS5Kf3EZviDO7cLklyzbfQxzfqXrejRfs6Ni4obPbFcshVfBCAUJ5mAhESb4w/FpYL
iW/4efs4QyqoQ14HVPQsCvBJJAWflMZ/PvWmku4VH5XKKhe+knJPtiThyYq8ZOW4phxIGkunrIqE
kRakb9nbDjv2rC6zA3ociQ5440ihLaiZyJ6OnVWvnWOmgMeNLbfbMIwgNTdv8ElihXHVO2ZPS5z4
UPXtzPRuJVI3fqLIXuz4t637/f6xK16AljwGOB5oYKrQAR0gw9+8FxmmcL2QVcIPJ9K1tRXLjin0
e/Qy2OKkxptgizUg2zMwuan/Z6vy7rPJIb7Du3uS1cWVgEsmsiwMbhot+X3HwYWLMwtpC6xWtBuy
4LBKYsFjjW/JF6MT+TeoQQQSA/gwLyyjgOegMw4/PZi8PuJ3vRGE3B13kaWXtnErGB2DZBZIUrrH
iqjuKbDm2iZPTjTPvBHFfmtHcyjjYrCCRAM0J2RGC5qf0I+YzZLlNUFoafB7s8WBl3dUH+7mgSXX
lFUtrP8L2KgqVKcyN1c1rs4EPWfvIyENPsrCI76ieoOVK94QGtKdz4XEEFEGg5kQHjASrquTZmIK
YTbc4L8qGPjlW1b0cGQUD6B/ywePnwvmv4a89pb83diaCXJKh9r+BG0MT4uaNip23+Bi3X0iMGcI
TyJMfoXDpRqXSUzAhz3zSK8SwWBFfvfLZA71qT+Y0g1qTm+5agpC3sNFgA3ryPHh/tUOV2RebuBn
q2B0l1Noz48QQCT8vhzSjhcX2DRAz3six+po7ccrwJiI1kCfRpqR84HCcI7fj5V3ymHAhMvLBdbA
089K//26jC6j2Ik+oMQ7FLp+pxfZHu5qec+81xlYYLDqTtzyVA2EWtTcAJxQXzX9fW6fJe2qpjXA
UtoIGXt16gmvm/9StnKyOp6f6aYnNEZY2HsDMlnpQOzr2sfx8MstKDO4itI4nCBYFhH0AnYHp4E0
vh7UVoJLg193oMhSQEEj2XZcPbA3OLk7+PDtDHIf0hEUv6miiEAg4FlkuIPQ5DkBL8d196EcL25U
HmHt1eT+8XHootTsYwxMGAx9HATHNpd21ztbkmOlWjyjR5bgsh9QxM8pIOd08bF6HFqKPT3/Ns/4
+O+lhnhjpHID0IH+ZWwdJEaL99Rkpfp4vesI4Q9sGaCxd/1pod6BG++Yqf+5Yy79MlHuSm47nXzt
VRSf875sl0FdGSBr0LTR2QNA3p7leD6fkvlFK5PO4gQZ38/uDLmyttj4Gkw+bYBm3fWSEyGRIuro
TK9M4Ax5BrB7qTFsMTnYgKAbDbEYyEW4AtK6B17wS2gdYXcWVdPm/cf+KfNr2fJURFFQZMDbmhuI
dlr2S+Jh5CFd4S/Cuk+4PPKwzVmn5xkmKsCVgIqwee+UC52zu4EjUN4XAhYMRJnGjpi9FBejKwZR
pMDQSdIzQATjQKTGcl6NNESaxrazA0eJRG0y6f6wuZAIdWrzuw+EQadgKkhBQvS/h+mezoXBolKM
QWDT+DdCosLpi7EJ4rHO3lT01VqyFmCHoKKwjvfr4fEAdd6ststs3RP+2OxPB4Ime/zncEk8SfNV
1Snl5h6DR+3T/vfkAm6HXfslFkIBzVTEiWtvd/GLMq0dIMK59qiwZrHmRFfntKL0bEOa+3RDaqXp
gv5rlfnOXPxsq0dp1gnfAaX4VB8OQ6zMBo+emSvyEfHTcGS28w51Hxc9qAghkzDufRaXhPsbl9ga
/6UW8PhF2Txb00p/zDyDtlwMpPkYypuIqPnbOjyrwBR31BxGVAQllIeNPnxtP0KuKi2fO9wvjGbR
bv3kNxv5wxmhmMVXL5vjgsYlwllj4i5+9sz5w9ySeFT4IbNY77yyy6VpVoWUTzWrAz/6YqtrfalT
VrVD5T7g2WZ2wpgtMIA57WvVdnIN5naU5HKrjoOG6aws1yxgKeXU7QJf+yvFjPbf0yenZbmDhpAy
GYHW0nd7g1TfyxF+nCS2DLhxQdeB6KNJmAeLjxooBGL5XVoX42v1dpgtwAi1jY+tbl0DT73N7Guv
LgPziHhXuit1ajuTsN7XQY9xM8KycEY49kRkIugNZghgsSJIqsadlILt7eS05rXlZglcH/kGx9Eq
pej8HnBUOTG97EvYVpPCbqgBmilWayUya5fBZO5oj7Gb5UXwhruD7dSqgNNciO9laabHceB/2Nvg
XJprd9HvduCPU+2+0H8CfUpUN6plizROjuhwienLp1SZ2Ac9YG5Ose8b0UVNcdWtpdjI1GtEnOBJ
1s8a9IH5mHysdzX8WDhnKJlYvYEQJptC7aivqU4RIroh146F0cLFk5op0arU4fITBUFPZ6t44kDo
JZE7ToUJmphYCA7Pmjk+SPUXWvAlWwLN94018ehOkxq1wKXU1qDz+cQnWEwfoBZ/NiaXzbovyZEI
vEA8QHYMAZqu4XZs83ETKJDvynZHDSo3Tx16gZAmQWn7Q5cwObFxvq4wmWww49jEF3pbqnmyouUt
WbIZi0eJZOl80O05Zcs5bJE1BDVuJkLOCQ81lhLP6+B5el8wfNnIvjX+ByRXe+ERBGhzLa1a6ksb
7KVN8aVAqXKpT4+53cgnp8/TPQDwr7Iv999Md7bEOq2Ah+D5Ff05pgxi4MsHBAi4BVN11BF1uL0K
iOkHEWeKvNzS4LvyPpPz6Ie33Kcc5T8T8aXalezEA/MIAXkRWqKJCEwiWojzSEC7Yl8i1JDERDzz
8ARP9MAu7xEHEZsfTVw0fMbCrB9+o50FsPkHoS+CdSdd3XECudgSsVGWGGAdYQhNEqpnHqZjhpim
9WdH2Yw/Kky3SAkRESW8zqKKA8KypCbwjzUIJ/6Mh7knWHZHxZfQDFYAI+Fs/n/uI2q98PkSvQzl
WuSWWRqPl8v1cN+loiTfNeBG92L7kq5De7jmyYQJCvQu131zU0wLDe35xM2mxdPKn17LjU7Zih5J
Yg6t1hiXFTMInJnXTzv/Yg8vqrocAnjQvXYZW3Pu+5OWlhwaTq+exgRlai1NmzaeGscR83j4OAB0
uVyuoF0uHtR1LqHa56KBSen+2MZR76OziL371P9/cKCG5LYfmDE8YR2QnDgSXltunFrVlEnzWZCG
BYbFLVX25mNPLP9JtK+hu4ub6dpn4H+Fc7Ccw+ef94Cb9/e4pet1seR2bQzhpF6pjTbaN5fxOyuQ
Xbh40wo408KFgI7XKBFWFUoV5LVROh4HgosPO3rbRATXkMxZtO4hkK7H+Yhcrg9svZjJ1Nos3O4r
q6Zjn08Jeef1rW+HI51VIs5He/Fy577Q6ycTZOO5EzMshqxgrZilxZOwORdNe9LN9CEvQ/SOsP93
JBG0Oj0smG11/hxAZdRUArHUr9shaCpI6OlIMeaVA0UgFr0bhX6ramr2tT0zc+Vs3qgp8MPDJsCW
B8Na02D8IHFlP5oAHN31lIkxxAsjRtnA+gsze46gvrJT2gFnZMtUQ63I90VmZDNHjTDYRjexUZQT
wiVh6FDRN/jG2TkEtOumJzrI2hGmHBPY127aQlS5EtSu0OXlZmdVrdbhA1c9wH1gPAn1BRsToKTK
1Mk4VTqfiYGQmjgBxZ9gCch6kagaXGZbNw2LUBLwGiKPc3ySW4GN2dWRzD3pI+P1xdVCO2ftdSMp
eYM4TIofkgp3ww8FpJMzeqzxr25LUs5OAK8gD4TxawC3lPCCl5xqN4hhNrVnmKtKln5HqBhrvtxz
7Hp4eKzhckP8Hf0czN8FE9sPhHKkOrT7buOBznJztO1oabsv1maxflmTjhkMb9LK3zSXpy4Q98KP
y5OEIuctW9VNbG88yU74GmfLIDL5JFwBFMRJCQHBbztWlAeCFlNg56r10Zo3jwCdXMxvkKWgDqDK
jTW8yKx4EzsbTLe3qpZ2eYgoevxKp/SS0fDar3vjJ/yJohvHZ5jBja7RLmVvD+F4AYnSPaUdA1dV
ajrTwwEV0wWgVIWW93umVcuAXyUzX+q6suRJG9YWBTn6BJ5VKype1LowMvJ22XsjBf1zZmpk0LeL
4d31yQY8kJUenh2Mv/EVUHLRfH+vuTtlFv71qvb2mThbluDrVW3sPAQVKYoM7jH1p8I78NXo2vya
NopGjGAdg/UzM+4mDqdrI9rrFfN1U+mrq0GWbvnlu6GPuumzjV12ywk4Ksm68g60UlwA9CbWzGq4
0T4KxtTsbpfNI1QfWO8=
`protect end_protected
