`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n+htNXLSuU/3gao+frgxmXUQTli29QIRNGyQ0887RUnAC3AgiCZ1gTIU8irsVFEuTDgov7CTyrTj2Th3NXOyHg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UbcfJmAknb0eMNrzWO9mJ/9n9LXBVNcGsvOe7dGu/MMuQ3wKFfbcqBiv67hG056/LbOiX9My9K1m6b5jrwJxHZv7pDEneNyz3ROEqGXsxM1LHtn5gxpp2xGFNHHV5Ne/gtos38uCA3KRqoHGNWFYPRiDaX06ie1jO10Pm5sz8QU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JWJ25mlKufPgj2BD4GZrJr+krJHhQtbZnSImx+Ec+bXn9m1xsBWMNPNCuOwAjRRKeYdcq1TxYNJPghCHFqavug7WWKXiFG+V0oZLVjK2WSbLfgKCX1KPe7NXzv8XzYanBNpUMQS94bs5TtjA4Wty7FPygFkV6+hsv8+FrNR/9uoqCOt71+osj6Rrx5YCr6V7iH/oYTpT/7mPaj3S/qEwHiLpAwmn1ldJyErDP0vl/duRAAlBDdTKlse0jidlelrneBD72uNocpqsCw2m5hhOY4bz1o05SXEj4SkZe2/9+V+raBDw0+uGO2GfROa+F8pVC6nyv7nRy6CJWVKE5dxFjg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XM4lPtCEPUqzCZeRfc6+LnEZSsDbFSdUOyNB5fRscGqoGTu4liwHIAjww9FDOwWx5Y+UaJJ1OjNkA54uhSiU4nja01ClJke6fn4Dkd60o2nwgMyAJBuW1ZxMEiPSLVWxg/tn2+201Tc98F0786FLtYXv1chWdrSMb2OCXuk0LZc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t77k8TCMmHVA34DrEnwSwCxHWP5bV+6cfbB3HhMOheSDBvYlLfgxdG6ggtGXuEd1pQQXT3vJHzQBsT9071csCfKqX0zC2Eh89yFueQVbWl1x4KWJwZstJV7OyXUPsl5LyCVbTd4Z2t/sIpIkaIX/Sw1cV2oJNlQqsU5cfdz/LtgRm6suXzVrN0UfK5HApKrT4TBtMOf9CGuB8W0l9QpCkiwIe024AIMGZxjG6gvr54aaRTnPKdcmOrU0V0hBh2CsQSjgZVta0chk/g0z4VtfXzpJ5/R0REjTMjtVedbmIDjVEj63cOQvC50VFgxHxpbUJiNM+B1gty2jwksCbbCZrA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 596442)
`protect data_block
43a+oqdy0senFSCugCyqMBRmkdA4/90SyNlos+N80cBfRa+tE4YrhX+ZjaqSX1+1c+P4FmjGZQTL
BNg3nGCiEp8VbaEkBA++/hg+rJDGnvsDvFtPWqQUxjy6ZZZkC336LMR7xsDZbn5pEd5cufKl0QX3
4nImRNysOn6CncRBegEsFchKwTyrKJFeqBhmduqOXtPi1H9qWYBu+DQJkIn8sU5aKfVCCj6CECzl
VfLmscd3wSKEFIgTFldzzzXWxEZvvVdGEM1bq6eyUWou/irdwia5WKYwniTp+06eGkmSqeUwvukc
3p5/rg+jip4CwIE296gwIkuJslhojwaS1xB5Zfn55xhjC4pKfpI8X0UazQmEbPri3kDB9vDlM4+M
ekNTFRVT86id8SA2gprJTokJneS6XTqY0Y9Bv5qFjqhBCKgEo0IPwqmDF8djJjJFbs82Xv+Ud0sW
F9YjA2mF9VvTB+m5bQ4fFjc0DL1h7BPs9EKoplw+riPkeYpceanRxHMx+FI5f8P2dOnKi3AdjT6g
o5WT9cnIN6/lCGB9vHKj66XbzJ6NSmgLLOwizQ+R+jNYRSdUQg4Y0leNmrr2r4ANYdaSGFjbgOi1
HCs9TuttkOEkPs81Ur1FpmjV+zmvPGJS22PeuIeQEXWeUQMFARdkuqIxa7+dPx6RZQ2Sr8um9srl
Om5n9PchsIS+1DbjfJXw7mJ60AIaEWLpDDA92xknRKUDwhHO4IRSg+msbX39KZp+BZXj7R8P8ZGx
MxgzVYvSXh6p1ZoHM53+g27IJCUQ+Of58RDVm4aIwzNkM18sALFXkSu8eCZbRXt9kCM1drhDPt6c
e6varaf/a3SfVoacDfTD2mM9UdLoAkf7+udf5loAwB1ukxkq1rArYobTdKFTDg7pScNHvG1Kzw/k
Fz8EMe5lpEbkZYEImXhgBlV5vo6TcF70THpdGpz229CMkBc4yqZABjyZTUVTA0y6//i7v28p0m6G
EQuw6NgP0ujlA7fdUuQ1gFaQYaTVgjN2k30ij0S6OazWDcczbPxeYyfg2lEoJ8MVFMTphPoKGML0
76nm6ff+vs/Ll8ep/9INAWskSctHWL+P6BMl/fWn/zWZAwnWFMcy9gUU51FeOoozj80WzB70bWBd
IC+5TeURt+jNEPPqFd45gA4ogPj3gaqMikasthlESS4SeBZ/WmNp5cgsYLNlxMqHxtWNh8K6P10i
GGj5gdRLYGhuqRHZJTLnj+L1qMdHgLpoCLTPYIwIpWVQP0dkFA7Yk9PMPjXoFpMPA/I3P8/C61yc
WBmgoXN1jG3e8RwWHryg4HW4/c7IT8sM/VPZ9jrVU+/58c8U0a8stkvPPP2Gz0VoeVsTiwJbdFuG
+RVcdT+3G45Gy6E+RJh9AlK0+P8WSZWrxoMafuUcJp5C/o9H1eCFbsPjTiG484oRKfsho2s12ZIs
d2t7sa/bSRvpU0AqxSEkHloDOXMeTKNC4lsfoNRRLMTyVLzoS4UepvuM1PaxX0Xa7cuF5qvR34Gc
Bm7Lf50t/YUWCoq7quGrx2mxjCg9Frzto1tKpCGa5dc6olnq09FczHlulQzay+R2XiN9bde06JMc
VBnrcdOKLXTkxBTDWg74C1W6QzQ5MN8fk6qWsyIP60I1vIBRNMXuWdWuVz9CoFKj/6bFWVtJtsmK
Lq020+fuNk0LHGnny49hZTylFso4bsoz+uLeybVTcjTk2ajLBB+31qeknZwxETigDEhMOwmtVxT9
BQ9OtrVXgtaSZ1c/EbM6FoULAHxjxCegSHd2BHpGs3p/arRBgFBlM+gH0EckzfIxxp2pXSAUUm91
p29k/3G1XZYDxgMZXkyWHMkPvKh1OoNb+W4ep97BzMrn6wGUIzQnbkGYevJOECbWPkb4nE4rhsd4
HSAKut3g0h2EGHCXVEHVMa3g+J6gXyFvoT2HEyQASjXym3FyGJrWiicUh7GJQ72fxQLRtBhlS4b5
TA0YNPk5KQYwhoPbqUuCU9v7A+9tkJmRXdB8uDjNYfYFdYsjujKYO2id7M+vO12InFk0izUMScQh
qB6ta8ZQo2oXxMOEDu4xlw9RfG+25jpp3XYmeapAlW/SRPb3+vQ3gGnqyYF3iGcPyPgrpPdLcwqD
h2CDXQNnpqH0eLs5/cmQeDQyVP4Dfg+PW1hWwBMOKRMgFQPdmZP8G+vIX1v+1qk1apLIyPToZBoJ
POn4WwFOEoLO4JTdYwIaB5rjqCG808vBVmM2OvibA1UAuafUr1c6+Z9uH1txznGtYUQbyJ71DSop
M5TK7ukhr6P7wqxDKu+x4l1kvxb6VVf2zfkV9dK0+eyW3oPpzFhko07noJw584+JtDZdZkURbxeT
5ouE3etlUmt0OPnisGKFFS8bii3QGfpBbyiG38Uqf+NGouvrJPP/uFPA8M/AkEUvGVfWPB8m8WR/
SoLaAd/CIMWp0clg6N6BIHLWHjYpa7sUQKFm4Ui7ZOAueXipqKDgU5gHo4g4b3vGieU4d9cqUKO0
e//fCioJ+upaQUp6HdmrpS1CxHmgbOpeNVaV+GybPI1qJHuOXMk9WGWo/INW4CfMa7hX52WYKToc
72FELKoa2zxq47ABZ15qYyX7yp0HjZXyBrNvM2Uza2ULcNdtaqtE5LdjxxEqW+t8yR9gItooVxpJ
phOlGu4k1ySkP/sjSNg6FpcC6EyavoRfqQAjSMu7sT136DXWpQQqzqeJ5DrhUK0k+5GP3sIKAcoy
eTmezRxVLLuVU6pgwfnOjTphwIlz0fv4DV8AGXtP7n03KvUtpn+qYstZaCrqMVf1AfKLqk5NXjTv
NHNg8Ub3ga64VqFH/+AP6A0P/cq7VRMDPS12gtcZNZRTDmETNhKZGLncvkbm97fxL/fKD9ZSZi7U
6M6slZDwLtrJ/0/n+P+uCp87FDo8Ae2apvS4hnrSZgUsjBzD+eYW5yGw/hXpnJdbejOz/8v5USat
fTOojodS1dgZDYUu+d0wzUe8zXiA1JHKm8RD+R/tqRL+38LsrsuklGf5QqM07tMzlnkQEaL41fWY
nNXtNupIDIaE6e63TBQafarO36wLFzrvu3bw7Ry06qAku9Ci1i1f/Tf2hv6AlD1HVrBJMr/g8Jcx
m4oLvRTTaojGClOa7Bq54hwEHOvXsocHmKF3Td8f06Jhz2WWRW25ic/kiTUL1gSBv9QhG5eNUEJr
weN7+Fd5w0B6g+VjDcZKhqtYLQb4m1thFxaGDjkF2ThRfYLZV/iH2Io2Q+SXlwfwtIRuxfyDCo/D
4d4PvljxxcnukCJ2KIlX8tl8PkO8G8GNHVdU+Y77VU87xpR5QWDlQpl3JclOmeywIge2bcw05ZwJ
6espHXdZbHMRDi7PC989nnRIM4OFScIz4yuEcBoDgU7x9KWO2aKBdV6jE7txI8vDgvOjJuNo7JQU
VRQPNxh+WSb35Al8ctIVHcqb5HKAgY5I9UX3pB4uRbxFJsRKB69coLZ+1IuGkS7v2BP+mcZ9bxCh
qKe/XlmOCaGqp4h1Sq0bJ/9bDJXwpu8dwZWftm3V2hIHvmT1+LtAZfzFQKQ1avsatY1dOqGn3Akb
XgrzvTt0uMelnFziSodAg6n9oQSUGQ2WYeLk3DSNNrqQPJyGhNo75MdyI/05dDzznzayXQPu9u9K
w7mj1uqswZ0xsHnPewvmXtT0sPeghHa62KIGiJkdKtM4Urt2B17XFrlw0Lce6QzKnpLO0q4atCLs
o+FMac+GpYjVe12xf3NxV8IGGBE7B7KHyX/qK2VfD/4FHZKp3IQYQCN8Bxu/SCRNXsNBwwOmpouL
2diWrhXnBKyB4qxegj4aExcG/MPnQkXvJVeodpaeDJU0e+sNnQbKj22G1so5QEylNePPWw9S3Pz/
87rgp6ZGs5Nyuunscxrn6eL44zMtZNEki61riOUWh/GFmrOkibcizQPvMVi8hB43BmWG/K+e0aPE
bpvO/8UkQvzJ6zJBZ8o9l8oUvGhs3ST9eEF+3YHb/RaEqfGtlBk1bxQE02FF5F7TRwMZguusA8Ew
eDCiPcX1jpFdoGFu3bn7ULOHidVs81SMPftqVSbdjjJKCsQn4FgmKj73eFxOd3ZAmA2BPZJ5IK/v
eEwS5KLgr5tXBxNYD9A5oEq0blhKpwL2FTsg+UzLglwLR1MVhlI/M4kImL8EbNvtCwu03oZkxgSC
+W9B6TbOvqkABMrinvDQ0KtG/9Q9mDOY1riGUQxH14Q+7RiF/gi29DNhwhmzxJxO+joVn11lBgTl
mjaMKSMskznVup3vk8WM0QtJWNKAClFYP17qTOGD0eEEQlnnlZLzxGbKFys4kV4XYz6rzQziOtU+
68NwFhtgv0WQOXL4XnZFS3tSTqBsTNv8W+EB96qVdoXwyYBoDsSd2VdWcIC9u68cBVGUS6SRFQRF
5kG+tGKqrqgpcy0yL2e65rclWVuCWPVnauF/+vSK/xFlC95qzjOLhOqxWGtgohrYITBFSEVso9hg
GAImf5bP8O3HXKlTxYb7zofiz1ANImuAYur6LhaGQ9uEAbw9fjfX36uJix7VVIc31M4ZmqcIDeZa
/C7XucR6ES5QLc6oYWFbOTQUY/RUyvb5JaYwN6jscHqpRsilfoFbF2fl5rt/897F/hnn4cF626Kk
PzAtheA1jy4sdBtEpqHI/BZN5oLePezCATxP9RvPPfnkyUd1wCE2Jp0ULs5T6oVWvacoJ+MXLuWA
tbDEnDlfFCmnOQzH1161zL3QFie696ydWHWg9nOMp+U54l6H5jZM0PqcoNUJWzP1c85OcoYsjDZ4
NT+8FGejzBZrPDOanSEZP9c/jVpJIPwL9Ejl6uBmkvr8bMVcXpxMNl1dTh9Mc7zEhQ3yCrST/PH1
C+49v4fmGDYphsR4Wzfx7mHLhCmCaR+NNJkxm1QSJU6MjEnIC5TlVH8PZgIV+FMvtCoQ8ySkhwXD
S8bfbBCMvqw8KulPbCnfzpANQJl3eMyoSDf31u2z9n61HbiiH/hrD/GH0MaP2uwOOfSBdC5QtIHk
zICAJWJpqn7l0N60VBJ4A47qaz8dggo6WrDNZ33fs+GuBI6wgu/RgRRBri8BlhDVZUkWPIkmdFZf
GxFVjXDRDer2V9I1gVG0z5fK+mCEZV+QJeG/cAzwWOEPr8C4jMicdhqHPZXx8V2QAG5vdaD48GmU
52lqun1USlX5rAAgQuwCVdo9KwiG2F/oQMXtX3kCq0hgaAurWbSTQUtFxDuP8RY/Z0skDlf93Sy8
gMu/Oo0dYsr+Efk7woa0vwRUvUkuAAFJkfsjL6GMXuRdSRg7ZZZLwzLQ6hVEDMQubzr+0JkOxvG/
k6NC8xcR9Ths9RVg3dG61sKgDgr6Cj/rXByaCz2+WHM4I79nJqvhucFbP2ZcoZqbOKUXKrsKRrNz
iWP7Sg5zzCh1OoUPSYU3ob5hYrSgGzvkGgZi6Hx7ZTzENtC06n99nQkK4OINTd6AJbDXimsc5Dkt
sRUKypQrHeuXNnFuTDncUIs7sUv/1RCG2UFpGt1dDdesZ/z3DIW+XWD+ChBy7m0NJCCfWlPl4Nju
ChUwNr6JEiqt5vb7OFhGDbmNOwKrilY0R+JdfFiuwqZzEcTkZuAOcB+szylJKUXAT1OHVJ5SdjT4
eADZLupfCdjUoF/nx4jDQV0I68ssY7ZoiVES1ymn735ss4/P8shZLtXFXFE5byCImpo/Mt/tjbj+
2+CPB8E24En6AINEU3C5RJae2Wqj9R63rTblBV8d3F0M69I9OwZxzwMaMZPqAILU+9yJPh55xCWe
ibujrH8wo1AtdaWJ9G9nRBlAvDtze6CQfmyQBArOePEL+DUl4B5khLXSDOb7kNObXBMIBMXKEUzw
8mpt/blQISBz7/O4bTgmmVVXvEApWePafLj0FlIx2cSWtv16DBbBY0gyY9h4wyrKZtioszIzaQAI
NHO51JaxqPUbF/I9ghPBUNDMP1l6iai0tBHyEYgSnZ4jS77giKu3xWWvOe3dblRJ0P/4HU2/v3KD
UkhSEkHlVnd0hob9g+wBhr+tf+EYf5E3vM8esqX+T3P3+rYgFHZ3HQ4S732s5c1QPh3XTkmNfHBY
rYFqUBrTFWOT5nCSxO7QplaBb0CPBu7usK0CIRht0mE4MCLnUxiA7hp5jPmHCNo3rlYf0SAE6sUt
pXhLX97ekcZoAkQC02z413vkU2VjG+ORtyJhm6xBggTBToBAR5Ykks0fJMB9KD6h75IrS9EPtKMl
Hz/dgSz7NOoB14q9taIjeQ4djB0ARWmP72L+bRbvlXoAhgL95lr2Ttcvcw/146MQTeIU4cso8nCg
DgMt+KMSXrktW0yCcVvGKlPJuw5ss2HV84qxbwW4y45Wofwx5e89R0euoi+re+mH5WJTAwjEfLhZ
mt5rnh9FqJp82LCHLiDPg3MzuGWtCHt/otY1TTLrdiEIv+m9R49jxBDoUM4flMu9gYAHP3A6vl+i
TVVvBYjAo2yUT5ZxsixUt6TLzPG7LrF/NqXt+KhsugZMwfTumPhxIbhZBJpdZu5/fuSprtvm5vZd
Obo7imxbn4AAdPY3Xb+k6K6MIgB4Aom/Pb4aii8SKCn2jRkohnAYTXgZNmBPCYtzAltwTU0rjGUA
4ZV9UaNbWM99vl3JWvEd478jkwafJlmRDY9qsGGsQS66SN7+nTdDrYHMLDr7es+++zxd+edTT/Iw
4trww7Kf/OlZEaR3pfgNmK6wb2mSaHICC1SrKTVz5r6Ea+oQmEaGttsnMflanyKZYOoYoJavLTfC
U33iXRk7Uk6tMYS4C1Uxoooye8KPssxFjvVFVdQj/pMpTe74ZJAOViG+NzOr2BIx6XT4oiRI/ANL
4bQujV03PrhmN7ojXUS0hi1sxKe5sb6X0fgoErOaeOm0jnjVokqUsgvmr1OJllv8AogvXw0yRZXN
9rbCGI+WdW4PQ2RshozunX1jouclvDZBEzyGic319fsn17XRRqmZRssdeMIHdbnWa7yPUw65mpD6
3a16kkBCkf2VFjs4MVzrcaKZ7nwkeMpw81XNvd+z1vFc33IcvuTcK9pwdNNvsmLUaAEsPRPrGy62
/RAZRdc3dbea106zvL/sWWWAucfhS85Zao/9u9qJiDVMVERYVQWd3sP28dX1LRcTnkCQkRS1ngGH
QZ0OdunXBZMMFFdWyoNQ6RretvnNhcMO18yeRhoPeepW5sP3Wov8Je0SIggAyL11p8imp22rpAzU
APi68F6/Y8B0+lDnLU5aTxz2laCwwipv4IxqyQYGEQnwau1gY13Ba2SQlWC45e5J375lUt0zYIhw
1UeiYcQTN6U1pDbz4sWwlektpyxa7ZlPIS42LYpK+SUv5fOG38H8G7Qaxhb+El3hLyRwkPNK7E9S
lQNI61cWPpumgkGMMT0GxY1uyxS8S2mOMHcdMHJDJrn72QrIsEBTqqfTUc4r/3uQlXoFCgpAuCUE
MoNA/tG4QY/ob0jfe9OKQNv3cLYSOpE0BNy2RvJsUL/apNgo8CF+lYR6oZ7m5ZmsIa2qBvyuEcfR
tY0shkO7dSLxUGUcVBkjgnGqSq4T1vyW2gRIkOJC2TmQnhlADxmzHJtdd8fuwiuRTB4qiFpDRh2K
pJeSR4QCXwRil3FHPxYiai60qhAfe/KVQbu/5vavNJZTO9vGVBFdaad0HBAj1EKfKUTLtwdE9ZVd
zvpGFwEd2asFz2N5TuuUwpW1x9dGrcgl9P5S+MAnyM+ZRNnCxWLPEei1TAwUlGfAv1YIu16komMM
IMXGtCN21GyQyF5weg3m7p7Hiz6RQeLxUfTcFDmPqAcgQOgVMR2TvYkmEDd2oG05GsMcIlvGhnrH
jFYQtr87GpGnz1aclx6Tb86mXwUnITEFXAFFwjGEDF6owmM7ivLgQX8teKA+Rmkj43EhhlFixQ14
GdBzd3RiWUfjDlDh45GwZto2bkGZduHVDrJ5NWqI3RC0Ff5dV9hpTWVNDFG86hg/0rIqKyIOLHvp
QwPe1ZLLZ3n7euQwQ59Ut4M+sLuqcAi1ZX9KxJ7PecIx/f3Qv2Ukkr0m7q+w+/7xhtNRHwFHiIsQ
+A8OvmJiL8qh9JaGMExs3pErj46NOIyKev5fNgZ56N/f21b28JxmHfUtM39fax4y8zIM4tjgSNCU
1MfPAkSL1cEc4znvgCZ4gwP8o10pZ3iUec9OLhW1J+6cZdJGQubLle7btjNibJel2xpYpmSLA0dM
Pqww0wrbn6fCZ5tTctqwWH1IhAuBBbzvPja4s8HSS6sCbciB+RfI7D1FmeEgt7WZBFEWGGi8vcZy
5DkT7Rugi8niZznOaeAGOYiMZSH+FRlAEFuaKBawBnGn9FOW1fdgr/npmhoxEeDCL+t/9xBgCneO
CuJ3UEgZTExVOwaTvAgS2WjuwZ0+iNNi1cPknSRrduwwEqcEi52mUc8WC9oKnuFubqEOzN1fSLMm
cTbqzHDHK2iaTwvhJpJLtCPHnXvmlb9MY97GKID6gz/NZuTgeea0UFWY9PEXtkvw8HfY5bks6OD2
ATAmgW0Pisf6uOFNv6R2K+QmutVbUsSi7wa++2oWvUGigV8hjs4O1YPKb3XfUWvPGvhnUhmsCTVt
zIOoVTpFqUqYgwtoFHkXyQrox2YdqRsBIXuhr+8vdLPfGP2OeAcaV3lsFefwMKL3M849AUBtDQ+R
dxvaW0/JCuYSWXTSTr9AGBegCp6KQxRCbeP8zKcwtaNyPJ1Q+w0Da38DYFGVAvsk28iO6E304Z2F
KHDFfB0qiHDrbw+exVNNpq3hlYiFjcadXW1riWpCo2ylrjFg7V9MptC+7d2MtRGwSiQrlRimjY5W
W7w7gCdJGs2mij0LNv4SEpCEJONgBrMFeclomTyUxBlapmawKBAOc6likpVHzgFz5cQBwMiT+fp7
g3KCxd1kBlg3vMCYsbzJmvkVocs41oGbIU6/tubEhFnMMn5pWE45oJJOrjXOYPTha34mpjFu5/zO
zPU+PHyADsxi2L4BqWa3RTWAawrUMQkET/W49vG4+mThCGBm4w7SK4o5crzrzGAptkO24Q9rtQto
pxg3lD6UwzvDOeLu7rBn7MjGcZ6pHmdYT2v9c2Ce0cxolb2aLo78kU45c9UkpfFUkVP9+ShimvFG
I3zFe0zYk/385PHxm1K1DZfWjac5M993KhYes5/q/jFoHb5h+KyXslbViJfq2ol7K8A8OIl9Q82o
fWKCsc9bQYiDdCdfBE/qcwbkNarCKaqGJiw9sLnWgwJ0Swu+wVEr94uCgNYdk0t++OTEoqhoE8ux
fxNiReooEJbnlfayKxow0W1QZhPsYljp7YiebL7uEd6GKO4kruWLbeF69iEncbR8Dm0rHlFppq8D
IMZBz7vXiuQ3wuZZMkUvUn+BVGxHX9YQlv4OtYUztAGfCjYfKYuBOX9QgXFuAssVy+mOA2yMBGvW
iwqv2QEPeYkA28KrbRlUMM5jtbpOY7t8lBDe+LqTjPoPmHXH3Juyen3aTjm06God2KhipuwUDbuQ
p/BYWbscUXbxHKgB0eAl5183vENqJd1gQ2zBKYzySkWVd8vr9tjDhiJs34SdxvasVS5CH1NGaRWw
7phVwscJMALaOZCsvNtKl4cPg66nzmbrVISqyW8hjeA84eEaqwiBihdIIthRmoO63U7iD8PrkJfg
9IL6izqsOUe+QwP0kYrMUv5MXFrlFzVeLlT8XxXo/x+nsaaXiZyZlfAr/ZKWcdvPDfRQAxzS7q8o
rNHUHpH/cq760n+qqKFiC1k9vBzKZXw3P2pAtclMXuqo7d2Y8eTbaPMbCmQ9wcppWMxakA5MDPxJ
I2m91SpEB/2D1mjsxOb/El9XFvGML2cvgMKJxLwwv3gywM5TZeTfyKX3biH7s3aTKm4K3OTRIavh
9MjbhLT+7INUoDBhcvuU3Rp0jZXlsgp+DvH7RmbueVNecvZOxwhOJE2VQ8ItsK54l5UYsHEJP/3L
BGv60b+eHonXsXxdyGbj9JcS+UCF4+070MYI2z9y6iNumDJLnwse9hF/TU5eTNTYasS6CWYLWMA7
82oePj9UFK+APkDdK4jCYLMDU91dbgvf1hgqnZJ8XH5CKPYwiu0Hi5hpUabyPZQRCfbSq/bgglc2
T3w5Zkf9rhAlcTbnmnnL3k3q3jbZojiEumiGAghak270t+XK1vqiG8tOG8pAuUCATg28hJEESbM7
RMlKG04AOntWMFAwOEWfykoLCLjmQNjbMM2PmjkCUs7nMqscj56DQ5mBDyFVPfqMhfuSyysTXFa7
R7y1LQPQSV9KLl0JTynXak3AGTYJgdtMNqB7PzikfmhB7arGZcswcK4uCnoZA3DnFYWtiju7ounk
aEj5D85tSyPfNVeStS++6vAc1A96NFlfwljjErkJ8HffjttFW5GuuSp4z5lCJz28i4zQC0sQtlYR
R6xrk8n6LpNVbEIfFLGYYX/XGQPizCiVdl4fJOpZv6cENQ8jXLWUlDO6MZiojs/8qU3khj3gIIQ9
x8CApy8liFnhlJIAdFgq0/HKhZ/XPCEKSfjkdkL6eQa7rw2SUHu2hNV3X5QZvlewabvgw8yJR8dA
ZNmtrLukzKPLjMeF+lotUQ+VDZtjzUe+JYimrI+04ksoyBNIHjD9la46GeDgZxjao5kOXTGVZqXU
+E9uGPIHwuGsC6rAZXUv4Iwz6RB6Nf8MNEL2JYWwb4deNZvx7QEzkjb/u0Bfo0Anbas6VzjqBjbk
x2JgbDrHOg/nOERm81RDYtCpT7RTRC3eg8PF1669GV7F/NTON0xIdCICvzaAnWfgbV0pXKSFeIQf
VSA1LXL6cMpX3y3QVm62FYuU+UYcBkftu1DurIN76tNH/eoRmpLctctnVL7R9Y4uV1XyvfF5hk2e
ubPsA9u8FzpCKF1q9K29W8apHnjXWK/UsTO/JPVdClj9kSfScE1NY+DEDxUBbhQVazRJCITqhTOR
bl2gK9oMNqSautk7NkkidtXRQEQTgyomhbmCavY0BfOe1oFUTvMYbzqZT3Q5yAxFvn6Ph8ysaFiG
dzx7xTI3iP4C6UnNHjZUxw3cNTH+mzuYL9sxqbIRBmmJBfRnQktPtyem4WdbSENooLvnZjJgFuq/
/E6VURS+fbkgloZBav04QX9aTH1+N2Pt0KxuFUxWAAgJ/HFXhJMm0ZKaxTuoXRji6FIBJEOZgG+w
btb5UvhHznncu2SlChkCvJICmyYV2Q8Qh6VCG4Uf2Vkon6fVs0aTfPUobWMz2Hj9/SyDJoYMM8IV
wx/it1TEhB04NpAsmio1U+Nv3dUklodMMK3qTjvxNBRvFjn6JbC+dbmpxyptf8waA/4rtIS8axRJ
SrC2KOmAfnEeuoF0GDD7Bp0rd9kU/KtTAxXf2uiez3kRBLvKnuRRt83KR6Dij72BFV8WZmsTXYuS
fpwiEYK3LIgC+QV4LDJkTVV4BlLGvAswLnJFA7NpfJzY1TZBWs/KrYtZF4ppWEs+qt7VP9VfC2m9
SyBhlARi1gJEiU8U2G/Cb7tc7fOyYzf6OuXcWz6Rg2/Li2G/gRVOJOqSjdFqPL+Sk0s18pu/t9b+
sZFupk4nz9UlGA/JRy+HgOqbA0RfuSwM4MJtAEEfrQ4JaQxJE9f4aI9JjHEqYcN33VemNCVfj1i8
JnpKUpznp/Xzjj3FVc2d8iBwmfjXmjyP+w0iEBAnt5advLp5fpkQ2D3fYmdK5J5klhOLXWyUfY87
nfrwEgieRibNyxanSiCGS7es+P7PapSsowdkMmD0JFlZPSywa0nEQPMAqQLMY0IYU5Ih+/BlVFrD
iq0vfAKmLRiPFzZHN3+MrES3W0iqKQsQeNaAcpWbQAObQWcrZIU+3RJBxwgmgqST1piXqgSCrt+1
GosdCJiI/9xgMOX171eeCuMRf+bDAGic85Q5F8H7vdEelX0lA8k6DTAc7CbZ2klySqy+U2sQlPb1
Ghbsmd8swwFMdhZGdBAB6VCtBcIEmtMvviECIqm9piUJ0UiqIzCUUZbKKXeunGFhyuTY92Xnf4vE
DYX7xTYb48HhBq7lVgTogibKaHyQ5znslTbYc2aZWv6OuzjkoyFn0v3tvlGy+esssCi47C3RibmR
Gzx9V8+TkJJ4PXOzAuGIHik4VPD+RG3MlJjn4R5vZngAGxESV0d+SOA2BzD2eZxck2fE7TzmvDoR
T9JItbWybGJ6DH5AAq98f2woOfEQ9eywc3PCFv6luKGk99H2UNuiIRivf21yUFTPyJypUqkhTl7/
AWkhLWnWYW04Y3pQvnmOhDgSdsAADaXiWZdukHDWCSEPP905gEIZ9pMujmvLt8hX8vxtA8LLc9PH
msR5X0eLmfNDGGTatQwDWic7OfebU7fxsJeQyEl5yr9rA8HEZ3fpQQ3wESEAtAtFigxRVBmh/YJ4
Vj/249nzX4R/P51TZTXeb2MwjKkpKildbzrOzKdb5/mnWLt89gXggmP6dzAWLN+AyRFKsZdI+Wyl
c+rTfkiIUeWNaFgze9n20jdHLSEg3NClfSUvKBjPZgGab/DPGtrw/6tLqRwBYg8Pr5uuTOjIQeM9
Jdiwgrq/XOWCWAXNc73yN2qL2EhnnYtQmDr1PrI9/+K1uX6NPVcnJRROVdMu2j7kPXWkKzvzX3ba
F1pAIgRwID+pPuaGcFXEW1NyYsAsdHlzO5MOQtWs6Ib+Z0mSoR7vYApCFegEA2J9BOEZ60OWLpOy
aBqDn5J3n0OUF8UJ9Qa4IJy19g0cbrKV5QLOXNAkKuKkB49aryTdJVQ1gHA37fBj6fbP17HS0AIt
2tq+KcZAf5fMpaEv8ZhRBjfw4sOA5ZHyiW9L6aBQDrMPbHLqlek9kAUKkXLc6ZCaY6VRKHTFL75u
1whSLIw4Cg/d3NaXGYlDCgMz5/VsFt1kFETxdo1273/i3J37IhaW2lK3SdCMOmKeW1vwZ3Z2XR7Q
eCrhpaQTRCj5q68320fMlJtjmoYs72ltrJwUEk/RoU5I2ttDFLE7IVtUf627qK8U+INRXlbCr1p/
oOWnjMAj6MFjQ2froWSTtbBq4O3etCfk/MMfyRRaRSkHdgeCOPRtWtrFyvthWF7w9uPMhUt/IBkR
FsIHaTFo8BJEO1dZTuEvAbSgB1N4IyigSF+Wy1NYIFHYD+SIVyixHeD2lbhzIuRvhRKqjPpmxs4C
gDBLJvpdnv/A2vmCKiIj4jpN2uZoTsJ7NpNe47sPBi2RfKXHM3lMnG+R9ZI6vZWPwyn8KnJ/MHq0
u5k7VFfI3CS5yx2npIJx/OsYb+Qiz3QpfjXgiyD4DSpWVnWaFO9CY4/G6ivNqrW4eyFZiAqu/qCD
E8x1MWixYatBn9e+Jyiqa4pDAj3JucY6kmNDYkXFO6uU8gFnUWq+4xka9k6aBlwSUpAJMHE0WmAd
vtLlfKw0aalH8xFXvyUx0cco69nEVotOFbEpUiWup+y4o1y4DEziJktkrcqFkNwjisR5SGUDaEAE
LJgZfMUVcGnA67ED6+WzMBIxXuYlZjh8tsrRNT3aDtFg/E0Ky6X+gGQoJkeNNarigXaZ0/WzjHUS
xBeQxPvFtEGM7Ygs4WcrWHSIq7w28mfotDpNVfyWf76EFsMWosX9ZGr4aC8lMyUapbDMSMxrI3Y/
hPTf+4QZAvw3S94mUjrDDq6yn59Gm5y3hACmYR4tdO6DHMKlX7y2jtrNd6AoPsFJ59tuTxm+TggU
fhUQYpl1bEjn3FVbZsrVt7BszXGydtd2xJcgF/8h/sTcPQ2vOuwL275cPPuj6NnwqkayngSlWZ1g
T7UaDFqdbOEDMphNtnIXUGuB+hzw4OK6qxQS2DcgitfM8uBUDFFmtfVXGTvRpJ3nXkXJRqZQ/iqe
0/n6ckX+EgmNdMuNbiiWn1HcEsQ/9+pUxp9+w4sMF3lKUSNYddS6NOiwgWfQSdyxUY/09sHHu1yZ
jQTeHY8QtioC4YgW+2CWwTkUZp1GIe7xPWvviVOAeOGg9B58HgCqZKHxeqPKlQ4bIVUS+8EIJSZM
D26JIiYo4kGvY69fH6Xl8JK5AWi4sxWwKL9eHMydRvPv2488R84adbR6z9Ixon0Dm/3XX+3egbu3
Sf/cv0wh/MrrkkYx78+3LaPgiAkiC72w/S0u6Y+i6l0bsOuBgDkyhsbhFUL3EyPytsip1AIi6L/M
i3XZQo6xzZPZWIDeSBoq64s+00sBumaBGwUgwegllF8lsUB0acWx83PuONqpM3zEMYnAsYNIKsr2
WMDRY3ugyIMb6YzmKEx3EMzhl+J0j86rT8beQynOHh3qK59c1v29+b6orjKBbt+H9moJkLE7feTU
dsJB3LHmc6K5P22/6G8pFvgOwlWpI6jE58xm1tkxGVOprpVLj5KuTCZbNY7CtWBIC1t5fU/yMrly
UkamIurbMU47A7ejjOFX2GtcTYrBCt17fm4E7EHh79uCLyzU4YPfYNHP1vWh1O6w5nMvsLHGIo2h
kRE49cuWXx5RmDJTRNwbTJystlxjPiwRbS/fjanot6ye2mXm/INCFU91z6mI7uugNwqUkT6txzsw
IdMdw6+PPqqhCYZo9c9vwfneH6H1++yApKxJHbCBjm8ljuRUxR3ybgt22T5wXSgmk30lK4D9cta6
iUwllodt0LBRbIxafUI/DajjDGpaU2uYKu9LZn0HvGp/MJB8Ar37DAn2gU815WJEsIE2nrLa7iyo
/uu49wIQjBB4PqzQqmFEgSDmg7El92wx1kXi3HrsmAZv9CpawY5esRVlXoqODdGC/LiXrPqN/EeT
MvtFpPfrnW5u/CsK9q95wSEF3j/ArLgbmzY/7ZuBL1jBB5vZVLKrFuae8rO3VauLPf8xUvnyPV24
urG7PLi7SNCNC2/juG4QC6xffD9rqSlwC4V8sYMl8lFwIH5RHVbFz/oBny8r5ltZflYR16jbNB/C
uaAFbGvnQ6Ya/3RVuX1oZOtpzto3cGLYdhp6emW5WU9ygbPUx8VsGlNbYLUGyKf3qgmbvnCX8FkB
HAXZ6CVTRI9wCb9g8hl7Zy3z/RWUNTTCwwVkukC4SFlIPTx8sNQltENw8sLTul5mgt623Q9ehSig
t2ktzFhSrylV8mVYiDBiWLVyJBN5jVu0+qwBFPYI6EZpoT7ioOviH9M+uCD68IgqvxSzOUfgiDKN
xJwmkPYuv8AsKxKYXU5+UkbtNO4Uf9f8ecaa5SfQvRY8+TSWlxLiTnqtpPCoH7r2T1696dHLcDoX
t+eZlyGAuM82wYo4nTwmX9qFP2w5d7U4VWshITyAkkHDpheIbORqQ1ieVx/UxGDBAaorEJC3yE6+
R5407BFZZmK7w0hE8vOypD5P3/W+J+7Oy6cGYXMr5Lubhu8+Fz8bbyw6zuLnMiPXJygCGqsXoib3
KocbHomr2xMbJQNdCY6/LAZ1kXiOiEVt2Ox1p+9Pdq5Wp1RzhUoVuEBHqb+0LHlG7N73OLIlWh9x
B8ANMq1LZ9Hc1X3UFHYp7cWBgHyOWTBL1YI5kcZdveZWkwj8NM/99V9TtP66EeJnfZLaEuhnTHu5
iMZp3UQnRZK8C1ZsSfPRBOfbCXkimRrAHvv8JCpRtSt+fiFzy0FTSbUnOaF37l7cU8mXV3Jdyp2r
VRVvLL0xL20K5NEO4tpzmkmFiVFEXel2e6K4JxfY+tZA/bu6rl3ea/mAKtH0CPkNuGiO93F4NDbQ
8r9x9gYH2wbdZoCP79cD9jblYyKAyxFgXg77x0j8u20HvjpOdKCJ2mPISRYnm2UiIHD1idxKASPp
nJ1Hd571QPnidr8MNp3Pn9lNxqa8QHKqkKxcomFZfDqebknEz/loDrBpdJVy22QhEy65RryF+Vbf
cJuSUClvAeIPcgENjLRIdBMWWUOuvylqnyz7RTkWF4TBIVHiVpx3RCgOMTGt4IgLmE7sCv4PXSOi
2LvpLMz1lY9ISrXKg9Q170/Dq9mGCHlJYCYGygTU8mPS1wK3vwXaKbxYnyuXPudwsdwSiuxS/YQ8
n2fLZM9w0wHtv7v0NXccSjNegkMtjjmwJU4bKKSt+Tp84qqDSBCfep3uDfrSSuUco7thF9xNR+5e
WhtHyFmHuAUKKRrMDrjEkLnPAvkkAYuheJkG12+RGVA77l0GvebiHRMGr/tIIG0KrfhLpDbn6b2/
xBAy9+wImyNAOTIfY043b8CiBiH5BAGxm9uD27enlxxHQichcSNpGOcB7CHQ4CPiOYa2I4mzlo3m
DPWLtpaZvlOPi70DAu8DJSIsk+18rrJPVcI5GlytXYlOvRNCwH+gJ5zXaEofapKH6P6ReD5dRLCQ
rU6AW1YTms/0rndT5q5e61ulct++aq9IbrR7jd0Y6oD9YSxQDlBRUjUcYwZXknnSSgBIDdzH6L0R
69AKS3QlBtXR+N4KO/STh6AfSJsUHNnpE3wztzDdwieovQtnr7BewqDwx/6vy7P8jf6dSCpxPZ33
mNjoIsGanuwDWcrCumstpnoT3ye/cAd5thwCop2pmt1gqM97r/gRs32toFCCb0SY5W4O1fJHNP+T
BPABlyKV+Cu8/a3up16mTDZ0Xe7sd+HK71Hvg1WBimDUFTkvsUeJmn9Az/ant7n/ao5kxIKaGByl
HAsP7uG96+AFEitypJ3N1eWG/wbduIFsQQVjw7+bQqVbEBeRmA5foaxH9JNrX0FOsw55nWLxINHc
NyKB0b6zJvuyWU/3rbZeppIojkaeLKKPWsxtqBaXWcHPwq25ZDyyKoEY7ljR4yBwCh9QtXzko1WW
7/JdQCwagNVdBUnO/QctF7qMveuPxH95Wo5r3IMcDeny+f7WpMqay23Hf/W7rNbd08wqgTAbBBbc
1/j0deiHZB4HYdQppf8EJI/4NW5K/sfiLS2piCTQEKcuOtemZWSGiVtzWQzJBfJtuZ8UeVf7nSQF
hwt4Vd2GtC9iZ3o4FTiIV1qchwLqaQyNuUzqQ8n9n9KXbz+OAEpTxgCoLmQhlw9nDlypdrgq+aJt
DJCKACICjDqdrnmMIlokaeYVpV3I+uneHaIFxU6Ipu5+rDSLN8NsIwLMwUpUYj72nnL1P58iH1Mu
N7bYuJuDRQAOQJDNUbyl0Xgd9vM2JVyNOk9J2sB/xLfh7c9MRbvLNAA5CwMU8v9sWOxBBExSuuAe
g2sNwUaiiHag8x9+FG5fnW8kBzSAXUuwiF7tgL56h8jBod15yfTkqVltevDqrH9NzRXAM5HQvHqd
Kk68pz93tOqftZC4lZbzBp7+wNmPaXsz48lJ4rAKTPI0LQjZcLMX8rjIQQbszQ3z4fVrrXFGxIu1
E9hjAVUn8zbk2mL3GN+Xr6x3pZPENKd3owtB/OiEPUly20rMybGQKipC2zjMEv2OtcAnLVlvWXL0
dziYUikehLZ8Xn0wmdfIKFkdPkwR53mO/d3FDOGMWYdb1I1euRjx5nGTVX92wjwSJQZNItTIyVaG
/5c+2gdIkPF5BKPSYcAuvcbr/cIdpSZ1GE3RRcsdKqvxzLQ/NIWss3o0gMRsVCY5OfdmJ/jz+QAz
qN2PNFdJM2mXyLwzdymLYh9C5jIJWJhxKAdLmPjtsKyZ58GU8qrR1jvgfyXRXl4Gb0fsMqGZy2w0
1/KZur2fxUaSeY5PT0piGuUHRo1ja9dI0K29YnrOzbWRSg78nUmKZYPRJu2DjFngwrrLL8iKeg+/
7wkeiwHZqfBcu/D0tdEkMSJkGHOqDDlM471QfU2S5XlxR6UZYYuf4qgLbmVdDBYj1qJMRHIK5GwA
/haUI1so4hY4pfWp8p1a9vRh27WHdhzbtvA8Z6x1XyTdpvtBK/l+U82G0pFtHwfDh6gtft/dAazz
Cr+oi4ZrkrVpWEdoUg6eY4RNBZwh5Fw+eEduIi6p7xG0lvr3OnZ3xO2IKzJ8aRfYo1WySnFASC0H
5j69UY49xIuEnuJ6DV1bmdDjlLNyg7hTRm8N/zFvlpFM4F1dorHRSNJSI/c+RrBiKSAXqO56EQf0
w3r+1KJj30WwNkkENOngtV52ERsITcrZEkZl7b1B5kjVEgkHVQJS5tkmEKIp7K8wzCj5uVhz4vk9
QqA7x2+6LuyTftm4xpliU5AlkEG4EbXN5mT/f0s8xffBzQmMPdWfRij84q/WddDnuBgjp0St3Kf/
QOdae+2W3z0BNiogt7u6EcpcAuak7V5NNeTFOixL6CG4+bL3JV2ED/Y7btmvpe+79PMM1HNxenJT
7TsQp3JDJ5u7rA7Qazas54WJex/KvKM+0liUmhrNa5f7V9nfKCHH63+8jzW/tIAx9YYIcGLfr7mt
z/cS1iZorsvPHtlbqET28osXhjypD7aFYyFf8axTwKpxTxT16r01XpKkh305C42rdvfwp4yuDp8P
y+Tg6aAVpu5c7qHVEuO59gVEMDxBjXN4yQZpQHwhc4uw8P9pyXhxiMS8hrqL5tJ9ivi4iSVQYqjR
EC6jM2LeAWYUL2JvkfrEPT/Bqbuy7Hd2tETy2knr4b6P5RIK3LKeJi0ekIE7Gvtcqf6DlPFqBC5b
8SRO9Qf0SSecOl1JWGAcKFkD99GIaYTh+pJIvTKOx65/ORr3ZDHb2DlkW6aL1z1XotmM5UekEAKI
nz3wOiOtmsqBiHF5uocblkETQisgzYlRwmDfvxg/wuXIbUeiKVZfNfojUh7jySmcwWOOD81n37K/
lmh7D0e71uDJGE4jZZyQ8YH6QPnseNH96pBzK0JODFSh9C6hEjEEuHElBxqruOltwrweY7p6YSTr
sPj4d4UhmAyj+ooytNM4lekPvUTftObX+jOSOO8Rs8G9vC7faN8JSo//w6kckyIBMiYVdKzoxQ58
bbfplomduw1VHQzPnJa4+vXJVKwH33Nxn0l+tXlmdAzx7PmH5KQDQuOvOb3mdJURCU4jqBl/7Rnn
hS1/bDM2SCBVDDF7cY6jZsINxxl6/9a5UZNNuWPPECSVXvVi3d1nIjY+OmY8I0Vk6frxsjCv59xV
s/BIvsywHSu+ApRMvj/RAIqivIJC6KFqUqpWEPPHDuB69lDtapuqaru/yOtUSyZvZRTdzlFehyep
CvFXnjzvMLBX96/2S2sUYdNzH5jWBtNNNXROI7P4uPbP6ehGMUUKnn+QdLEmL21sT1euaC6HWbT3
lzc5PsNH12hDcdKeMMMamSdcZ+s25/ZfKK3YTI5hudXFYTXZLFM0HVtOPcye+sXWqPDJOo+08DVj
gOVaxkbsX2VxJXf3/6f8foOVhD3/2gZr5l2IvcV9zuXnmDiEw+rYkyBv8qCZKEL4WzkKdVPvLUxA
yjrNTBWthfZbOS63qU1bHlVZMkHqGKf85we2tcCI0/9QZs0WDAgxgR1szRfvUHTR5BNuQChl5VIg
75Xwz/DTSoOWavOLmXNYclHv1v/FcGb9EPmIyiBzRJujSSmhCUF5TjdqiExXiPSQfrNwl7X84CoQ
DZ1e9TtELsyn29kz6XCcueZjqkDk+Lc1wmpeKuu+LfGRnDyVyVK+ebFgLG/8NdSHv732+567n6Us
eTys3JBLm9G3aINiDuJaEqYxsuVa0RNr4DeqSxVdNpBqun5/1/UF1RLQeFaSdLu/ohAhD7xxHH8s
6BDcs75ktIVMLawwWPF+S1+2LOeU/Y+KeBDJiDr6Hy3dV56yY0SmooZ/4mtM5OYU0+B7FpDUykxM
k95+FHWBC0uCQZMMASz4Si8gpH5aQnwWWfocokzPgUrZn5EELzTBgCQBAahTu69tlBL3WUSnmqI9
9Y+KpjtKZQvGbjNhFxnNSz9Alo0U2qq/6QyLP0Dmw+4ikQF4qvf2+5kWqwk4ybjzYtrinA45QATC
W4uzGRCxdbC8HxH3bRnRCHobKFRVLDA1UX7Kn4jUfp+0afszgP7LnrqwEdMk4Ipgi6ra1PFWHPRo
4B8sRsBup6AcdnmX+1lriicTyIoL9bYIctdLj6bOZTzaPw14Md0u/TbmBc4APxDU6yeoxO6hedup
XG66WwgqoVt2dl75/i4g5HfmyLApplcvuknQhz/2ne2VxrAo29tOY2bGuowntpyZ1s6rbjV1oBAE
YiF51kHLiZhDnO7SiVE27QOUo2o4T/F+ZiXp4EnYoKwxvuCPUAH5OCLDJ+pH6hm29RerYGJlwQ+E
3WvnAICqbp0INmGYJkQcFtm7lP823FhMeirtA/GcO/4Q9JRNHd4CcqqNBH2G8Hggfm1Tu/ZxkWoH
WGEhHjo4NBGusq66nDKQaj2oJhI3phPn1TB6sWoBHQB9qFCSIyFS74F25wqju6DRviYoQVvcGkpa
eg8B+wbfj9xBSza/hfGQv/9NtJB6+LeeZZ6dL8uFmNqztbiJxlUp67ciEaPmSkqUlFwX53VeK1nZ
/gV3g24gKxW8ZgaJZXLpSRcvZ0gLSH1pvFUM9L4go6sca13Qq+To4OjRSnWh1UsmadQ671OBtH2z
Hjuh9RsA4qOHcEM5VWPdq1C3XgHGAEH0g0J1Nn6zTpi70KbV2syV92pVegN+tsuLl4onk7h4glkP
/h1Ps3O6VPwFZXKQnGijsA8ahl5Qekr51AYLby4unU2FWUY4QJ7xWRHt9zZFDwJXasW6IuxFGBeL
XMY2ry5NCqDQW05v7w+j5KtL7udHRfV5aiCh4HkV8Shj1ipycUGOP//JULRxdltCnVGQX/R9WcWZ
UMCOWDBAUlnmjD/gq1KUBf7D90RJfD1KOSGvxYKaIZ6TAvALd97Ie8VQoHtRuvbMLVNZr27krkbQ
DXsx8hB3RCwVZW0uzba0i75n5lHSoL/R4Mx33qD2dovGCRGV5dmi10D8JeIcBOhebrshg8I0KqDT
PpKSxQX0vPPyoTczk4Zxlga/YC5OpmVB8MXlsfrntUnTyc4bVVaY/SKs3zTRo7oE7p9KlXe+0zfB
U0OWJhWAnMBcp66xsGbUc1Nar4ymjMJsApqnMOWIxqOTxk2Qh7fcmHZ+8jSCDiClcATrr39cXt0F
xf/lrxjAn0DYEGubukB0lXzVw1Kn2Pmz7O9aTj6fpTfXHt0QVHi43JIl/AK4WF0EbRjpDxwGF5Iz
zcrIKNrACfGOS/mXPkYPh5DX3MHReKOURs52/RofocJHEzabjrtPfBNwp8V7zNHs1L17sBOxvnct
jwsc2zg+U2GXvoBPyojdR+fGDD76UNanlIDXR11SIq+rMDaksMB17j5YouORi+JV/BMcRqp77Y7I
iqil8zxEruEWDbEvzeM7s/UWe7XykmQ2L2mX06eBGFHgOsmtSXGQQ1uV1WwslE7RM/I7LW5kxCiZ
wAPMttopYXzGVZuQyOe7CtmF7kLrPZ23pnwryTjQRcxnNoO0vnOHyhrLqgf7h3WNSEh4xpUE0w91
rJFyu755Jf2d5+9TC6XX23F5eQD9OzR74DlWR92XjnHEeIQpMen90Y8dzR4CvUfTZrLlbgqFczAI
xnfb+pDEfXEgHQQTJHfPqNFDR8j6iA7hy3WGg+2pTeNMoxQJU6Mo2XR6n7qLJCpWUdIzJiqeORHb
lqMsBZmZMTQIaLTfdHtmlbYZfDV6Yy6ly8RkfKdAb4Z1EXiSt3gklXbZfWCBjpylOtAgmw0qJlZR
IFcJZjUAfvMfSfy2w6OJnHHyOgL+r6gO94x44YItDnZMKkwXOfdGYgDteNJ0BQPZ5ZioXo+r3g/U
RbRqIjRneVTQKN3ayl9GWi8NTZ7xwxj6/RlskBYAYjVS70sca7YWgm+q5FR1XJOs1BrkLqtcTN0U
ZUf6Nvm3Oe4QY9u3h0J4W423AASCoSQ3M9inf8SEd0P7OCr1+xalaNsvgPjUeOX8SrKNe3CrbMVA
D3jWJoGwhLdZxwz6K6FDnLJ9+36jKP3FeY5SCfhgpvfbaZlusyFSXvoMSD7H+RFNiKfdAO+3x1+w
djDU4mneY6tbpgL9DanycltLy0Zo0X1tADZf6Gwsdb2hEQOM/EPcvB+19Pj/qPEC8gkUo74mZN7S
vEKzzpsbBK99lqmAoiLGP1d6gpd9wyWawpZw8uyHpAleyNt73FKEf9efNLw/bu7vpXF5/xXbIXrJ
JEMXu/w3PtW8gi6B3RrvyTRt8Cw2dPQTlLdi+fHFXXNxevwhuz6edGZsz/P9FZU/a2TiDyaw5Ecv
Ccj37Rh7h4NC1zhpSuHg4cHZhcRvZxbo9byLfQtZxSW67Cx7t4QO8LUKJoJXUnyE0IBTBLJO9e1x
e5I4Hh2idlVOVhf6HXmgXDdcdOhwzm2wCj0TaHI+wUBYqQd6pr4qwDZKd3bpeG0pYv7K6JnWpAtw
Nvk/qZlzQZedxZHiWerfsX4pXQU8VAiyt0MCIszwI77fv8UpWw0arU3m9v9nowtKFjEE4GWXize4
Z/9bEPE8AkoQ0RTKrKiBRhYCZQLMV1GCXKg7ek0bYmO+p2gJyGR+nDazwj9YegoBrJmP72fXq/4R
Sd8JE8Wz2LBI1UN+Yw4qD0kk8ERTRy8JkBs9tSt2K+QlsHfvv7YpiwyNBlHYHGsntTx5ZLKr6n//
KpO8Rw7PkyWXdsomJsq98eIqvss/L0cmHTrxbaLZQIHFpVSHkZ/8jHyFe8P3XZnBG6C5kiJxzPcX
6JoJ7ewhQwpX9/REJiNKls43jCsu8eW/wJJKjYpV3asBXnaMBYzDo0YZzV5yMSHXKuUQVxzbXHb4
1FqPOgwM6AarQ/kYKrRMwgWHQPzQbM/P+0cP4f6mjs7tnzS0plM5BLDI+MhXber3YstWuCDY99Za
fCRSAWRa/visNvg+yxZLJNiXTLtCTC2nB87lyY3BGE7YX4oSHk5ItU9+aB5voMzh8FHYQfq7WKwE
cWwe8SMGbefwOKguEX8RUPOw600/+XAz96t+1ANH2fWJZIMarDBe+dtjmaaxZpee1uBpFLY2pq0d
9AC+fpcYmm4BPppFklK0ilRb6b6+0fCvbdr096Zkty6dV+l172tyRBjFJ9hrZcdTfH5GyoEYckHu
dAc+BQQnLH234pAPIPJROR0ypR5zFh0bVUrotJDOSrIL3R21Ss/4P2il0z6sn5vJF+6JG+cMTLoa
eNAKIX8LrK6UtJf3RDSKWO57QopCjKg5f4pZFatouEDk+/3oW5OuGCeGHccayipG6PT2YVTfLG9i
CfDNtgkqN93rBVivgMv0s9cQjrB/BvgUETXj861Xlj1uiRI5SRT23a/DHunpSS3JbsYfIHuvnRY1
LBpbwHRGinbw/hfalOUSN908bBjAXRkeXWSKBXAFICD19SZKGarAGcoEUZTPJKlYl/SEKc7Qo2QX
rWOsbmEpM2vpOXSZ2cLQgdaWCffC74H2yfNFhXxAYTSf6OqkJWUj52kYEwOhmZwePIhlIUrQcoGw
YzNBuqUl/cSI8Cwv7zt03HKt8rN+tblhqFwv2/mUk7HOiYeCeRh1du4azvaBfmMJ1NNYv24EOUCT
xPDPv8bWy83tUzbsiUzw3gOEyMPK4a3j+fyEJoPT/1U2hPzq7reoSCNVBs61oC3tGh96iyrPmuQ5
dDo/3hs44QY3VxA7MrdqiOPv+LfS/Lqf45jb8dy1FWzVpktzJ3iBAVHLhZ8ZmHws6QhCY5ERXgat
TAe6cK0dSWsiHOtq+tNt6nrKnlxYEXrAN1oX1RV627VPrGJAK6gE5d/1sgzr51YjtV9dQymZghby
wRvP8psirKCilwlMEj1CWa/H36gXEeci6xHPksKKO0gOg2ImrHb7nyEymHX/t+dSP3tWmlEci566
e3yoc+j9VsaQa1qjGe418zeTdOIK4bjabscvZ0rQb6N8ofeDCsKBzfF2fXOT0NiRflR/DtIHErv2
w5QsIKuAAUAoze95FWuwIkpHC2LcKIiiPGGdovNj1ni5aFriwOBiUk02+jbpfLennIapP55FQUtc
P1pGm7x/TVL/fZRZ+tLKmNpIgygqs6D5h6KejJ3giI4gWKkobE2dppFgFXYve8wRaxi6sxAy4SPf
QZC7r4i3YfHO+/cFWEr6jZAwJQStXKED408Ymc+/vBFlwcdkpHfOGhV/x8cEGCfCJ3aBGZ2IddZJ
wnWOQ0HpbYuFFcCFD5rBt9rclDmsgklcPM0kNsVAlBgTvOBSAoSVE+C+oap0nOsNskrbJk2wRdkI
T7jNLZlHPiQ1/9GTAnrgrCTWU9bR4uh9diOMFgxGK7yXzwRR0Q9ZKuKZyjC4dMqGTHEwReJ9hicR
jgYmo/SKX2r3ou3D0e+/FONYdsQf7HzhyBTigBjqgoZ2xekgBYgmQWLNGGQnB1OPSqfnwmEY7Gxr
EaA0OFZcT6m+och5usutB22E8oLVPtB4ctaPgo2GXN4A+RY673VU9MFc/Sh+89QxsQGCBsjJB31J
pD9rpq+kBeQZlwJzk6J3n5MSHyte0eOlEmFsALbcoET9waFse6TQQjZyUYGcO1X74n5+3wqVFWwa
k5qpQd8IP4Celo5KF656hd3axA4J48HH41gzmZz3yFI8gWB0JmmEeUTzj8EXKodIGj9Aowm/a4PD
RdsZyPOaL5nOzcKKd5s+2/iQAQGFLODFog4T4x6X/09dUibS8mQEf+iy/H93XdSGuxADrcTMQ+73
d3a0fFt2hoPwD1mFM6KsQtQa068RD8o7d0jZmb52KxNZDRTXTT825EQY8txtoDQbYsq71zJueSg/
lkAVGJleoe5sLGKQJATyDwacFp/hU5Lsrb1kGQxrrdeXJOChEmbOSzQlS1erFunikT5uSz+pGEZR
JD6DsPMEOTwe2wWkpAdHbGgQqe3oc7QBA79zdsyopdb85pSAiy+sOtrBug4EK2nA05+unNFolJMf
MxbcxMLzchmM6tihkHZxHL3c51vn5ig52LxgvFu05kgA+CIeO1abprkA3ZDiD2NEAJVwtByN2xE4
XeTAE4gBKS/j1EOeQAWF08tFU5djJyTgnLtLd7uTdkQyN+BVFgmEGgRf2AWVnGrOKwTynmyiGh+0
7gwatlwuCs3hw1cJevmvcgssUPkRDJlOaauhLKqlVK8Rjc4im/BegIDBjwUXqp0JnvgRXwgjR9ej
+dFJfaZWvy8hJwe4DXk58nNddtaOaJUnyQWzpn6A5d8SVTrzv59ULev+1SISGsUI8+PGhcKwVduW
CZc+ib8vCWxtdWyFLCZgJPXAuIj+MYASRb6SMZQKQNmd8W566MSsQci7uWoOS7X97ymeqRH0i14o
wTwrB1rqstYBB/3ddx3nMAShZsoVyqimTj/8qyvMiVWNwEMSlxeozabY+BGWhLwoEWqEq1CVai7t
LMXaaI717fB6lOkd3Xjdt2tDcUnyBYqLaOgFSsdxrvkvNfCrAfmAOYtqgl+jhigdD8+wXbipGtIF
fcDtA685xl4M9Ty1sGeefs+xRDhS2fZbCE7QO3VkE30wnhReZkKsYMDdy+AHRbCzvmDRA/IQPTzr
6fi06k2mETx6RI4L9sPXEjDZja8cSJ4aK/3W0gpaptcGclanBi9S5JKUkwLhAGtFPuc1fNRm/omU
UW1tS+ZqTEV1QawqyC9f2NInt3XRgKgWiwFALOATTa1COXSzTp8Y+zrK53umFjy384Vp0pzVSuWm
Q3FdLaJRreNBWw6M4IVeCA0KmX7GwfGWTOpvZGJh0Mu3EoMyOhTb3u8CsBwsoND3ZVGeQ0PP2+q1
hR8rJMV3UlTcbI2u9C0o+KSGF41LqLY6jLWSRPKQryKyWZcptXBx53GUESAnlIzOBwJAvCI3iPlR
x0eRb/HLJ/q7ZhTDH1MVWBAWdee5nftK1klUcKyumVx8j0Too0z8gwO7jr9UVDBgD342MhBtE3sa
BFaEzSrZesucJjvMwSwE5Sx+y3DYyfb6eqorhUUoNmERKw4DM9H4Tv9a0y0lWnWkC06ZtNAai0aM
clHP7OQhowGsucnSgbbygwjuEIWpVsW4Ti6WmlsmrMhFVjgGt6jb9fRQ8I5uqpvmuKw+vYA9qJql
VU0x4adEHwaPsbo0Z4HKvvRSunBBGpLvG548ELVOB0gLsejWiEhVAEjILIN7Yd2y0eLgSYzToJd7
4x46rjvS7NOCWnX8c5a6ebzeF9qNwPjMp3rSwOwrHjfZDxEvwKxvPQa2xkH/IvJxutuSs5Jpcp70
+FnsKyIDG8pGk0uH3Vb3zJxQC3spdv//U2sRPT40b4hKcVEhlPT3ERBi8MnMjPnpvrZnUVvlxNbj
leDzk6MF4XgLnZB2v0PH4G+IGMa3WQg5GN2AQz+ZyaN6mXtTsD41qXC0LlKDUJhjSTEfuMA2s1VK
53J3Vc52otzO2h6Ggm9j6JPelBXlYfk9XqWS7r7PN0NVeJbXnu0QrPe5zeMc2qi0rEJU5bqzcoId
yalrvJxce6KK4XpMISMggYmkHXls/RkQCtDQBRfUGDFRyqHkwweU5wHNG2Qx6rjoHgv84FnCO0zI
XwXHi0s2eLQjytH8H/Luie2DHhF7BTIUHHkVJ9GWpcf5sRlNdkXqmJXclXXu/bBjHCc/d4fuQXJ4
gUFP/I+S+v4YzxPhlX99Ig2gZ7/xYK0xY3R8LUOxq3JnkdwyKwAhGklSFPp8lkbUCZ6AJX/o1+y7
O7htRPO0P+5EsgqlJz2DVjZmHebsv6F9M+s9sx8unYAn2EnGC1TOmfp1g8nDUToy3J2x9JB7aRSY
apXF0JEA1sHjUamdkNm6j9+X5QilXsRyDQl8GEEGRlDINH1Ei/ea2qMxuHBy8ut54AK1Mz9W2SU7
6CHoEsEehxIrIlcJBqfVCFM4UE0zJ7CjCVElYJLrAKpY3lCTNAtu8v04uLBtVb2ETD7vDGz2ljv6
cl8tc3lTWXu/m8VXCBDmMP6ORNVNkfivsSHIWeqnSI0b0p/PUvt+uNG9R6PjCpFZG9y+P/P3D2VZ
2Z/D+tJX0dpCz4SeuwrySkfhdeIkgdcV5m4kdQXvihytrKYHGaNRkYh774IuHLmVIWiXK43Xuh1z
YaOaVABBjLlxzmzOLk5KnltN6+9sMI873Ioo7XJSQwPvG6Aod6W9YnvaQ5I0w5o7mOAsNeskheLb
ZsLZFmzKge/ZRSNrSaaXyJhaNT95daSWJlDghgXt5CBqSyIK41/8DBcDFe+D+/7gXiPxSOPpqq+c
y2nUCXHvdAAt5K0vIp8x36rl4UD9wRDo1aW1OHll/UUx6LhjzlHZf783UA10xJWmOgCg65TZuE1z
dcK7Bctzf/o6KVucB/aQefUbDvlL1BziHtE06K6jdlIXl86P3iu9R8S5W0JRsU0Zv68p4As9oUAW
s2YbOIvjz/WWeePt9mtldfDJmp13EMduW7fghyAKzBPzFUbC06QcmwwQD2Dt6/T0DUPkpS2aG+uX
eDvAfiAdjG88hgAU8IVG0ttj6WNQAPaK4L0v0HQA8SocMdWl329Y/jEmXp/XeDLQ5pwsjRryip0K
Tv64PxydmeoT102TqzHeEgIZDHWWj9iuFhvoZJoXSIamdGhxg1o9bxkgbLkzZhglT4QY2Azg5j/q
SVjU/0QoJ/y7oH3AkNlOByrY+PUKVpBURWGgNIIlmvSzPIGPiImXF+2FeDEkHlNMLrNS4aUEmH42
fB5V7Sbh+jmfyLFq0K19fgkAhq3OrRv0gnhKKmgohaLGDDI6IBwviOlhWrcNeOQdQmDIkZ0IYjRT
xFnaGdER3R3CHJ9acngY9Hn54s+lWft6e0LZdZQ/PfhYYE4W6/eqHkbtU7a/oAB8ddimSJvU0TXY
xigRzibHDqUiUs0vy5F7/ppRD5u0Yxnul3y2p01Y9U6CZuIXx9XsBEAMFfj8Dc9Ybf30ZrLlY6Nz
RkA2Qf7b24yx/1b3hGWHlyjETmiKRJsmfZz1WdWSDkZ45EPC3GLXxSZ9AAaR7uxd2X4nYIr6wv+r
y0MXKeMqH5K3YT24tX9DionIXzbaJOgRNVjs0N8BIcX+rZNEI+Hcx4tJsRvMtaH5N6YKvebm8pF6
HDf7PICFTb89zidXtRTpr5cF+1nbpQpdKA0pH0kQcNrL0fwHzeIyJm8h5DeFyUY2dpRVbzbnP/Wd
ZMsdDZfkaUL3oSdn2pAwXUMb11gWBDlU2FodR8mXhLsDUf21lpU96TcAWkDRPHPDHeQY4nj9LIuN
nQWLayjd+hFEy2v7PXTkEBop5JICwxJtKxFIqMvJboYm2VYgWgSGD2Az6TQ5uXxrCoLPLvaG+IES
S1CyWU/M+egw+JM5MDtDQE7qNl2bOOKXz/4vQSb+5maIq4PA9RiBdmhE+DW4MC/rgiWhboI80mKi
MrrZIiavuUGPkhmFRxPtDsCrPcRpPXTIvRM8uaDpwklr+sIQrXzbim0hOilG9o/KOxXqhMNILR4m
Fu/wZ2kcXvK9oZWcnraHq15sopaIMSLdSCNnNSkYe02d95xiMBf/MtLxF+kD6Il2ss1OmT+os/6r
RekbWjFnXBNSSkdf6QsacDQykMU3KpSdg0Har/+NmWe1rN5iGlZpsZ5Wo6bIGGLfGUa/JD1XZiaf
gsxc8gwvbUfFg3jFKrw50Xcl1ARys8qKwYLfzJnNwbyXXuQziCM4guK0H70WXhauKYPKTnCU40x/
WNEXvshNpm0IcaO4WA++3mZnwkwESG+eGNl7Ls//1XpVoS98E2fcByNcN2urBtyA8uulgnPYKaJE
+DCboDaJ2vl5zYS3k2+wVg0KDq5iRunbMUzJjKihM1fgp1qpCAY1ZYZSVudKwAcKZXlEyPNevR0Q
J9jr4jIRow3zH5WiHBqa6Xkyd2pWEELVfK69Uek1J0JkAWZj9GwsijMdSTIK3M0XO5VIA2vs66PR
KrI9BWvjuP0cO+bai1pm+IA4qKrLOy0Q1asvx5RmnwuZXYgHCK8fg9Cmr0TDnu2++mrcYSsDJ/tS
Dd7ZUEQ+2/0aYf2SUIDTZwabOnWizaEJYJ1hijvmLwswK1ZO6N3pCMMaJJxofdazUkrgAwWWf0pX
cS8qXLkNc34d78oozZlji/izggv0Ije3dqLM97u3Y6i6pbSFaYrcMbwyXU6+LftXg0AZck1HCrJK
REUJeKzCM76THP2nDfL4StxIFn67ODuI3wECTenxjY50Da0tHihTeKkLj3d+3spau06Mc1zs2XbS
rQzOgstVXP6//LiyBPK6hDNuHzk74/zePxM6J8y5i6qQkTmuU4g2w/GgbysXxrts026LsYTZoo8I
+XwE9Gte11UKU6axJOMMkPq3kiFIsuepotmdkdLNZGawO9nT+edpAlbFoketCIUr12AblC98RuSA
SZ5HpLwrZk2iJ5PJeLxzv5zrN5CEBtaWcPb7gzMwMySoAbBFnk7UIi0e3UyoMAIXNitQUOUgwhUf
b/pSKsbJe0+3p0LJQ2QlxWJUeC5DF5RowmwhEzg0DAzbTYIlk/FUt4rXC/WGdra0ZyVrdIfqFpQH
np4gGJNfd6kjQZQSXuC+/sbKuWhV2QIPlT9sGNs2cOuxiZmw3Erb/ULVBzLUKMd3LrkmWUA86Tgk
uzejQDkrV5Udp2EOBqu3B3/aL5UvY+gHWF62h5SotAtwnAwGeU5qzw1lVhbVa0BGe7DgTdP1ISKq
ePylkGitP0MrQNKUWUsX6NXkj1m4ludO1qgAZW/aPS3rXabtDhq5ZzQ2MeoIjCi3NQn45S4GvAub
5/iStQIwsGcVOP7dTjaGMn+OEIrQ4FhYKCNHrFleo77bFQ0EFYNChOA/+qxL3ltptlggiKJKB3oI
GMBqmNNwZdZ7XPEPAD9Qb5U+rrwGFIs8LVm7mxyfCe1WVKTPI2yPawlWahyq2u3UbFJmZPpjgMZt
dIBaztIvG2uolVcrEKMH6yRXl+xZ7hTRAYHAkvrq8uzyxRw/yFXRL7m5FB3/ltfIgAtR1dymVcoY
JrVMG7XlU5kESqhvz6NlRyyvR/B6YXix04rSoW2ycsRHVeK0Sd8SzV3H8XKJdsnIJ8bM1HOOlNaE
fU2MOhJ6kOcZZapz4HBY3Xxl+bNCcdtdtKGg6CsQDiaXxajN4yQ7Zjet/GR+k84hBB9ELAUqr1Yr
fuyy5XPspTDtq0b/u0EDDAv7mv8ssaOvHFNdbHM/ABmsJWjEyAHmtHylLE0I6x7Z1L8HS/Zp5PTF
UdpKqK6j3zjVA3ZeI1oSnjmISgyG2EMB8WRUfdUgbtJ2mTnYMipFAl0kxvFCs7sao3Z2e/5JgoOf
zeA1odWMMGalZEuMwYlbws2d0G6KJj9HektcaAr7npaTQRprdRkJkRnvbOII2sH0iWKx5gpai8dk
KXHQKjyOHchePGKabxdAk9rjoHluJbdAw1cAMk2DZFgQFigYPaT8ZKJ+PA563fyXeh5+upA4nFER
SZOdSpAZvoXiqzv73AqIrZVAHPlK3BmzmgnfFRyF/syiHoXPLggzDFy49EeW9zkGD/9BA+g3dZFN
08cSrgZKZ7v1why3TdCfYDVkk+sesM2FJoNDl+fuXMiBt6mwzKjypqa7GEEwCRQ0MghQt+HEmdrs
BpfetuM0ZR1SMC6ylhjTIWuuVD2EhF/ytqdURWPAd/g6aNaveS1ad0sPb8vPKQkgipTeNhiIVsq6
naJPg4TkAb6JMMZ2TkyBEMsz5BKGcXzKi0BoqigNqR8a5ySgQT/2A3mmiilgP1bdna8nxcCcrn2b
5GF1Ihz+fh6dOx2RsGJ2ja7+/2AQKttw1zaCg9q24npeD+yVNGre4Pes4vpiGrf3qzk/WwuqUnRs
XvtoXrJu4YXLjB7XLauAUT23aeiG4K3XnXPFMumoPorm5MPMmkFz8z8Emw5DAEUrriTuuRgB9Xyl
13PAebGzX84voQAUjrnue8pXvRTAhA6Xzhs4J+1mm4lo+8g9GYQc4iPvd+uN2xNMHlO9pKNhKYMq
LI22omKC1NDKWlwSr5FxY0NIEGoi7TAvcF/xA8P0Q+8la/elDkC3mM+PL7yLrHm2wJOrUVHtgMWx
teu9wAreK7Dt+kAaJyYY8NWMpnWb6YwSvey9tTQgRCKPO43x3pVcE++F/frtSe6AtPYfGIZSkWRx
RyUpVcPOlPLXVpkixd+za58zUbCgX765V7ggiwIUXMaA/0vzmHLZ+NIZyL+QumySCl2lRFIumrJL
hnH0GRAvOk+ejlwfvnIvZz4ebBkk/HgYHV5N0dewvFidMJ+Cb/4/VfJkSH6osP1q20ZGqGkraA93
kH3+z3FG9wWHVmWDsWfgWhuud/qaMmAMg7uXWs1gVP91J5P6zqRSXJiISYmqg9Kc3PEeBSFLoz5K
h8DJL/9oVBt68wt7SOmwMQynOBXhst+n3vUdvCSKB1ud8PzyJ5YgusLbLhTBUAgF7kc5BowvJYQO
8GbbYbeaEUX9TAKGxJprJiI6zsOaoKujw9dyaX4Q+sz0f0ntpQ3094giBCmNE13sRxDKsE57swN3
l5ILu1dVCqPob7AF9h5gERKkbcqLyGf64Odkj7tbtBWOEpgzMS/wD7GXBEXXHreUr5JMBfVKZwtj
tlzG88ZUozt5uY1drETzaM7RbAlz99UsFFxhQkh9T0dQjVTBzEqhb07Y/9xPQYt9sPzmqLDA0FvW
94NesWEmnKnPOeRmxhe03Z4ZkOLPPp9jr1+E6S2p4sljX8LG0wP7QMY7tuxlvzBTu48w54c1o4ee
fYXmMCWoi5ll+O+TnuvJ+OwG2dsYaG9TDhLyJf78vPn6xN08CNJ5fkzYddWgezqnOiIZVr0ymEnN
46U6KyUevFtisfFkJaFXJ0TxYFrS95zHvhfn76tHRNYVyPyrQLFA/DBTLYSStgvkIOjjnyWPIs5Z
bPvb7GZUXFIWP8Gcc0zP4QZn+2PH053VhSqCjZui8kta9pjJPGPeVaEAsAGgJLs3s51LF3UcIm7X
9DVaxjw4gDDl3XsNybMcJirTG6mr0LWyh8njKVVJaVap6ABUa5PaUxggy79dsYaaaYEuOSQeGldP
PqBuVAA2gSP59drHRTIv13ka6IgqKMqbbbTWDu4nP3v12p+zK9O/eY3i+jQPR+Y2wMsP1zXEQQr1
WqYnBwHzwP+kxrgUGnbFiUIEb4DtaFz+CuZsmcvmOS1ktVxdxqXYJEY7Qm32RCGTTwCkmWp4rB6c
jksDeHdDpYuaAkF/mZJthLS4FAuANYaX7fCb2mwpkZx3mDnAlRSSIdyDLCF1Yp5XLtYIKs4plr54
og4ixCIobt3Hn0cKkAN3f1H3L3IOYw23KZH/ZB6W80u+c9d6V3BeyBfU85QwJnaS1V4dLEXnWANM
iNm3edDjpJ92eO85ehIp1UsZazE9l0Jdw/9XkPdjZ2n6c6GIDAwnp6swirqCa0GcjcDnH2lgl8a4
kvfST69Ao9YB7Wc6TZiU3IciOgPqyrNJThF6GCq/152ks7hthXsE4myawNiViBNGJMZPtRh119qk
N10wezulVHYt/oEpfr68J5XMMark5vKWR9GTfk2l9j4gjtBVno5qQbFMKHu+KUwcR1E9YEb1TiC4
s1jXciQr2eU8Hhhp11KYCfYnw0DjYr7FfHO8+W5k5SyEpP7d5T9U7WjyfExndWuLvJr4Lr8KOR6W
LtRwYJaor7pKJABDZO7xCsAjgM0UNcnMGD+ux245eVNyN9m7Jt5f+nuL52ZzMa2K/dsf36j8qRTX
5FVVcvfvTngw5Mz3Gin6w9TGsYnf3ADdPdaldxmonmbGt0fjIYXpIqwAULmM2ygmJ/CIPAvsDGKG
oRXDXgbk+89a4CN9tR9xrtdvR7l5GzGueTmD/aW+iYVS7rr94MD15rPdXS4R0eXR+D93lvaTRpEO
CXeY+Yr1RqvoMVTenXEdxeuXER+YZOqaMMnodDW5M8TrvbrDp8Fvsnk3VRm2vfRKwF0K7i7mth+k
n6qkeqcKOMVhKRAgaIrs7vKAFHWXZRDG842lAaHoQY4MMCAbcF0jtnk/dK+Yl+oYn9YQZVKZM23Y
bUl7i+E/9c41xuUi9utBFqpK+DmwwS5eUsTHnK10Y5c6NLBWXtKXPouYszvciRuNLqev9cCcjVMm
fdKAMkIrPKQwL+cg9kt3vx+A8Eebzpb7S/g5vy/6PVwdsHrxVYSpg06Ce4ux+vXmPxpMBKWYcler
n/EdSvb1xdnIFDex6IH1eU5h56XS0HIlJNxFq9fEPzpRLMg7ZrEz9qjd5dtpNIbUzIf8ugBG4KXr
thDCNGg+u2W/nIyP67cgryVDZjVF3xFLkW5eEz5afO49Vp+4CI8R1Tfk22fo2JmFom3/6QSnJnTM
F4MoDfHOHStAgnxOc2tkSFRY6FE5c208YEh9yXyeDd4N7yTMKW9sX3+v5w3lz8R6WGiIibZBV8dQ
nWQS2nykpNzwXoYIQuZrPeEHPPeab0M+H+IpfED5kPFY4yqW+x/bzS4q2XIV3SipczaixsLzqXr9
hOEzlIBlfRqHASD6tZXV56SVwAGwYQXUIPluctyjLrTamkfxX1ujb8ekLVrf0kdEPeoW4wKsHibR
6lANaDsOf8ntissaHn9FlIh0llSPbtlVOF3O1d17uitEkmcwWoysjOrQTWOB4D+H0cKNZSGs77Rm
WzaJp75M3KsREBugfwy2etyqoPgFPiqKrr9mxoesH6mags4q3C1AMVyRnG/tk/w9aqN+ElZH9KL+
CUMwtCtFr0in7PJ0P4p9SwbUXrx018/kKzQNfDYb44HUN7lR7gSJEiHLN7AsVRT2ENEUkfIdI8tN
oFCoWqLsbQsekvolwQ7ntL+7Z4aLb38lL6PxW84quWetuZolGsILa7YTBwo66uAuletO98dcTL7R
L19N/4IK5QXr86NXWk/ByD1k07uOXL7uikefOXIEzbABAl2p5RWowtrb3ttw5xALuRGSolufU+HJ
rBcRz8ZIbyjmFSrpQXnAaZPsRuh/PTrKb0i4Um3oavSBh0zb3Y5txjWYbcpDvhXeVWShp6eVNGeb
tc7DvnFOYqdvi+uD99Offw2OcLAToV5KEv93hSlz7KQQrvxjpbWfAlygfzMNBIn+Oh9CPtkIFojK
jIdjpaZelgE1TpTLof4AD/NAsdRDxOr13pkhbLC6owBbf4M+WwaE47XEtNwUL0FOUb2pFiLomKWB
jTwjRbjzbxoQ8XtKsNS5OTAYraaTFJQlWcCHNVZ0pXFGGwkD5RckcTJXcqztucYOTV93bjHP0YPT
lj4fMiYCBsVEDuMb5ljb1rkKs5FV3uF2F1+Z718gQ0vMXYNwz9f9VqKW88F/uAha6gUpDN3QkR0t
AhDQcCerdxx8ThKqb4/qodRzgdOiLM4DBsLgm/zQFQj2PLZsS/JLfI1CIqYXKqN9PEWsQ0krKi8o
z+/fubiEvjrMQrGVqyleY/mEOfco+MeyeS3nmTM5g5u42nSAef0v1Twv1UId7xiXMRsJ/JTW0NIB
W8rRLq84y5xSABgdq/6v1FdYY2WhAF5lUM4ZbghHZMe3gBpCMWhzZ8ldsrJucMcNPp4Wqeiogy+m
2kqlyQ7yMUVXfnbHbKZDjBwIdHHSm4fN77ZJFdqAdJa2fp8S5zPa0ACOTF2GZhQ+sUNAIlmRib5q
C66QUSX9VJSAGpXjizRkvYqEzRWz4ES3iKstpVlFaWoQzlvH9sc2Dn9FAeEI4PpD5bjF5GViDQ5I
+4If1DftReQXzqzKvsty30WRL309KFj4uwRszHmarwncyaMbnrPcIc5qdNYc2facoXtdenXsun9s
8PLx3AYBxnDLsx2gLt2zsYlKVFt6vTJ35HyN/kLpTZ9dzlUUMYBfkcEHlYQng91TuNiTSc41vZXv
cDm8AL1RvcYUUWtmPn3bWJgL0EvWm/F/vHR/uw9YZrCovB9t6r53P12FimuJsNpe145Qimw6EkCf
7ITAZdrhm3ilSdnUBHQ9nSVQUCeJMdZW+3ezExFnCpYJPKBsyhxoMrzicdaEsZd0EToaqjhZSLFL
qL0sYZmzj864V6CPkM2YgyawPfRVMjrebqsaFoPSeRFl08pHaJ2QHkTxvg1jgT+7ZBHlSJAZBDnf
y7dOtsAAvBo5Zi5awLSvOFQW1q3s1nrqYt4rVHBvg4TBANOj1bCgEgfnHrnNzgeNepca+0aGsrRi
/mZpvzI8UsxXR5+tkWsx41t8jLmNMT7GknMlFd1hkNa+++PWwXb6ZzpzSS9xxixu8tTO8ztVrGac
m83HVpNnc7xFlsohaO/Vv1LHJ8ttTEJPGUj5PGOrg70fltisSrM4A6ia+ckAvMP4nyCSDPOhOp8y
NVjrTk3nn+o6JP4lQEtIF2v7phGSVIuoQoMf+soDvIx/eMlsYwNovZL+6w0YgTg4sngIoYPSVXEx
WBm3D22UvIO967R24oHmRgh1iM57w8l7TPVyxLRW7GxhaPwJsHTuliCiP1LUo6i9Dqrc7z0vAWdI
F733GUrDSS5Dxa54FocXBL1ubFgBvCB0lq3nJlq8Y1ZTxL1fz9tL4FqgwsSsxqZP3WxovSorlr2e
i53hDLmJn+BQNq6QWs3+c1iB5rDR9onxlmbnhmjjC94BzJ/0gnQI1gCSE8kvLBGynW4M+/Lw6ITS
UZ/qr3ev0QSqpCC0FDgAt5a06jmfRTzmu4/ZimaCPxCKwOyehOyTW3SKjTXM9Ikczb0i+/ISxsSF
js56SxHhotV5bYUYkP/jVBNUT1OY2p6uryaH5OF0quMvWhM+lQcivudJ6xSqhyJm+fP8ruVLFLKq
kZO1PCkmf3AGpEN841yQg0BqKKH3PzGBYG7YxdGEJZ5gzjnVfZn42HTHR0lMnVfqFRqIXD18KP1z
PkeA499ogBtE5Vwe/eU5a2LyCp31liW6YKcsV/bZamyYUKoJyd7zIcFpaZnS5krObKsIETo242x3
CHHMvW1RrywqDD+9x9cDdIBYl7FWVaHflV6K5w8+n14dChij+ktMW0NtbiebKzIKYuCrdpZp5/Wi
L0JrcXRc765WnXPo9GMExWMNzacqn9RPCwqhZR1MPU66a6u8w8bMavtCFC4vjqqrz0SWmrQndIYU
KbJU7NTrz6G3PdRWFFdYNxG3XsceqQr0E69fYDJazBJ/xTjy7dg1o6yOfCEw7BUG+P9bDcwJAfxW
SMRlZoEMEaVfNxE3osEQM+nEiwJzz8ZD4EG0s/37BgBLfMhkpEfbWtur2U8Dm43lvHy+TZIWJLOR
iZuoJnY8NNM7nTNz8rlhiULy/202i1kHQUZsMpWvdXAupLmvcUenp2T1fAk0kjTflvf+0mFpe+5R
RD8vmZbn3P4ABB99ulmG+gz//QlphjQIQfXCCsbxMhl0T8g950psSLpZwsfqETVDhx2OWwgXP1Tg
YXD5OgY+MKz52KEqd/HPhC7EXbYJuaAJuF1n0dQwa57JzXEU07Lsu2rusJcGZrPID+HiKSgGRyom
FkZAvbkVB9MWHnacdUTppwmD1kYRT5EmKcVrwx9yHbqt1cmR/EQcZddrOx+i+oxX/PSWIbXg5k2C
MeFeh9sOQ06Tj+F2Z4bfkg0XgXgNDX5O29IF7Z3eNCxFlOMyOlDO67DgZrN1D/k3WV4jfZ7BV6tJ
pEccH2QMXBQB6LYVvHIf3iXIQ3dZ2UcoF12ZT/uyx4hhaKaIvWcBLB+sq+Mhp1kEEx80zo6KloG8
U+Anx8bOlV9sMN1mPIOS1PvYpvm1sbu/hOJxgDzmVzd3F5ip+fphT+2Yn/nF/5FSoSJ4i/n6WeHu
DCvRnImf3esJNea/W2tPSx45S0zsuULqRSvFJS6lSCcQ87RlOjKlQigsbCAgRGbN5A8BskjVNG9M
pKPUz4RkYLoB/jUqszP5nd+KPY1vNDZwY2IzoG/41ZicVKy4mU2yV5BXv5ii1WAl+1JEtcWWonuS
11FEzQK/RokgTCAg0dWQIGIK0ieMscMh33xBHKSHnwQO3CF94XiVVW4sLPYxyFatNrtFimZ5I1hS
nwjM2gRpNh5YTxmUuRz0HKC0xArcBkk5q8necNZ1mUOmAOevWUw68rImvyZFEcHVgNVQVKISKvD5
+SdDhJ547h3VwDR6weeWufZwiR0YQE56we4ZYDiAwhqbnd910TZNgedVbJAX8oPK2YaOeFqOpyuS
1Yr/UPvkZjf03NbQELiA8RVpHIkTtM/IrjSb+1sKVvMH26OJ8s/4FemFKPgIUGEwKjIDlB7SrQ7Z
zNwLvIoNYsrHOs+6ZkawvRMioRmVtpnDEpsLVVvfE+bT39u+/6EqB0uWG62oin8ASY9zXFwrRXNI
oHSRLpxYj8V5uB5OcPZU8oVntAr/q40/LsjZcuMDHpkuXq5FocDOdOsyQRj0hR+fhnIorylRthhi
L4GYbb4r9c04rfZA9Q8JF2GM97aQHO93Az+usy7+g/KAJQddnWMPeTv+PRqlirGU5M62YhVQbS/T
ips24horPqyYCYfmzB02PE7/Qtwf2CZIzgWvmHW8qbeZOK9oX2Zkm0mzQLmSmescu7f1wemc3FBa
1IzW73ivR2Z7FcgvwdMBCz9zoqiMNxv6kF0awg1Nb7R9a/OmbDFuxUmD7Xg84UZnxUOnJLqakbcR
jZ8vNw8WFqyQXHrj4r1R1Cm482nGFiVqsTLdkOIjv8bAItY0azvhPtom0i2V59TKSOeR46Ohfm1Q
4sxZlhhHkq1B0nw8LdeA+62eEt4J8DkavlMzzQMQlcG5U6m5aPVcWtuBmWWRb0ntOOd2E8GNIJ07
ILlRBKiQJVGnDJCNOZWuJlXvkYCmvepgw3XStipy4fRsVwhlq5TGsdezD2Ny7/Ibtet7oW0de1Pz
29SO+ZN1Qe86MdGct73ZqF5Hetrg/NvQio/JBGxqd3u2wuYbK5EGDqZ5/ihldFfLH7GCq4hjxn8j
P+eYahKRB6s/fqvIXZgykgV+byOw2AEtl1QIblF5WRPo+w0TAlQsdPXqGqWkYmrvVCkEQ+WiG9CG
m+MTmle7/NZS5YBN6xZeObZ822adH8iMbJZqPHRPmPPWur2K/mNf8wD4xzZkelt44fPsz+6oRinv
81DwmVKEyVNZ2Qbofx8183jxdQulZcYWvf0ng4nBlumNP0UoPQkpbXR0QJUPQhnIHXqZTaX2MWal
LQ8rr8vrg0DtVvBi93T0PKP440MVCv0oavETBT6c84ec7mfmknncQ2IrY783WNcRs4D+9ccNHxlH
PhOEOHOJIarDiezmXX8wwCrlvtQ4D8aIG6PAdX4jRl9YbgD6V2bhiSWPLwTWUokh3NyblhQzq+m0
QBsaR0FNB0tRbn5DbY3ONVawC1V1nq2+M37n5ySPsasvDoLm7EtAvoDBOdAt9MqTxQO9goEv9pzS
t2Yml0g5PBF/DSTrD0RK0R6vT67QBADAT4vyFZ/eunRc34ypn9k6ru6Lazi43Ld7hVm23jaEWoQJ
P1G4AG7LE4ETZZW2OLQFU8evdYGyKzJjbpFtpVlVvt7tAn7aHBRENQQlcomnPyI8XVH/CpGtQTzB
M1gyC+/b48SLpdrU1MhTxGKBRm64JSMvJtoCIcmABEGjhi3Y+jy0jX7OlKNH3q38FwKU35NzJuak
oSqF/hnmUsF9uqYkjRVuOhRX0nwwfeQrWf8Z8MZQ9z1EJTUYCAtcM4Fy/NjXb4FW+0GbPBl+s+oK
klAyFeTIQlL0XIhGymYnFgOqmavOdIqhwdA/601PJyQXq57K4inEqF/IB91vslZJtpg8hGEnRt9F
RxjoSE9gsxSjO4NqQAdgf05VpghaOCdylebrn6+I0TNvZN6HyZyKKT3LLI907qFX/z87w05U5tus
sjb83K6M4mBswAYtBNsf2xguFV3rSX1M+VL6Sh6VfsGM7oYKWkg4RDyoNVKp+4sNu0aeKrSlJOoS
wpUN/dg+VTb4u/LRWtv96I2JZ7ArQCLSD1neyxjmgzTGviZAeSJ+nhCnsNxr7YX8oHiDpeTtoPhp
s5RdMNQtILvajR16wNgKbUrRJV4mYSGHBfHtaZA6XgOId2INfY/5h6LulsgUAopGjX3F/8LuDuSC
6QB1pA6rjrOms2LmyqbROcf1OenrfnLaP7vb8cCPFw8up06WPcqVY1uhsu88BTuQvxWe0iT2TOF4
WHroez56Vdt8Qko8pKJof2YUt1h4BYMbzBHed5txHInS53hGU4+uY0NUhf0JAnwSFWazQrQEfhip
9Us7KulMKFgzPjF1uq5vqkRy4U0FyqQM4dDxQhuE1op8KTL5LM7L/tDlzVA2Qo8OEZhMIww21FGX
g9VykWWefmSdXTqNtalHx7CpLuEgPZm6FNWH3cdE/bDOfeEagmoePknybbo0ZZRX/EZUOylcbcKT
ipIm1gcpT/E7PIMd0JoPEOcUVCrEuvJFaKlzK2IJM5LpzWmCqmYJcYQ+9RqemlQWFOENmed59IdZ
e1xHd6N/ZuI1NK/25qVe9YPeVll//MDgfrCTdKdbdFxA4nqUcEsWsSr33SlBv0jiKCvMujbfPGmI
w+fKUdJlY39TQ4o4quN8a15MFkAG8Zf3BraIA8+M86p37om92HdqY85mTM+ZCE18TMIwFzs9twWc
vtdJL/CdUEItXpgdR+ZV0hzw+neYT8S9UH8anPpeW3aQJyIYkxeC2gtYOxGavmEz1AnDKM/sEIO2
Sdd7CGVeppmXAf7HL2WLI5BIu26G0IylBOGyP8RFNN5qV35XxzU/w4pKoniuE6ff9re1rKZlpvkR
F0t95+0ohdmOZ3ztucsOKSCYDexTCUvuWWudBXLAxeAvEOc1Xwlptc9w6xNlL2LgJPx8QFTnaN5l
9j1IIZOmJv+MdNh3ax46hfyJn2qR42xGhBt/KI7v6Sc6TOAn2Gzt50zkByci94R+Cva908U+DAp9
fZDWtuU9I9/R+Kbj/Gk+KZ8G5kl+Li6tO9iJde4X/hj5ybzFYKLReQkuX8W0BYkyU4+CI3jhx/Bz
mM6FIwyHwcsezoU+d7w7Gin5FedxDUT/pLsnXsLAOK95Va7dng/JxRK/mQ7rMEaHJnJeXt/nEqvJ
jerqXz50BwwKFGAU2Q8b7DoqcJc6h98+nhSAzSrtQFZq5G0L/uxuAuJg9dEWFz58HVGCNJ1r+yNM
2zAlMNj/Ay8OHVQr2AGkavlmbPWYkvaeW5bP7tM0i62nl0J8RrGLZbougUHxjJrzBssmmGBeyDf1
oTj3CVf0vDdgMeCm2/xSD5RALNYKcyY00MO4YUDDG1D5PfE+3/f8Itt1mlOUSgw/CYyUu2bjjZwQ
+3YWxFMBvAaAMWs8GJYd0cPsmpMHKkPErlefpNaEkwk+XCQeTZ7W180060cQ7WgWT5SAXhoiVYJB
5d/fpFL8SE64m/slEGJ0d+pPasjqC5b5QDpOLLG8IJk7OwgvfE/Xft1QtPKpsUMWPffKR/ImQ/n1
Wmd3ks7OFIq+FiGV6b1wJYMsD7GG2EBGUMSuQriVfb0JaP8Bd6pKmfDbFHIu4QgZ9uZsHXPCMRJU
dIl9rE3R32pVw9QBFNy5IrGjvttyE+lWS/wICNq2Ihjxl7DJqOFf5KugJZM+mL/lUN5rXckFVFyU
eBnjEB7pmazW+LmaDVKhH5ztDZPtEB/Qn3XJAcdqVsU7kNfXGKOqL93CzavMX1gCwVE3vebh9Bpv
8U5dgYTZ8uG6my11t7uQsJ/vdZAvyqi9FVeIXfaFO6t+kyp+IY/wCX1cAIEZiEKo53VkZzZZA5es
kUoDJdNeMx5R2sPo285W4npRpr1hhxXum7Kxrz4XhCYT09xIMfAQauzrnAzWK28esVQkQYuqGdO4
KxjSV2dW5icV9de5sKS7EGRGXJc/YdyyG4xOzi27WVbXl/ziiELt1774Vy2WQyMYtisn5OP01aK2
41twDj+8hEpBXuxkUR4AzNgkOYTuO0VG4+IOvS88nh720JKZqeyXAjWBfHK/0BFtu1PPGaQh9xl5
12tPW36gNl4Jp5bKZCSaXsJYc/0nqasWlp4BeQ3TXhcXi+mKwY2LNtw7NBjYBD/wyU5uMXCRPknz
aKVJ8R8/ghVbCb7sw1krSql55pRHRpWbUgb6U5jRwODqdfSeUe/PPg+72tU3MZE8Z3mwrKHwvQu1
8pNcHciQYn3xD/Xtk7B6FNo3V4zLYhWQIwbusKQytWDFFU3jwhDZBrgoYzzoCFPHbH5runBL4FRm
UNTctyRq6hLWdcN/4PC+7+FhbLYiGwNuq8RKkfaf78Iy5JBV+Kvxblo9B3dn/5rhMO0zpVcHlXEP
yOgVc59VPxsLmQhZ1LZ/+lB3aUrNxHrkd4TbBXNVG7QxxCWd4gZMSqlKybdB6IhaxqIDQXXQg37A
bLvztsZHs9vdDkby5ZpY49N3Io2D0JVjErP9QvTtoYs2Gd7CekiLIyFFYKkLMjHBoK6u9g3gw/Up
qWfennPnL+ueOoKMjrikRYYhdnMasyGtwQeUqrpV1EU7DQIxVlUzVBAU0KYBDqMhbXkQn69dEKsL
wTJSloSH2hINy4qs2nQ+eMMGbUybbmfoTAroYx2R24f8elhADRLvQQK+C8pjyNsoeNedampNXWxr
ygs4yZlnsyGSHkAb8yY00pP/UogFVhuF9FfWue12WYbv2qsP4sa7OZsQuA5iX3+DAks3o73HiYN2
eQJIIzLSA+gDhxgxvBoV8MlbPUVOwWtEUAgb8WFBBwb+EQvYSqjo/TqhKUlgkEKk9BE8zrljhZ2W
ybSVFMfGqxPbyMyhvfeB09GwpjfFmaCfudJzyqfPRPDkJC4/Ess2DA9GwsnXn7p9/4av9/r05MmX
8m6VN5Pzs5UDO1Lci0hKqnnXjmY/C7mIfHYhYhr4kCLQOnSFtKxnopSEHrobDyzlfqgm8Sxak9NM
Hs8NqV/ko3CvWonzMxdiNZaVaaif6eIwDqO/C5MyI2wa9uAp2IVafYe6JHCoh0QmQdB/MUxIaZKg
2xr0F7qsmz+z8ZpEQzwY5nsJWK8XPmpt1NawHc9iMi7qaFyBuXf/t8LwS06tGDbYqMQ+hhONNSSo
r9FyeSfoToWrGfwtZv2i0EvTJ7mIAMmuyCKCv+6DTvZMrTyOj8uyhIOLIT8hAgHQ0oFvISOKyCNx
gd1aShr2PBlhLJ7iPG8a22LYmhcB6woLeVjqfWYvQf1jfI/14PQr5YsvBUyhXkbkWJ+bvSrts9Xq
xbcm8UHbzfALuFOI256PkM1GBvONmFswDVVzkQXSLwwStszFPukZS/yZleVR4xwhayu/28jyRSXT
rPq1ewyWyFdpuCHZXSaWcyjAAW7kKyyJc3v3DqBFf6/SF1EBE6T2sO0nogNH+wETi3YUyxYP4Dc7
iLYdYakwojciMwgWOqb2myD1GUP5jlNtl3dGdS0RGsYjDm3eTEHEc6fMsaUMMRj2ZPcjYl69Y7mI
1QkgsvwpazEwExv6ZG6KTgYNvOry5oqjkeK7XuYsrpFIWQ2u+FMbmY8Pf3e3Gf7ftzK/oR9s2Xn8
2dmkoYBhrkUByW6GyaElCak8QR1ehVpkxXq2vDJrRerWQ+masZPzf97EriFxrGoyjcNYqhGBzwVv
mhdeUd2MhIm0WwPJHYcyKdwyNCQ9RA0zMmehc2wtP2vzGaUwnMmaM24pSnuiIoVttNT6FmKXZHx4
eJNIV4/1wpga4PDAac2bVENZU7BIy/fwzf/5lPk6913al70WOK6jSLg/4jPQzJZPhGD1+tDA5dGi
Pa+U5Lg3UIPJdgV43L+iKceqOkDRIzLJD8qOm6RsX9IC9DYpkmy05lOVQ8Bxjf+bweP8flvGfLmP
i73oXsRK0yGz6RU9lV7E0vuq8AMfCqyQmqDpEXlDt3nrfXQW0kpaGwf3fnPjkvkNyiJPLgHem89M
haOU3Izlp8DJcug3Y5gkZJXbHCaqNE8V/cSSdzky8l2KfagRRrOah0t5mLmke7Bx+LSs3W4VEVbM
ASAVzoRAnETzjiXR/Ip46mjsgWgxu7GQZ5051vbK8khPyCQHRdqzkyHVn7Ujxfn6ilayprh63aP4
9RhZoVpA5YZE+bhbgJW5MNi6uqIEflHEjBXBGfXtD0/fFo/pu5luwQUopZz+r7Rl6rYamfBY735S
/D6SS2GTK7iXWa8V1Jw83na62+ztL0tDFSEMH1QxIg/nkvKyUgUKGp4yqTmNT1pdbZKxlNCIvxA5
WHm2nH3dlme1dtJxrSKaGtLoCIGy7ZzsFJO611g6pVAfaAmhKt0Pmc5Pb8m96KxdL9oy090fqAoS
ci5FFt+jey/MaCvH3eug2DpFwT3UUaYMR7dRBCeozy68DgVMfm+dELF5tPKyW7o7rPJs+ComYHdi
Ozvta0rvWRWZAQakh8e0xwTAY0GiSKpu26ntoXf56g1OF0yPoD99hT80hSmcWR1hARaJ0OfaEdPB
z0Ncmig79t7xcURQ9db1ZPEIk4vf+hhxksYS0thBf0hUl6KvbiXIgP//m+5RGQgXO4zDnmjlqm9/
zQWvBe5EwPrF0uXGN4o/bPZ9Z5V+qLf5FVFiPxX3rx8BBQPTTKpmz1tyXWgi3EuUDJnfmux6QPyw
CnKTQ9zfhbUFikyIWI9h925YuXNakGfFDiLnWim0X8kd+DNEIRpwSuQuwRLK6brMpDfr6X28GzF3
0zP/ctvjPQ2f47tkjK+K81fdLJWq93VTCXtPkOW4+Vnnho++3ebQeLkMBLmCpp4jqTDWAjyJruW0
oeEuwIniIeZy1xXo6lj8+h6Z3vadmb2A7I5Fk6MrGCqwNkkSczpQJ/0da7ysY5+yNlW9eaV47y/n
bFA/muKu+nyLB9JegSF9wl3hdoVlZT5yKJb/QBS6ig31iKKLpnq9FXym04APQ4vfVm5B8NykO2av
4MdMLDZ5wzCK4WHWi3R7iO1Mn8KzdSdFPUUh9iKDw9z8UJN4lG5PJvUJWN7blj6ZxbOqkTjEFxeW
Sgo34bdjK26ESIpPqDv8PmUEaO57wOBcJGtZNrb5J/apKi0Ua3C9AKpTv9k2f9jbjQDit465faQa
3Y5WpDm3GFfEm66AxX3yTcES//PAVuDjUe4uwI0Lnykp+BEEjS18og/teZdAQNkzKwIxcWvypTtl
72VIjXW42nOW2nSDF7vP3sDFVc2jflrv+CLOKwwWkf+VjeEOw/6D4Hc/L+uGE/M9JfZlQfaPdl2j
Q10oPE7drQgtd8hW8ly/A1TKEh491+EW/KeQBOzOpGXg76LurkxBgmetpIdL9nGzd2RgwGUuX1DV
5p5F1jppYU98nZwM0wx0mThS2VbUyrUNL+1UUK941qmaJ57aDz5pE89cFRf4b6u0NlG5eYo+7P4+
DREn7s0AU14X7BbMg1zRWEFw1h6c1wIeqid3mY8CkIht/Wum7+pWOHkMRe1EAobS1ByVdxr7ypnA
e9zM2odlHVQDElR52Os4lFuTlN9uR3bJtVl9Z97LaAUdY0M82zR1gm11Ymz66fUauvFn51x9ZTjd
V/+qO/qc51+fPxzdhb+AtD2Nn2igKwHdj+RAfNEFAh0/iSIEFyZDTORYsOgvgvq1Qk64oL399OgL
Uy5HQQyHNmkDoRbHr2CXRHQjBEHZ7TBBb3MnsgqjzdKnwwOLaf1/b4PgJMtPQzis6RIgG70Ciycj
qWTDYtC/DCfWBCPTwL6WrMijtlw0anRP8/plK3Ep4sFLp/Z9lOO/1IbqfpI4CKt3o0F/tIfU+nwI
ynre4AVYYqO8pT+5XUe3GDYGPyASeCTYuZPjoTxA8nCJGhwQzCqCTeA8nmRFP8VgmPuX3RTxVThM
WOVrf54o9mNPU3cHgmu2IzQARaA5aNZL02b9hQS+QBtS1Q7LKDKqDm3px2TMPWlDexUCpyevN7nn
u/iK4SN5VBD9JE9N2v6lS+SFZpVD6bb+zOk8P1JQOa1J3PJOZWg/ypZtXoNG2OpcOZ7vwhGMILrd
YEyr/F6s6GJIOcyVeec/rpxkcNU+YuxK0B4XFwinGYq0HNXrYDQCTNFYM1vSW8zt+Ka7ly5WeBmZ
tj0y6ADW2Mr6rYYIWqXfX4gGsDxYWzDJnwSVRVbOviniYYL41tL9iYEZmV9huL5AZgmowLhc1A1u
JJ8w2YynVuG1mvpXGK09xGnTIp7OAkCM5bH5KDgbn0KZgLlR4b3UdTlyWXJngGhYsBwvPWNztp3F
vCwBUKo6ZpV3aydNFD1WK4rVYnPMAopXi/PlQM1Zj2CJrNFLcpK+ZniFFD1FS7sGwg3SR+X23ulH
SZAZpPr9Z7ahQYIt26qF8QUA2+YL3mQE8sCgKBg45lNAn3oCV5pcEkcVw+yDWmKMAuVzjP1g/aaM
4w04Kv75AVT7QXxIMRxVKtbMj657nKXeOjeZAXZQhKwDF6r/7lgy5Lrl4PX5Pobdx6go2p0/5N0P
NG/bpwH4CYFS/S79qVv96Qs6SRchj+yx1BjbJGZTwxXMC+XbthuEUjuKOAYfJ6RShc8jJBitJq/5
KYL5ojTJPjsSHlRR9jV0tw6oAF6IYX198ap3GBsZelFSGxSiU8rpWY/ltCH5+tsfGvnOBydIwTWr
vbg/LiaFiKA+PYrmKdB6n4Z+pl/jLpQ25z9aimZTZhlvRALZunBI3P/APmIswXZToIwNtl2lDlXf
D6gj2LQB8AjL3bis1I00ieumpMkudtvzujW76crxJNVLPwAYg6nrYwkC66Wx03LMP22yeYVgLqRi
CvpfgKzqi2UdB66ZlsHbbE8nOFlQVuJmP4cJZXCzO/fnUWsjwkpzEf90soo4K9MDJviTsKGpb7l+
iAGzgTfwotFqFkepmJuM1nykO7/sqcUEBdIuZoqfIrbirzcxn5X/tWXcq1fEtokNaMzqc7Hx4oKV
UWukq3q8GLlELjR3L1eASRVILzpCY6QHN4RH/yVYtp1XHRKZE80Aye0M02l7Pi6iGtg/+x1dyxSY
Yp3VjXwdZJ18IVBIUmrBLi1XlOWqnRcmZtbBF/G6IStn72WzXnPtgoai/HjM98U9R5nmC9O5d8z4
/yyAtDFXFmKOVCA10YCccfFfB+oXJPqk7SlmTido69TNwp8//ESiepR5v46czfFwcfrSRRJ1BaEq
jXpzrySbGgTGILLlq3+NbBE1b87iYjwjImBsQ1W6zqKjS4hev6ZKlF1yom3G61DttFB81+/qH5hY
mFdSlKl/vup5eI/lClVGHFY/JO6UwXgS6Zm6aA9eq2/2RM4vJTUxGbqrg1+xiHomE8PU82Zqwnet
fgRB/mp1AO2i7hGq8lAIukf8k1ZC+usk83bGMWsMFtDssGZDxWhug0bkeDw01PcURZKksWxfhdjy
hw1Jq/oFkMa1Satb/gGQQ9HxU7JyA603x78naKjDmBbHF/71/zP9Lo0pj1CDTxI8R4D+L10KUTS4
YyGqxDkA4Db+/ftvWWl+eRjT4GhujIjLTUMWfloINTUbALz2sfhCxG6miVoMqtXsDNoD5UtK5B6w
JqoUce3vJmu3q5ci2/7O1YETYeArtjTpWgWk4MOKL4nci0dySAf6xSHBmCPMmZojSQfFrBy2y5ci
OSgqcCXd9lmj0XaWx90ZwPiBJdVUOkO1jyQEv/dYT2lrBBSMrE12/joeRhd6nALEa7eFmRv84dbJ
g/jbNVOoS8mHP/+YlkKnTIg7hQfYy42zEOF32Bw8VrrrzcCdeaWiStA0JrvYm98mGm8FR5aN5Wo8
g4y3PfpZq/41tsNFoilwY4b9NIK+VcPuUyRjAw+yVhNLYif/u0KCRhKhPFUbujlUqpgIaY9iCPVH
6N+SaowIZgw5L3E/jaeX/U9MmBj2l5o2CsKBoE0sDmgyREzz0H9equOr0heN2dH+0xX23b+bWKtc
0fW2gPCPG5zrmgDnA7zf3+22Q+GydNaS3ThkHftLA0fcHApV955XoycDfYzNDeK9HIh6pMlYWUwb
ULcXHqkJFe67ze8PxhNLgmqapxiFYYqdFxuSMsHiQbUQ3BSqlyGmE4ix0kfKmbU1KS8cMa7nTgb9
3i6XODoannkAInwdcnHhDVglobpXBv78rBXixhKax7EZKokhXMI+nn2jLaqotu2uX2LouTVIAiGc
dmLOzUF1VFqk/X135bF1woUNyA5TXFoqRJWf2IRhyXELE0c9Gu99aVe9C0LOLpEEP1dvePCyBFtb
dCxILBABcLalruwdA+QHH1HkD1WrYVJHmFBNI6nwtsoUFbxNH+KMNVzOacuE4nVCYNkeLo5IkDBw
raUYN5zXj3qfWtBnOBFy8mupYTRWo5cKjnYrDKYmEy5LoG1fwi1isqRV8RC8T7+5ZjiJzBv5vSO4
bxqW66N9KRGOSW+apY58AieQHImBAJ7/L4FJNBbf50kDj16y47nKEIvoJiFQIvMkmvzoa2BsXwcE
jvNTX1nqkQhy+HWn8pJ1+BIZsKa2JxYagLpxOWwd2eH5PC7OSwVv9ahsDHRzJr61WwRP37Ifq8me
mYqq+9gNLyEurC9VTBskCSIJ+BTxzuK80PUMCJWQRT5TYw6FeqJuAIMx3TkJJWQYpiN2Bk7wqgCw
sGwPK9em+CQRPRgQ6K6STHjyBCL965tZ70FlYti2U4MQWoWxQnkCIpKMSZPjwbx8MjVzB9ut+cre
BCslI7KTh+OVP09T/0RcFaiJr28My4rf1/QDtTO2q9+WtbTN6O6dcMKn+czchk1tmQ/6w75Vg+nW
u2gwKFX0B21Z+Eb/4XYXTKk4cg+H2zXsnF4oYeg/wLL/L8pCg655tuC4e8K6OFWU7I4mQbP7Vw6j
drkyGg+YQn46j2+zIPkQwamlZBsWdmri6tmOOe78Dck8cdPbw1tc+ZSNh/NPqxVi6MJB/9/Z2SgO
ufqldbpTnHRxIyb1inWXmmVx00oE5MaDJBAzRObBUuu3JLs5eZT7GbSRcK7wQNy6CH6DLa38LaN4
a6+fFM/3uIpznFoX6vKY4olwHq0NAehyv9Uw3HANxdXoJZLWI1fq1Br7ate3iZv3JJ1gQCbfFpTo
DgNVz2aefn678qg19HfD7+go0AwjDoWycjtTFBpLTtmfB+UCGhiFiGcxBqNtQrctm/o14hP3S+6+
3680vOAxPjsCHnm8IOAx7lK3NDVp1S73n6ghDAV7RUSxYlKLEPht4QB0Ar44adTZj/OnYByHo553
Iz58afERGgny9GUI+sVKxgrDsGNWFqAC8rA6TR0VjvsWZKdmSjFvLne9Keqi9LpiFbgIHSStK+8c
zg7rFnMkXB66VnatvsVx2vDBxwVvTR/1QOnoKY7KZ3lFY6iA53gWJ9mkx+08TzWh9Umke6Pyv1Pw
kGGbevMiI9IhGIC/UusdlUd6SzdS9NmHYA90RHW5g7EgDXgH1M4SYUzHSrW3/sdtqiNO9Gq0+gY3
MxfgOIb/64fPxnuObV86tbWKZxjxKjpJwJdWp4mLIfytKTTS+TNG8tBYNckBr8dUELXB/q+J5fgC
BMbjd0OKRJ0lspAU9VtWMAusESEwQJ6t9eiTKRE8+gZ+eaz2EqIAr0Bw77d1eR1w6Voy6DmzYKtx
N5lIhR83W5eC7NHl51Aj7SMNi/Zm6HQCNesuUoznW/ZR6zm/0kAmlZMA9JGBsttOQmsk0dio35da
PoAeNvCNxwpnnmSOx+AiI8TtqsO89KAdUFwos3bwzx4ORSzSxYp+BfX5FcA2u5O1PjjUYGUiGvOi
Pq80meaHhPONHUs9o/NGWeQHk14Cg3OtF9vrMmPSYnR5ijCZJp+hBhFIhuW9++ruLR4ToFipSoY+
xNTkMlayPbI7L3JtOmBNieWxKZ1vfGXNhAfHIrpqorSanMfHEhCwGyvmhaTM1D1/rRgheT1g+xh1
QyWkft6g496QdYBwg88rM7yQRVFDHzBU2nb6P+XSjtAjaQ4GvBYFl9U45Pnn4teJGY2/wIwhW5nV
AMsNIriYDb13mHOIJE1/cvQdg0MgRh3pspe0dSNxz1wHrVDWQmuifJl3IUE/HZyj1Ddzjt3B9X22
WqTz5C+vSiCRIpWVMLCdJHl8zOHmIoYejULfQMM80tTsgnJjMvp84s4Bw+UxCqx/CMTyGVwDCEaC
bOAq84pRdQl4mtM5syDmP6miOYwuSCft0i59igf4JqXsQJpio+qFrOc2Tbc/DxJ5jRiUVg0qeoyi
hTMSDO6bh7vVe7ntFVr6ce5s1Tb5GTsFq6yVwHgwLW+3FVrFSJWCLw3CLcGQkyNTFf/79q736eyQ
M3v9vn9pDt6p+KEY1xpS+6hSpVo1iQ74FMDqD3sc05o9rh8thHY96WBIYe9Z1OrvgDZhJUTkGumm
2vsiYmTFGhl7UwS1NXXJyjSsJeJTRAgNv5OL9DOBH0jeKiS0PivpjtSJUrmkh4ojaBZUm1G38OjP
+qDeAOzesJafFPPk8QhHjuDlfVWUEyEifPUDXbnj8TcW+NkBErkslF9bV7b7DuLxoF3VKsES4PUO
VsmhU4c6s98Qs2EI57tOC7l4b7JpSjERcOyeW7b5S3gARMwPdDIe+/kG5VG+PFqqV2TR9zVE+j3y
tpy1YGOD51xHsCi5AOmQh0+yLN10U1ocEHYDXvC4hi7j1jlbX0w88+eOjExamwChp6IQ/IJKvtcS
iEPQ85zsrR3yBQsTarCj+zlVY2EEWqC3+JPSkN54P9pyQ0gCohC7HMrNUt5eDbErd1oZFqZru9Bj
Dt7wxI6kah/ZsInT67H1XFexfDDcgcnbZrhayfMrG1hh8lWce5TNnnw7lu3T/ieRSPxyTM5uUlMI
Wsj7rXOHxdQyWS0BPSV8lSla66lfSepryfYFkA4bXKJryYZ1eerCd0jPd6HxJ5jSCmrve24I+qQ1
VAYmWBXao1UZZp5dKKZ8fcZB5QAydnRGlkr9M3qtrrtOdaBqC7IlYAZWi5//aPdJ59ZD+PM1nyNm
ilhf1EU5DFVqlPFR0bGyXZvYnA+2rUyMBgbePbGq3Cu3CvSsopZwQ49YJfHgCZWlnfgPZvR+NFHT
D6/SvebnjgteVlynghRWdgIUAHtk8txRznjpXGZiiSbS5fRAPigRHrIYixi0ru76VZzxL9ALIdf9
rCxQVBLwkIb+5ML256g8dTCYmjQ/f+3qI8fui5TVwCtNb9rswH0OD2WTkLBYbKosZ02VB5X43oR9
xKWX57y2VMo01vc/Z6Vf+tzDackMl/4AZALefqDSNFIg5sRzgQ7PA3dbXS3QfexSmgr96ygCa9eY
FzrUUXflL8t8UDQJDSoQSlvN10nT16CgWpQ7u3q7fCNSJDak/8o3Sl/6EkuTvWicfz7dUpJPgxPc
/nk8+m0hwdU6wq5iPsSjuZbpz6Pc4MxttiB99CJ+3AvNQW8eVHS/uz4GJaUDha+LDsFUoRqIiS3J
RB5w3MPIK4GhJpq/mWzXSsG9FQ53pO9Nddfcx0rM3aXyQ1CvkEQ0XIDjK8E0ACzN9DpB+zGs8KgH
cJn4cBu9KhwwMDscMSZxoC0xkGiVMLd0jqukLfSTJhami2mKR5RPtjfWMQJeTVxRxd9NikkR0bVk
/IGu/fW0AEIi1tCmiASaxezgaerEnI0yh+LvIQJKcBRuJkInVYWpwsCzyUnS4dLQ95bxIiwMttEF
81r0WH2KgkwuXhP3M4AHgN8b6H4kBnB3U9YH6UAEV/wE9vzZk/BLp5eEm6BZ2SgDmHGeNA77ErBm
f65eOBoN8rUFNte1xJfHAV2tJB19boJMAr6HZpmV4+VwVeIzb2g8F+VyKOIZCPQszq5qj4iVf1B/
MWnO++3BpOh9U+N9ql41MgnrbfWUfbYBuhZHYVv+sWwbxU5F0g2NGUjV8Etncch9XeF8bq6GYee5
u4lltX+HMQyYBJsRvudNE0BKKl7YFa3NU2AxDn6AQsSwc9IaOzhZYc4TQsFP2PUnxZkJyZ+A3grY
rcktxrIG2oCIkJ1g62hQmIYcrw0LxgM2DUUgsEFB6BlRVaitQX9HfKD2APkcPYL7gJnPrEZJ0L3/
GBVLyvnKLJpqxoJwI4uN0naLiyotjVAt7MarlhHpESmnqp6VdAaBVO3I/Rm6B0LyvdA8OIauB3Qe
0tZTbja67mdRVs1urWf8nP0dOZOAStDUiKg/9LJtUllnmbgBYJ29C17SGzQz8tZ/mo81m4gqvqIi
TRPQ/Vl3t1Cm36iF2lk6qMM4sxQZM4iGhpP/GpaPBqxTSQ5mTdyBEw8GG5BjSrTbhnxK/hjvwCdu
kpDS/pOU26J1nk5jY7WQN/OtS17VJ/67tdmdw6Y/gEpgyN1uygbxsQYV2O9/UNNjEaiytRYn18UA
y9lYPZn2X6/GUw3QpctR2DnS2dxxgGOmH8OTdAnKPw+MtH257jNVmUYj5e6/vC2l6cf0oS88HdQu
ugwwTWTgvwWl1uTdnvlUCDaxaGhVxXSQ/UXcmGRMSoDilef1lCny4KSOO6NT8Ib+DOUQLPykUg5x
RHVJgahcl3PDmnKVoYfh7K2iXlkLywZOkWmWuDWJjJFY6JXzVWGPzZXPBIuEZvO/qOyIDPl4GdMI
TC0mNEz/f78aKNIrYds7TtE9fuCjNkyZpql/HKcmRb3ApBUo9yZ5J6fP2+wI6YVUfyPPRQAjMUcK
SzSJolQC/EgwMGR5VtpuwK0C+77xGJpQMJqGjftiW1mrjCQS+WEGtrN0jVqDFRAf9jbJ/wR0KS/W
d2aThUAgmYPcXRxmsRl0O5bLbKE4/KQl6GAw2hdGMby7a41OR0/uzqvwpyqOQschSmM46in4eqDc
AQ+istUoRNeXaa65O+f1ebC9U+1seRujX77GaaIbvu9LnfO6SBeXVT3LIABsAgDpNSixgiKS/t6a
FtJeajOucCvSZ3Hc1+Deapd4GxAbm77phG3wZccDxTI+MtrQCLgMgL+QFrsbqgST/8/q1vtzsn8O
9yBglK6ND08sFoCa3cPyycQcdcVJTs231pGIzpTBZvpc6L2pIoG0IPHbenFrQ6k3onrgbmT2Y76M
EToAnogVJig7hgzN9FM5BOlQY5IrNL6nYGEwlPk+LVBfPZl5J7eFEEJGZlEvtA/FAA6cML0fDf0w
sQ6bYFORSxQ4BVlbrQd16P9cc6a/5OEt3FPDWqJrFUwoxiaW/djgOPA9Kc1NkkNAySTp0hrJdZDc
+jN9KBjBeO5XW9c4iq/ORfP1xZHv7QBS30ZoTJEzLhufLG+sok36/0B9htsMUHk4F7Z5U+ZTTQod
a1UPR6Wxd+AKrtScYNrgnByyNdyhDFoXQtqwv4B6ryTVC4sNJsPA9DbrQXIbjzsI8zPPnefrSLyX
9SaMKlTOZdeR9JK/W4IcOQxJKFVKjTDL0zGW/jAI2Je3ytlDvLEXxiD47dqLdQhNkaSlhacuvqXI
3M0dHUascuHuJnbZqEWn/ciYi6pmjNee24HKWR3E2+XP52H0b6geWvrMlDHX1eEm1YBVeCZ+v1yP
8Hys32YwG1gd96ShLnWFASV51j+0BGUI57HZtLzTFd22H3NZ20fTfy6ofEV8fzGqxVjcSjHnzj/L
w78rhfLH3J7y+SEr0m8sP0oS/rGxecUQ4TbIoj47Vszhf5gAzsQ2Jotmdvy4BYGWDpCgjZjaZTf7
IXUddEeEhfzKtMEJJxMgM5d6ZLDv4fI7K6H/ZlaAJsAakBiUPh1AuJdMH04Q3pFp8UskCTNMhB9B
OGg2upIguSvW6kDj5JAMCDjUwQ85w4Xw/SGQFioUBtD2HP5IYrRCMn725VAGKxAD+BkgABXOKkJS
G48dFgAnZSHJhegSm8LUq96RfJ/C2wWw46/mrUDewXkbnv5SB+QNHlJIvD0+KNPKkBTgwig41DN4
ryxF1U4aQs2toUXwuwHix/hyl/kKSxYkW1AB335LQw1KfFpkKCuSRQfjk7HePiDDL6oWveaonHf/
6grRsI4ejWLMxbiICOVV1MuErFcDf9ltj1p34hGOpuQ3V+0/O52TOC9I1U42RDNWTn/Psik+e/3n
9SOB8HSxjy05zDKYbv3OX9dfwqc0O3nSNSDyvd/I3/tObkyFeGuI3WgL47o2XbSGn959EtgvtNai
IT+aHRzKoHP9fDEgbRSPmtCOr8gqym1+P7akxPfO6Ec1/2XMDVSvedTZAow+B1qtqxcPN0gpLfKk
8vAokYSdr/pFW0amLYSWfGP/ArHMQymmC2nmXw4otlQgmbO227H71qPbLv8EiQPcFp1CEIkdnOMD
MK8hEiQ8QhHCYiW8Rrpgf4k/68MSfCZNVubBBM4a9ThuCwNtv8mD407HrKJHzr/SdstloRYmMIDV
UeAgxXT6+5+WmhEaCYfr8DbAS/8YM7Ey1w0SHs4prUQRpGUD5meiYv/Ee800JalZXVMJyRdCDCPK
uGryvaYX+AzWeFga96b5oMABtDWKEWP/dNHxyIXCxBcasVq4h9ThqOgRoAOogT2h9TWsfGiwJIUC
zCFSsXzzqcZT2IlmddHm+YYapSqfWCO0GOPcLqIMCuDHSrK+ke1Iln90OGTlWVxVziZOKc3vIrNP
G4232LEi3a4YR31poUfPqBtSJwjq5pHeE97tChNW/HApLx5pY2/OIFRhNIY8JcjGqaGQ/rspvaPb
qKUQTpNVDvk6uTe+Fn1StD4qGIf5swC85KITZrHXJK1XEK40JlGTZLZy3PNNe+dtHED2jNW6zvZW
tzzkktas1QDlKvIt0Uj/IhiY5gnwXna9e+WCwvbbTafadSQfbejt+fqw/4HS8ykarBwTnA6jcz+5
ZyCpi6L/xHyUk8KWOEyVIxEMiWSwVJyvevnA3ZICqoH5zNJsmshvWANkvaUwc6ByXJ1wHefpykaj
E9Xx/YnT6vYkUySQS1Z1aPEwXEYs2NCvElQqFsUMIc+Q26w6iYLejW6NwAMbxCKKp0VJpVbf3nGI
g+Hn3jrCeOz0bj+KWKc+w4459NweN4iu3lhACnU3jS5wxXUiSNnBFUHhbcf8C8JYTP6HfhAGSTkz
nPcCgPNfB7XqFwSoxrLQ21v+hjPz1/K9v7OKE0dzrqFdFzOr+R9aI83KBmvm/DkvDY/j/Xpuyndl
36SxNFfCTip72uFTeqnGcifop3bgAG7SjFBk1EfvDigPeVk0jWSfdj5Z7sQafSF1Ouob5WLMQ1Q7
G6YLl4BIir6cdYRwwoihLZwUiw5b/t1++JYYVvcd8ACqUDY1ngMfs8kX2aZQ3s+XSonAhUBcGAWE
qcvNyWZ7KDcsh2B4Apa/M1fXe/qJaLqvZnpIKKJ4iEwD+slyo+lQThFki5ueoLbVS7DDmBgBYq2l
gyy1ZsUUQrrPYv7qFSaeq29AuA3duLRYn+TD9QhnDq79PPDR267H0KCfGwUdxY0XbBpW3Ta1nKJ/
l0xDiJ6eEjG4sTrVGH5XKDf8A6tAQBcK/j80rstG+U9W0gVj8GoQhpDOcWjlRiKlPHShkJCAP2ub
y/6qYP0haUyj2h6y7abwl6AI55AJazlWLn8Yes3Im2+JrTvbCVzcoXvCHV4A6nWIsS7OneM9c60q
B+wFxhFYJpIt2p/GGsCWtKi+O0rwhmMpsjU3Tw8oxTQPSgXDvUMNj0qXLSH/V07RJygebjust2+K
LTECLiwwy1tzgBnLG6E7brLiSh4wLsi5ENEevhxKac7g1mvUtKmAvsmX82qzk20p7rUPisi1KbCZ
SDMz3z3/6ToWPpTg7qnPRzTfvJscizAXnxxmXN/ejnFr31YMdrAFv4qmq3K494+2ZW1tiFA/Eg/x
HxlJmwgCsh87UKVwDjaonYwXGsNZlTw4bQxA8tTdTbUfJRntAxb/1I12i3CUm3+xYyhOXwgYSZIM
reedQAKu08WLA+4ComIjXuvgvIHiPNyNEiA/pPkNC0yAZorc6RKiB915N09+hArwtuMzCvAgt6sE
EzZP0vJ2vy/I6HffHtXSRPqeLhFje6ryWuXGkNQvIEiUniK8pcd7N4Okjhjn74mkPnkeyD021e+0
LcLQf0A1LPdiPAullOrDzL91JUnkwPG+e6hKdPscvWAdLlNMQJETpGDZQ7vO8DI/ihCSDos4dEPM
BvCFVk43IkGIk70611kqPf8ItwWeaFQISLXFydyW8SstdItjR9ZfKM4XYqdxDNQJO/oCAKy+7nr5
hcCQ4veirINxV/lyxvYTuFGhdpTbtcjqwwVIaWN9JJUB3k5hNFYV6u8yfla/XHai/fk+GY6aC6KG
gzcrV6xxgXSKsT6HkabBEPDgeDFNyCwAoKSLLi12QcywBcBJddzmuIF4qOkJxvsOyWimxEKwaaLR
0WCULFD+keozO5THqO1bnFK12UAIT9ThJRappW0Su9TYOXKfCN/jAsjjclqQhURm7ceQMMk1sT91
zMOil0J4g8uaapAKVOIcz68Sq1W0k6s69YipoA/s8JdtNbtYu18gXnndLGAz3BS997Ll9mR50DCC
plkOYLEIEC8QXHpkaeepSjCJAPR7iVc4u/i6rXJI52oLyXZOVDmhfLtOZRhmBNun0peaNPqs34N7
Xuci9c+yhi20h/Fu2jnzkJ0q7lVUtlOLt7NgEt/PDPwdLUncKbQhyXs2V3JWYsHThXoO0zwSlZA1
QhrmSmMxiWC6DH9Q9FPFzQ39BxCGBv78CYWs4YGBqsXxUA6HzEcAAs+ta+0qQu9JLRlxtGBKbq2h
mx8tSmkNoTXxApjqh6JagfE/2yyD9UsQQ5wcxDPA0T0Fw6+96iYGmsJPSZuPMuxGHBDO9eoclf6F
f6M8n4mTzlIlNsC3zSE7XUOylRaYNyp7eLySB3ezYUaGlV1SMeyFLh95hRFz2rSIlPkmBd2eDRbJ
+iqOW31n/6nXS9HEaX7w8uXhEnfknycBcaZ4CTBRYWsoozzejQVE07O3c5tEeiCfPCRMbF2ApWBN
u7gEbYkn03pdGofAcpX33HW/K2AeFthWBrYpXg4/Kkby+AyMm3RJehJmOaCyjdD6BdQFRlMt8O/7
/K50A0CEurWT9+Q1GMr8s2NWFgAhktsV3NCHKafsT7kEFQQUYXCx/seeRjNIlWm8O3ynRiLyi2i9
GkiBxIb/zFIzo30m27YtuAkuycW+2I9IVR1dZycmyaZUKmGYwQe5E/95PNuKbq18xq1TJGbAPlf1
8DKV/bTRErV0DKnJgWMBmU/x8B6Kz3t0Z940aP4PCGsS+VgCQiaI+ctwLXv5OJnPmPNPLAFkoAId
he3h5nLgVRqT7FVpcfddEbSf6qWgi8Lek9/c29GIu/nEOeNqSSJR6x44WSzbVc7QUC+owNPs2Opc
GCocGexrLlelWbuIoFtlIZijqH1azQkx8F65idvA/wjQlw4qyk3BtLtMjEVCzSGbeSaH1FW8w617
ciLhQ7mnrICmuzEkcNzZFT1Dt/mMbXnO8C/UGWEYaWqd71bFhBjS+F1OKJ7ig8qNlZvln7S460ou
53+4bDUrgtiXUfA0T0/wiqspL+rQTkOuBUYNkBNK6CKHC8GQdPBDA8EI/k/bqxPQx3c4QWtAeGp3
RCJ8xNHPVKq4JZZ4Lql7H0yzLB8zwU3l3hNJ1gELojO2fBrgrUD43Sk+YUScnqZgb04c3Jokouyk
DJ/v9aM+OX82FESjOne7y4M18aye33nhI3wPmy7ryEY4SLW2GEw4+K8xtPVSrDItHjjX/oZlyjI+
ZOluA8INOSyY2yEIYoCT1n2o8U23WEDrctPuTK5B4NrTza2aHhuxKLGnPSn4areH5NaRPbnjSaKk
UA4sAx88E9gVg7fhJfq8+g1sBpfzWWQxTTGvu6x1zwS4Bb5uVsj1bj+LyEa/Ne9MyRfDjfeXpOt6
cjJZMoNc+vJpv/UVUGisOtJqeP0pfzORkfXELHZ914PD2pUGRrAVV/P/5rBHvP4G0He1NM8MIXLt
HWRsHexnmhj1xnJi5UAzd+uPc7rF6e6x+ym6sgaLz2KN+PnATBSioqZftXvDcfWff38OchL/zvn0
jcg7JgdpOeMIQm/DQRyp/bIXIpWla5yZYDgVE+YnUPhF/+ik6Vo9DqQ67WTMKPq9zl0CO0zqcZhX
bbD/XLuIN9dhO4I7ckQOicRoY74jd/sJLdt3tnjTQMQjKYx620PUikhXiz6TLBvAK/kZEqKkStKn
E/Dqd9heTNB+xWmF7+9ptan+EYFSxZHLNHr6VJjcDfqd5PS/fDQItzTQjwde8kwPj8H85LetIlaS
0gSiphS23t72pwivTeToxjLy34h9/y9YIE1sf1jxHeIMLRaVH3d3YuED+3usCxTU5bA7Xw0uhnKn
pjR29mlr9z7PBoYmGT+l6m77tRhdKsR8MnlxzudUj4j3b9FYO+hQyNsym8TkZeiG1be2M12tvmUR
hUZKJ351IuesDmOwTU4enk5BpjQI3ROImNZkZx562GOYHn6+Hu227zJSOYmuomPTtxBgZOn22Tp+
pRjDS+M/2WkgBxtrNRndFc2+au/jiVyoeTHx3D8UH7cS3s2d8i0SaMs1tWJ3FPiPNcHIkCtKr6kR
vsS03ssrxznaOCyNRzgs0aB12T75OnfXm3+nmcmn8TRaadlgwLKXcl80SRb3tLRu0EGU7puoR/rr
X1VoZkt0EZGpr2Y3I2Qe1zpFtCfJJIOJZAfoE1j2kKqjjVjpdcDYrLunenACsiuj4NZS/JvgoWjw
pLyTa+Uf4rv6WczHA4wUg5GlyHhnQMXnqOj+PjSlgb4yXHBANS77Pco1o9mgbW8EAmzyK0DWA3Vo
zRBgWX06kl4NqF4XzIu6vtAt6O6QBEq/AY3GmYTCZ1Xrrqik3WgNgLjo2U75GB/Yymr21D3rc5K+
Odw6ogzwn9DyWdFJ5tdBmU0YIu1KrN69m4hMejkTVPxcelF95nYMHG8aoV5a9AhvHEISIxKaONv5
0f3R/F/d8QO6+I4PbO2iJKqGXJaeQ+z0WBvDQlXQX2UBXKRfRodp3d63oUn/GvdAXdABDuvE9Am3
rutvlw8N1LFQVE5ogWYpg1zeItcc8l03lfW0BcVqW+PvTRBvZXXjxj0OGQmDG5igXcBdmb89QeTT
UyAsybzt/0tzw13bqzSFnf6GKfxRRoyJbqNWYOq3KmzrivRjUo5lcU6t/YqKvnPHHILoVCkTjQru
fTaa3DFKwpoOkTsEmAsJExCx/VeeCaCDpcFvfqtvDMqNZQxwq5YwxZa43aSBRs3BmcZVb+T1i9OT
uuF4kaA9I0TGy6pJ1AUolhGILDY0XF1eNQSxYGDCy+rDAFz35+bjQXqP+04LNTR6+ypRvqWBuO5u
LkVXwb3NK/AcEDmj4fF1RwaJbHCFeTYqv0yFWoC+xtnGuoM5gJGRzTAuhtPILvrbhPgS+ObJYm3K
BRlsF0o1klKjXIv5VrS2WEjQj3Q9nsF8r4LLKLNVs6EbYaxh6aNvq5xPKFwwWLCEG1inQhNVnIJZ
nYQkiopMWu0k8ObAszEfrbF+kXzfZbjkhVFwKBEpX+3kCJYBnAa8AGfmk3sjt2ECHOc+TsUwEb/N
gRW14efSptEo3e1c0mVwGLADCunMpbYOoCZZF95rzyLSnorcr4S/T6q4EvPwcaG4SY2fGJ25mDGx
9F7QazkbEr/ITdLwMkc00CFAgw+KUWEsO6tPr+8CbcIbb3ESit6bikTxQlC/8mS9N+kDrmqDED4a
VQK9o5rGL2TEKxXthMutyr0yCI3cg/5GelFD/vAas8S749DPGI7+Qgn7EGT60/3yvGNeG4adU47Y
mGNWQJQhjRIZ2pXGIKdMfzQk+C9OAKCzOyQ9jGzOvEcDuK3APK81IWWHAB9vvdunmu329AOORDqw
hBqZCTeBoDRv8/ER4bbSLq8NJWHC62LiyavCMdfFxlX3PPA7e1Geqc2Am4au1335DxgLCIjMfA1Z
8ZXjakQ2Vj9ZRRBB6MbQ0AqovmW7LsqMy0PIfIhfewfZSnASJ4b6DzVHS5Ewb70Ve29FDcBR6vIv
/jpvmbbdSc+yehOV7GU2Ihp9U9ONXB5DzRIfkqjt/6tbdQKwcNRD4hxTkhCjNWdfKBvp8+N7zUHt
fTPT32MMTiIr0QXximXdk2Vv23pfl4dc3w4jnd8Ea3RCmxgIkCQ8FIwaOCUgm4AMAgi/T6hmFKHG
z2keSsdOqAK590I6iXRAjCjWCr1gxs2UCzSDgq8NQ1zmVbXN/G2Dc3E5yeo30LDkExhJY4iXXwCm
s0McLefOcqhDqPyaYlKjxd4V2kIUVtEm6Z03iBC9H52xutUgguqfec+zAWRuWG5dpTqgXnlNI2BR
gMmY/FCJS7IrL0XAlJFJJWM8BWfBIKFwLJWMIvXcq211wph3gMC46wSs4/WrZet7T88tsWiL4dXk
kPmgzBtLnyNsqzmNvdza2GB5Op8IoAAKLxUadMVGXTjlOtxpef0C8i2EaE3czyLauA6qfkdjM6Cf
wWeKQw7lJJrHN8vr0WIJV3vq+hpLcEutDOt4q7PDoRSXK+oUfiMIPX7vVk0PBkOyMrXcRxVOCnBP
YAHSEEwofuAxgHF9GZwYxCBPg2Ma1aIwaQJDNkMjvd6IeVgHhSH6nGP15zxBKYa02uo8EEKDqt10
+n/IjyyNbxTQDTf4zbH4CKu2UZiFuey1w+MJKliowR0z0hI6a4+/mbtiVI00jO2Xt/r6PA5qnzu7
0Wlq/H+RhklrXe0VouoyKijd6zGzR8NadhhO29p7pitINw7InnwJ3b4ycRhN/VCOFvYQX1PFqkHc
/u0BS9wR8CbQFwaYWnB7T1tC1yTGLnQn7709Nu1XkFqH6GKcJpBFEwpCh0qouH/iPVey3/5Pm6OI
3sDdoMY6rfrceA2JSgsDqTf/jhn5MCduR8NXVBQtf9Y3hUKFA56XS19k337D245l90dXKE3pO1vn
QH6EaAjkGOtJbdKxesFfP7i7pIIrUPCrmiIBnzjEhHdGpRWQx51wEjPXJgNQ67J8aMIeaWdcTTJT
YcYDqJG7s89ZDFD1o7lmNDXZDdz4Kmn6Bf5oT+FkZT1yyS3b6UR0FBGD6m47s3uh5kShGKZopJfI
tGkd11NkVEY4v5sq8A8DZyDq1X/hnATdERKTaBB625CaEsbJvSHm5kqaD7lLPk5jWIzSVhja5Bg+
Pod3fY9ym0vUPnw9d1Kkj4hyvJCmQfYV/ipweGJCgLjNowtNqLI4FcI7ECae7gORzcc9Ap3D8LR/
obYajr+nBsO157ra10kDM3MDaVXMatt0T2tdP7XpW52aMvCNRoMnHOqZ4nY3bWzr2Hhw11zXgyH9
4GvFxPYzOpaaSuDCUapku8pKusyXnzCsYFcEVWmr/1Sd5RYkk7zu4thr8v14ypHKWRU+VBqsiugf
SPb4Mg2BT9h0SfZwBx/+nbxdF5VafxtcahD9JvFzPBXlQgMpt1ANENdTFRVUfvGWtcryKVs/Wo4w
jg7yJchWabI24bR01+0o529LnHWiAc7AZqc0QJ3qAjoXnRLZWXdDly8mcWOM++XHjU93JULpOMmr
5/Vbap1ma0GYfdrBvcITirnfkUh3wPV+pJESFy33e2h6jKG6BauYy0TkeEQ4xGN6XS8iXyEf2V43
JKeJHm6lxN75HBPG8KYOMOROK39uwQVSswWgFLBsjW6WE8HqkzyYRPBZdoBVZOgw/8Ax730sCKHV
CDumm/XVseqWp+25qP11Wom+5DoCFEUwTBSMC62cYw9hZYRaUCRDJ5ak0e8N9bDybimswmcArcnT
pcib5iMBT+CJQvMCWINc0zhPUykDw+Hg5CAB5IKQvni53xFWaWirLxvjDR8pZ2oOEoQbDaCLMuox
P/vEl7gtMbBt2VCZXGAy936FfQI8FnNFsBa1gUVW3chyLIcYIK0Wyze7DCZnaIE6kmpuOd5VxGfM
eVntlGUsQ9kvcDz/ftSVR5Rj/3SDMYyiBB602xXFgT86qj2YjzoZ42nvDRPYNunWdFaIMvWI2/bJ
ew6p3oSJqDxDrQDECbiTDsVIN7ZDxWvajlyjipLbFvpgwdQ7sr/ocmK/PByx9MiWUIAkQs7youlZ
2iRKh71exJ6+Zt8CCfBJM3fiQhcUGDSITT+9sjY43thQIkMjrklZ+xmlgZ7SBKkiFt23/lV5+04G
WshaHMReZSCE2DHef9qAJftWMZRi+suC/WbLU6WlU1G5YnAh/R27PnEe2B9WBmeA7LA8FqLlHRNx
M2wkSLXlM26gqOsKSfaz2MOswLNFkMEsRnbHCf4Pd/QL6kpVIlFfnuNxSzJOB0XkrlLYLS+EDMWF
0V8H4zU9QW0VCJ9iUUCK8t5fefk0Bd51AawLnBuQMln+zfySi2nLrjHrbvaIfNOBUVfO08BF4c17
jzD5Se2icCa0iiwullJvbLF3DfiUPncaIktV1V225Mf7NfBYsE9eMsCPBsF4SbbAQ+czcuyaiSEE
S2OzU72K2bzXM/ZmZnMpQrVfBJOc/M3Y+JlF5WziR7BtU9+9oIdhVNYtXU95b/99P261/rlwVgea
IEpQNsjK61NOf5/k5wSBo+hTC5VleAfsdy6K5rqv+n0gZk4/duy/3bhSsKYyi8EPCha+EGxn1FQs
IRyxjhBkPS6cxGEv69XaJWbf6FzMa20Sj2r61TNScrTe5Pqu79q/ZBA35bF52MWW9s+xPPrcJVCe
CTv/vxFMgY2yKUBWZsCU1JOhn7r6WKqzPI/vojExMTt6VSrWW2Wq1QdLZ+SPVKz8FWMoIbKNV8Ds
nAvPXF+zk7H/Mdqy1IGyy+fT4ziGqz9mRPJhfXqYxBQ+NDjK+fzENUrhBVXr0Cr6kv8wkFLZO1Xc
bdiaPZLEMM+Kcbz/Hn6CdfoCIc9n5/XntIZLmrc/gmlhE/GuYMI9Lek3cdjBe8NVF/lpZC9xxk64
SM7fQ11hv6f0h+xgGp/g9S0fHbWUQxt52TnGO7/5bFtLPgLRmA5Oul0OMBK0H+iofx66SqyYo7pR
4WBDLYbYttYCeszUwmTNAnAs9RFGKTfTwsTgAuPAaFCh4i6sshttzs4dmjTQb+kEySpE6S+/2UGb
PBtlhdbM6s5fo9ytfmbGAJEOgNrcynbEeA+o7VJAsDAbsdWhYfzjBOVAMEXJ2p0296TRn6XzW0se
jvFUXVOHmxQ7gEYA0FZTtPglB50lA3QYJu2bXDNIVe1onXZIaFctt2sY5TclnL/L7vrQM3ftR3nE
mOVoQZkQ4p8jgf9+EtDthx21tWbEhtQU87eJQaWQ/izh5ujNfnBuxGwaulhSPH9CcYDTbqRCbfRd
7tgGouSLsH94RuECAiByLxYO/hBikpze0W8EpbYFYmPn2m0h54KDTLRIWk6W0T95T6GLXJubZfeu
9ToGErfxIReVWGxb6UnuTSptRV+HjQkxqcfyx1yy17D6QlxRb0ccH8CitlwPSsaDtIlCqM2gxGAP
AY8MUrktqyJ49CUFUIjLnLrKV0zjU9Ad+9Zsm+xcWYPMRKKTPpb5nuBMSlVK4zNfSTXQ4aWAxjBx
R+OTGivXEPV/AvUoaPEjuWLYy1XFo5fAWt/cRR437OAfsT9AlrhHes4s10th3UluOYOdaOMo7pXW
yglGAx5A/l++Xl0+d0LPvgQc/DLSZhx5aKNN7ADemC5X4DaK4llhsRvw6gG8XLAqc+gQG5l9ECYb
gR/UQAa0usiup+rd9/WSsA8kiZzonOh+UPCBaPLA4VkS/AAcxSD1GHFaOQSqkrtA2+OGm7PnyB/E
k6UCYz4CIZdWK4zf1qCstYJJmGv/Zm4Zavd594BfMyDGxtpUxTYnsWbmk8R+RXG/x3EnYbEStDNY
vR9RDmdCCF3rrQ+qXzQCCpae4vks3s0xu+++mztCtlOSMXm7BH47HDnXYU9saoTqD1ioDO7NWRu/
Hw6ryDR5RbQ6SKQWY+LXgbkae9b9eQUx+esQoA5fXfwRY3DoKtpDDpT1Xbdi6PJOWvxLs0fFxQG5
UwXqoHXg7elkfPAOoQj5zzlz91ojTjtAqkzX5Dt3TGlJgU6ITtU2lo/775W9CJ5y+vos+l5fR2Dq
7LkkmsfGjSP2549XjxTdH7Tx+mgWzySKLH0kBuC/UXVE8Bnq1NlqQtu+jDxskL5xl1AqI2vT5Pqy
q51l/lFOnNIvygMQJ9gzgsqwD/P2T4SgRmtUWtdNCS983AayNxD5RtgD+aKwrJffw5O+danCC7jT
tLbPU04r8kP64m4GdKha6SQN0gPe65H4sy6ixjUB8gjEFpLTkRBFBsht82ujiTo9OKzS7OIwzIDg
EaBu6bnQ/Y9TormyNXsV8Y9Vt/SGnELvva8AzcpRkEKK+5izM5QVM6/OloRTIvJr5zy3JnQXWie/
n9B+/jimT4ktP3EzprBWDGeqwVBnXbucdWfAbNUrZ2P1DaADYDpUVeyqdD9CjsUg2NG8GWKb6qHm
8cQqwRFL9pdyAwaikmOTI7pm/VH7dL1vbFGMNddbh9heOlhShP/mDKNY1KbFNXHcYfbuDlihWwb7
GQ9+RwW7p53P+3pw0BAwKerfSI3uY8mDJSD+tCkvyq3fPlRWQXxs+WxkpClZW+e/sTGTPzUg6OSO
50PH+oSG0C+xNWI4k3AhsVcXaRJAYn9zfWxbPSpJhUp/iK1kmdxlcOdWl8eZT63ug5u5QhtQzqza
eneETMZ5Vzx5dzptyHCMVTBo9nplWv2OT0m+SbJvWUsWftiQfc6+OGCzwaCLuQwvQdEWikvoCkM0
84M3wW5tV4M1YCTqRDte9t4A7isWNg33iX1LMYglTzI5tVWHSo/H1xv5ZfpMT/6z2tNWPFuPMCCJ
iD3cCR0S5bFdVMWGGi+bl5pZtoa6+J46M6c354Y4gBD9bTAIG4yQ8RaaBc8+jtb7d07QuAD+GPMZ
T6uyKL+UL/EJhJEhkZWUWQ/yLbrLzEi6eOvjqbGC92+cNvCxN6DEAD0YOJ/sfG3Xgps2qHbVDZWm
0Zpc+YVcbKak/mtB0hUXPQaTha8d6eueVVgK4DuOcxV7mUQC68XKlXaygmqH8030FTRN56okxJpl
3PN8F761eE0ckSSrHqKNdP+ATXrQu6E0NSzUbwoXitcY6MMsZaq09Z3gMtNcoFrGRIn45tlWSftX
4CzZ66D+kTYuWO2cMpnBiZZebCssCnWTJ8wgexdkrxqdIg5MS9JIsu0f/YvI66QKjmUPv+c33Xv9
lx6BgFxPb+TyoRlxEc0F67ypigtK3Fu14KD9P4uviGfSEp8rjO+cX+XTXiLZcqw9MfEIG6kWzbqe
fJJEMlmsPiYxZGhrUfwkslgg6wgYSzD4fVTi2ObVHaUPVXSm/HUMsp4cf5DfObmHcELZpfG8U/CP
RWb8o6GhbFJvxlQm2AzurXeE3bjTAtUqOhrccoveX+I//gEJICwbTiP5FoRWkGhhdp1U2zIylBck
UrJDnlOkf8eHU5uWIgRNqg6FnAHLyTBazagCPmAnOKJNQTX+q0EynNQ1fEGj6Mkux2l+IqM9+is5
MKeDCA2k4b4H6JtlVT2oAPWuU3VOztfQe2a2+YT9gTTDmVc8clAqwG87WlNqskFLaVrUY/pAyUHo
YEb74NkVXOnEhXvpkHbBcPrYSYYlznHlcumcxFPZNn5VuZM1iuZJTFzlwlutLO4a35n1JkMxKw9O
HL6aSjD1FiYi165voX6TPfE6Tqe+ijpmFIH4LfuGWAsJc43PGuaEJD0ZoTGRyXnvZh9B3y43XlOM
nbcnUqSqT3guTj8hRv88vJGI6ZbznpQM6FkTiTUI7o93v0nVI7BQM5NiRxinlbqpdxHNTkUjsPyu
0d/UyHR9E3f9l1hTtgLNxfZymyldbQTndJbKhmvIoljNKIs7V/jsP7Shcl1Xs+YQXnroNYn/ExFR
kwZvYFSULZS4AFRQVjL/NHasilGzn+DsNFknbbzHfDNamLGkkBT1TdpUCn4OW8r8NRyOKuRB/cqW
Rdy/PPksNGAu+9h45274xqAiwkxsLi7UQXD5ZM7QUh8qwLEkgxG02SOK71OFvBTzZ4m/dW2smBMg
MhPbE1eWa4Gm27XOIIkPttmxayl9PrB2xDCUvguTYuCLBwXo7KydTNkl/BmoKeSeURcoZUgxZ9bg
TnsJYf9BF0n76agTpiNs9WQjYc+QRwJEqzX0Eb6G2O1xnjjl1iAVwr27BLG++CR+w8yaoyJnWMfj
s1QGA2Wu8NLAtXP5UjOyeIVukWBSuVLcdjgh0A791sq7JpOc3CHvjSJHhv24oh/AinzcXAqXVliP
LjQG08w2b71o4km3d0bhfhrZI//eQ95sko2Yw7k30DDj2j6Gg/FMMJMBSds3tZ5EAPmRgr91n77f
ocLP9j6M+zI6dNYdpSmGWYlkgWTCuw02Pb8UIHxkwC2SaYbdRGmCx4W5WfDzUEXbOqrdyxurXWYu
dylyOMhrbRE8jf9XU8EcWIkIoAsULRbetxyw6TVC80t9gBqNsVA1YAZBrXpNR7jIjWcLLuhyhobw
c7uDPIAkmGy3AR++pLPN0022tlHU/VE06GDVuhzvjWXyQhXU1XOR/1HH3KXL/8CRKlTokO/7cuPy
CcLHpa8s26ZQCUWZnzgeH9N5QezHGjuIpql+dzWVvzUyU2LAJPAxz417DN9vgs5XkHBqdLw4Qtvp
6zRv+auLgrTXRTKEDLh9cDRXxlcgFK2zBuW+Gu9ksipBjTGJAB4O4oCXQVf/oe9pq2ewG3HJDgX/
CpsQ5/6MffmtmUotrViR+r/4U5i2zgM2K44HxMAe9BtrkxHsSnkbTB9x+KhfPZ+k0pMiv4yI6pKk
tGcjr2YVtIwNXpYYpYfTdDOwdIo6+/E0s8ZDl23/YLdfP/u3G2KEZJY6tMepGQCha0BV5Fs3TpCy
WX83uTLo7dMlhRr2QRoot4KjWww499bHwzLpnS1I95CBPd9VEsEhhs3DWF1GomZV8PtPShaQO2d2
atx/h1ZFcRjNsb6yPEI8SbCXjcaVyJWMqYgKYHMf17K3Rd3YJMfGZNeuYmYXpFHD6FTZrWvxuWbX
UyGhGuRgRq7CQu3WrdqCkJ+K/0GQddn+JNaSkHng3wvEWqXjtVve8UYqGxnH3wDpXtc5t7LDHUdZ
/HhPJOzZzaeVYTQXt3P4F9d4NS3ep097RfawatlpPvnddL2zjgnp7FfX1JR0TYObZYk13o6mJNjp
j8DDCoepgIJsf7qems/qFKIiUaCGMkdalGy7tNNmbjYUk7ivXv5NjhC+rhbgV0z0L2u3MGesTfrm
JtEO4u0UGouqo8JmxDeaODmW0AO3yU+KutPimPdJqRvhGqXvbRgrQ2Ku2eiIOqoHeFGFeO/JATIE
lOt1pF5/1TSmzb+TjgPLAZmk5CdAUSAdPtdDxadTROLN3NhdOFeGF3MGkUFcpdDdO3MxZO0lmzz9
cxpJOs4d4DKUHgQujC2mRLjYKxepDxCsSUUnQq+DX+FV4sLGIE3hcXpS9vQd4h/3maHboniOJGnR
XlPqWTTgUowKhq6saZJn6CInAYE9w/3MrkFr91autnMOxEh17NJ1YDCnPiIC6mopy9mCi1bbyv2x
gImQfLav9X9SUG4ksQ1HieetxXOSVokxSZcSPaX7ryqrQ9Gl3k8fRmmErygIHgWpee3AGUEeLp96
/J5EC066Sj/KHTBkWGB+za7v0fi6EWNOHpopyrTtN83cu6d+yMqNFTWIkCc6A6aeR7rHzguCXfX/
jNlldRDwKsmcnXUcXJCjHdyzzaqJZtdA0/NfQe7iji4uo5crMwj0LlmMlcW05xGUUUTrhimRwsp9
bBm2R0T2D3oFolON80z00FeJhhUspSw0yCgY0NE11/bmyqKr11GgVsC660r5e+658sTFQLltrVVu
87Fu6Plx/XCHMwS4nbA6h0GbY/7Ol6uWibx3XSyEMMInQa88DpKnWW8z1cpYb47FPSIwsXVLLw5i
l04/XNq7kLH318K+xJBMg6US7gfM/n8Ske3Ng7ePTGw5xGRm4mumaxOZOX2xX3o+IlMAz/G4Kv8f
LesfjGKusw+3yrnd8NZaL7Y+ZZ8DyjWtQMIIJnoPgh2MjpYIoJsNKDY+heD9/DOEFPuDYl8WtP0J
Ib3bVc2dHIyO/YvHTUgG87iOem9tD7LR3yOH4352NNlj/qNmvMJRnM2S8H4dqAWwWNy/jA1i6qG3
z7AjlHeon2pjz4l+tXX+cZmSEHiyKwJd4b/lVjvbPFiQuv/iNjmVtj9uBvr1Ksac3ZNo10ee9Aag
4xasOI7CA8/Ihl9q4mnSqBFZVT8dj5vfS5QhtorzvrCpiEPkSZiNvBEA7spAVdPhEyTkqLtGmx8n
+mDhk688MaubGSNfYerGErKPXcvlSC4d7eKehdaCPKW8Bl+RtpnuUtdXRxrpnPUWXxF1RbRsjusI
OcKy+5TC/w9fEPNla9dWH64cBg+nVpU5dL67wIVQZyBR+gsbjsB5gVmyDrqdPkfr12OsHOAzsVEQ
/OgX3JjPr82I6MqUukpFSJhZAI5AWvKi5vj+dGTQuMGnPs04Uz3UHm3FSxKglYDOg02rvrJfSeSR
MzEHLJ7Fun1GdLXtlb3WaQqwlZwHEh6VZxJrapO7DS3Hnj11SBYvoYwOcGF3s7F/KzaUR0IfC5eq
JXSGjSMZk8pHYthEoK9WKMYHUnZdX8giX7AId8qj8C/t7rxYyoDsn4ZSC0zaAbXFWvG7Lj4YvDB1
B1bqymNc5YSAa29gupbyME0wmlgu9eOJse79it3Llc2SjOEpiZ9Yzew27Xn7dM3ha8gYoLFk19Ez
grYACv20Eo0bgLMol9+3dHvfcHYunC6GEBi2nPBrH/ykgijh5j7+Uo6vt///nADX9TGtuLAy4IO7
MCYIlZm73gKdBRoLIPhpxGZKjuU6RIM5bpye19aUdB+BX3qhIDSPtiidiPLqWP7vmOX1GnqNdua5
P+OTGc5ppboClp8L9nj8CCe/NOW7BMiVdmAGJj/J8R8ZlBPHxMu+Z42bfjYk4glRjmGaePEmQnGs
2xgGyy2IbgGWASyw6FPQ5GD0DLkWST+HwppX8kupM5Si3CGSWdMRlPhztxLRhlenHzzaSFXjbrmQ
dkJRcVpZwdRaQAnkuRjvuAQwoXzCNzygYieyi91XuF1yw39Q6TEs6wBoEPPcgO/F2tsKQVUXHjhn
M3bd7/jLio/3eDR0ooS9v5Q7MkWtjSv9+Lp2QMaT9vsDFZUoWXV50dqusHT5DgIuyNsK3ByDqLIx
mPEiQPrsJaVQJ+/znfy7E9z0IXQSncoBWHeErnzL6e5OO4IsyjKIr55WqCIP2t8Qi7WSyGjHxiPl
Ys+Ez/aeOXiXYrcoHqIgGX5iVGVpeca/DfmtEQ01S6FDKJSriB6Z3zRmhGBZNsNXZDWdc4SkOiuM
zfO9gcDA7iy2sXFMhNlTdrG8lzSkz6lpOcibQmfNw+29nPlxahiM/oeBR4qoGX5Xdwo3KLW/NU6i
/661fADvQO2i8QICrazmGUxT1TGwvMv8+fEPnw49+sDfwEPfxyqPXgNi7TqYsk/1WjGm5UGB1JSD
Ck8BVhWQoQPO13BnG0u3F6YnybNoszUOwj1Jp+3PmoXbfal8YQV2cSPKA4QgK8JshsI9lDYFKi5z
qeeqmrFweax3XaBxlduNiiDdH6D7RKJV5tGdziCno6NAC391WpVQnEIiP6W1zTm8O5IlBpmCdmff
cLcC8hoAUY8n/fGpbnYpfm5YYtL3KzZ43O95FU0EFZCLKv4E/cxSQdPxrGnovd26C5RUdRCdEz5Q
R+uqeuEDRYtr9VyoY6ZMwaAjyaAad67xAByIfwB/pPvdFG6sgLjqyHpQRdYIhuVd5zKgsYirluEb
iqy62Lp6ytYF8s9PlpJ34BxWIjCl+COK3mzj3LzfZ5u4iV/JQ7FWOOgl3SkWgYTPPi4Nr6UbgMN6
U2KSasskOWANl/9tA3XuxkNt2/2z6/4af/9JpinDq/r4l+7zSJ5w/kPJTmob6vzUio2xu1hWQS5g
CC6dppEe6nAVV2oRFQUvkCa9FkAGslgNgz7c+fy8MKV7T00YuY0/dxjhln5LUKfu3hcBwkEing/+
h5bzWf4iFxxp70LQWwC/N+eaOcSN1jfFiHjASP/MWY8It1DxATLTYJSN4UxxkscNmexChBbtQZ5H
TT2o/5wEVh76pM7GP2a33irNcfZ2iVO4QDSsNkxRxchavpOhxPWtmFL7D6D6wBSpNOPfRE+QlMn5
Kej5x4SMz4Y18TICB1KvPWZYTVUmXzSEzXSAraK2cx2GZAFiY67okHtumEs3xkzj4le3/zMIoscf
xonvMkUacYDkYiqPvqOf1oPHI4bvzFMfWPIbbV23NFaLnJf0q4mJ0UrC6Edw/h1KZwyrJlIynCDi
fAUyx+/sNygL4DzkrhhCWjN+ijDBtzP0iacguhyB5dbLNG+7P33ozdlGdyPvL1TQclFjT881yBpe
tBYHqO6a6OgTt1fS4maDJ7tsXWEiKRehO6JeUD3o0ylUzFqCzC+BuwZv5z5LnnuGWPKHtV3JaPi4
AEaHjvPCE9GJ7Ji8jogaC1AoAxgpv9N8d+xsO6LiC2sLmCMgHeC5+j/76PLbUM6MCj1chiHPGnsk
guCCy02TXvsgVoHZxmiRficfQwQjPEBc9kIQ5X80KjtDUnlcHxccVvUsWDwmkRzsOynlOLP9YU01
2wCtU6setddk3mUeGAG97/nvsrj3KYanrOsnDNnxfUAJRWoXseerMRq9iMi4pYfMAFyYpo78Kj1C
elJgLOkH5/vCZal65mWDsigWZfXdHF7epMYiW8PRnS7fAHBF1CP8Crm2KN0WkXLh4pm+ys9KSjXy
N6+UDpnjTGG8IpZn4XrAhIXbFuwi75qBiF3ybXPhaUzJZDkTBkj2wNF+IhIH6naCZaymgLfz8FKV
Rzdjd9ADVutNNUM11VFX4bxKL618SGL/VJ7mglLR9dtHSWpG/LT0ioyyFkT0bL3yp0fv1YEO+gQ0
UCwJ2MQasyRhEw1c18j/L9nDwN/LbhtPaexUdrhbBxRHd20yxjW5lbBM8bfcJdAGl8f9B8znCWVZ
5WEELKW0WlY+J0CeTYp93vVvMCTQSmJfqjYCN0swQMpWE6GOYfHBxVbGgVt+wmj5OeSMl7ydxear
MBgaB3+BL0ScmRHu41KrV8bEsPH82fq9Ua0CXb8tdWGQkuX7hEa+PQijv5DjyAwHbKfOy0vo3rdB
coBiXP5XiABmGMUPuZHg0dq83oEwVetC0zero9n6Wf8bJ+YH7TGz33PM0pwEcY93tU/qFiwkBpdL
oE7NGQA2eXBhLOQUZbpb+4PFVLKgU6bS2hml2l5iG/wFScwiMSX45HokE2dH6k0n3XuknLPbuZVs
CWNxp+y6Kzs8gOK0GtLt2QnXAvZ+EQ+XNRHX52M/VTiNKkaPZO2RwyMGPxE5QDm+CJ5e6kUqZ7Jw
AM4eP0c1GINCPSznT4hsC3cmAzjY25tTh3/dqR/cP+L5CzYWptJMA9/YXn7oSqI7gg43zHCUr+m1
R8WSsFG10oE12eqtfuW3cOD4PwNqXHjwa3UtDG6XY3ARFezXT+NQadweICuZixAOn8xEx/mlmX63
LEHqomp2lB6Fn0BJYV5oY6wnqrF2iE+I6GB1h3cl/1k5pHzIcHaUF6LOa4Rou58QJx0xMv2n7K48
cYqdH0I/H6jFBG4qajzse5WEu+6deoYWt3nxLNXiEzpYmNqryuZfbIY7qfqpqRgsmSa0jWhLisnH
/SK8vLuH7MPbqhk0grBelEAqwMlUxUmrmQy9MuAsv60uDTeWWNaXOZIXVzi1LpGBw3YhlmcNBK0n
FCnQQmoT54qDXEdfo16SLQ7WIXpLS5krTk8GjHPuYHvn+jwaNVPt3ZiX6wiJxF71dS+GwLspTgvh
Ky/hL2xpZ71Ok+J+PSpa1SpVdqnSQ8RC0kh92NhJG0PXohOOXO7R+AqyUH4ek42RDn6SASGbbPb6
6IlttXX3KWNzX/Gxa7703T3YMyjHT80t4wbc5GHLswD7rxyo1tpj/iN6AckcgSwgrRTCdz9bBEI7
1rbQXqyzBV103HPgUEs6jXVOXQphJQqD9t9cd34tBXbAzlamoTu2hZ0Ix95DrlOobTyVVe7GYXyv
/fA6n0av5P08FtqFIj0YqAlF5jwE5gkq87IYKhQ5n4IaLdmFS8qPUbaF3QI0gsLn3OqK3cL43/17
7Ml97qLzNJKHi91h3qwR/CkaiC6AiykOiNulzU0T+jstVs/hlOE41uCK0Lm07xg333BJqLsRp3+K
EcG2AgaUcE/eCpa3nxhkpKNwGp8HCM8xvm0P0Z9g0HF3dnrs3/3KhRolQpe+X8JMsO+YD2HOcKct
GykLxhnqGXu7s3MVEhRJMDTrLQWWnhIcL6G82ZAqvhHQ/S7J60oBRemg4QzxVencIkM8hJhnfuy/
2+7QgL29BvnJpdFQ2CoHipxw8b8TYAEjcB6aKvcvF0C/3vGG6aBMXLxK0s4dqZKrZy05pPYgHRya
smHYuv2MVSw/klHc3McgY3O+pWi1owGQ5oJsPRIeJ3Zke0MZ0SxztkMDPl/dZGXHLJtqQfIZbf56
y5/NKt24fpijbYzJtACOvI0LhN5j7SeF8ay//N2Wenhqw5VGe7E7FaDmRwQTWik96wz12izNLxEr
Oa1j6UrvKTJYx8lbwzP3OgWM8P7FcPS1MSxLjPTe3MFZmHptgLd+5nFVzY/TugeyR9sTVoNp5i0i
OTOzUvPDttMQkWDJotcG/SjcsRhHaRwr88bTwOvy23BxLAjTLwM0YMohJMzDcJ1wY6FAYgnyoD5m
hyP7CZN+DMHs9vATcEz0XEYbsDSkK88j62J0ERh2Aac2OHITl7e5NfhRGCWKDjAHA3cW31X1nHdr
YbvXFdiyWIDIInCDdG7rJRgMOOQ+qk6Dwf059VwW9p8PiyqDP/N78QqNioeM4EPE1V0RKalsAHsu
coQRXfypYC1ll4JBLZEYp2p/JP0NBRedy4dHG4Iu3zNQ7XavUnsS8sf273443lgXVYovRqlY+6JC
bPMejLvdfp3ZuDJs02lE5FtL2PZ6jeFrErf8O/VMfhrj1bTJqgHVAeJ0UeXjOLHsHiTDnOgaR2ca
sQj6b+8tkiXQmfVdaK3RkyQz//7rp59Yv8NULS+WyCRr03bvVDCv3ajeGq6vI69hUeqPNfCKP7t8
+gOh54hTgNcjxAEt48/25V/iKv/Q0ID4bEypD+qj3f1zh3hQQud/OBPLU/JoIz81TxsZGEcHhTSG
i4tVpnbo/aYnnhXCe9B6OWPXkuOVPJHMkVFktOh2oGNsvNac+puxGM3ow9cwCrfvoA3bk8fVUFS4
tWUoGJ8WKdNp9ewRnxicBJB5uFMdcCjNZHFFBvzGVUmDmin+GQb9+YDvs8mypuvWZVgtgmd8g2GE
nbdUnWr58wwAXMwPkDvZ05VWe+U5B+nQlueNjaxlWL0UMmPHyb4P6yx+7moi4YgaW5mg+fTcbT+P
CEkc8DUeoz/NS308TDZDPyqOn7N79pde5in6TjSrtyYgjre5EH/Ts7CIRaCaFryHMSpVgOKn1CiO
fH6clbM4mJfOuZKyZvo344zZxU3WlWyy6PqNpTIMMzTzyB2bMXiIPTfZ3S51968wWmB3V04m9rDW
2dekK0P3ylQB28L6hXQZLcQS09p8dqXAFIz+jMFvLA8IxDWEPYCVEvPuCEIfmxb8dOWZ5R7btXrQ
AAjTCka5QLl2jtExEZNWYOO8dyKg+2yoqhOOhbooHDCmq9mtVGo0QUijUrZuvjYViV77kYY28/7Q
r0gG0QfTFyeL4VQIiWHncaFebYfOjA0wP9EdXrnSXGS44jGXAhlccVzzwYZ18A/5G5NdHKkvmDqm
MMv86hPps4pOT8MD5ShgD95zOBoKTZwHAM3mEwdDMW+DaukWT5qF/VqXmc73OtfX0DGzGcKqsycc
HtffUg3tm1OUGJmGkvyqbFFz6DlEP8TX3VwqfnkfNO42U0xq1nZnQxgvwbqM4f2yIeLRKX3WKjKQ
poHZ0Vz5qYgaD7YTzEQyutbJVoVd3kDcqR6G9yfXau1bTwu9T7wl57yjqMjDOyBgr0rXgq8M3SNu
nNhcH0yYJHW/nbUOWumVCqJntXdwZL/6eaFumVQ/5o9u45jofrClUipwHXqm32YO631l5SwzS0rd
hQaGFQJzpDvwcsFYU1/G94JUuEfQz04HIsw71joYXSsjMhWoFa+w+tjjs2WiZWD8WLkK8UtGNeJg
/4DlWlvp4ic/BeGvc2HxJ9BMpLEQxbnLrJimS/MXncIwC3uwLC092vf45lGkqJBF1q3/ncpp6icv
eQHCu7612O55RDneyZzsSsVgsdlv2fHoQPhQgwM8F3s8xcQ9UP5PGLZ48LoK7/1Vq1bGW3HAkcHw
83DGetyfrz9PW/OkRxWtWDEYxePxKrJAyhUH3qS4f7J5YNb9rScGH3pzLSoidyWQTtsPrJik2VMa
K/r5xvkJphA7wFd0fz4yRr74Eekafv+NYtCxtru+kBVpCRqCq424pXNYiLU8KlXCZ/Ml3EdmP2jB
iENBBKmMU4p1prNv1Qzr7etek5m4Lb7PSJxK7NHDrtbqbFRAbkqYvh1MBfx00MRp0YQM2kw5zjlJ
JlNQQkqO2SEnsLf0XULHdJuarc1s+nVBWqwiHQNxckpOLyLQGi0DcLS1ufEip2hJ5BWsEiSwSOh4
OaMNk7XhmJssa0BoxmCVZ4j/c0gQsmSorSCqJW5dORk/7zTmyeI5NGtS/t5Y4Y30xm67cs+PrUg9
52hNcoYxVpj/GoFBGBawQ+mAZHazConsjPuNja7cB7aksNsGo+TeK4sNUNm6S8Fl4U+XTNIHlftO
vcwb47mUaI13eKsV7Kv3Cxrwaoy96Eu8bKVowgcT85ehgNvPjMQdxoTDPtPI/P3w3atDPct/4NCL
vl0w2JXIcLKdeYbE2/O8mExuwoB/S3wjheh7KhZAKsZWSwAjx2fB/Q7mERJ6bjP+C6BCZrPidQiW
DLzXMW8hm69ATsoRBTkBkOJ7OdrEoVfGokTKA+g+Tth7H3AUsNwUk9u2p2aQsfeGWZaEAz6/S7SC
tCSOA4kNQ2ngMHjhIGMY6W3a6jtmwXuo/9PAMkvFF7QF/ADFsrC+EM726wUmXvlxBcaypGjzHZAU
HVGcN8sy7i45TSaIak0Q/OQpWXZO8tR18Bi1XlEKOAFgC/nQSgao4Myj/bV1MWJnyofIe896+3pl
Kneu03rc2cw0GCO6qogVOVbHZa3nQ16xBNE/5ehqcOnvV6053LGKzgPZIoU1asaosYc5exmJ7LxA
2Wy1a01J/h/oFosP89xTDw1LIH8wVhtPxQ2NvLU2tHHuZwo7CcC6+BcNlMinIbAZf7j72Vmw7Fb9
tJFsAVoQDqqId27jl2HRutIZsNQSUegwaXZAUWv49N2gqzof7/nuSp2yq094lQ6ETm6VwEchCyjr
UHOwe9KnVHJfUGMt3XPi5RH3hPBHqD3+qZVpnrewYYCLnd91b7axs6LoTSGCIf2BseXiOTLvyXmf
KNFZdcfuJAv7QUO1CYBt+GqvnRV3Ltiox4ADR1jJCy4u7OuXkruJT5GgGE+lnolWPsv2wOfbTFdW
3dXtm+zak1z3KeZLLM5GhXT34uiMBONxr8BOS7m0MlOmQADbNXrosP1WjVvoJ697yXBK+GKC1a4s
Hj3hb3zbqWNvjoTfBmGnBCJo9dKkGZo75yZDluXDxmbmWayPJ7l8vs3ylyknDF6TNIdFTm3jbT1m
aFauHOcfrlxKcOr/MwmT6BkRQYUpAj5Vzdd2194aK4FM5ylWPdxWLbQFlgCPWhSiH7Zl2awZhjWP
FyaRYI7GZ/fNqtPnKX9Z7sLzf3XgpV00OoklTAsQOwXFAhk8elY9Ku+FMAeh+jqh1Gc7JfJpGwQn
fxoIG4d7ofWW6WLqzIk6B/XgnvruUTUGDjyFcUyPJe/yAf5FwFHOgTMBq/Ob5KKBa2VfhoKC4KlK
nsw3fDDvyH1KLCpRJJbV+bCF8y+12QP6ove0Rb9N5kjGDbLm76XEkkbAnXt4LJIZQDl1iuS0mwRM
FUUp2+Y5j1dsph7mgXTkavlT6ao7x8SU1etDzKrOa02ieqm5mePOt1FcVfEVCWngexwjzLJcLyXh
wUPKHv7sZ+GygNvyfcn+pw+RxV/2yPItHxaMtZHbFaNqZTIifTv6SPEgAWruhG55fiPqRPUjwpFf
4Ho8jkNoKDelkCd+nOxbIY2LC5mQ0v2KuSZLhAWHiOE71fttwEyVXdEu6ONblfqzKqj6OkwuF0+u
o/R5l3k7ogJTkFDfhK63RMCwZDwGD1T3yhPiRMc8A8k96pmzbbcqi72qXEpwN7tpiSKAALVkiQHd
NiXx/A3DB4HGHkgy5dxdouhXyFQqGH/ayV1trk6wvMqcF8l3T+LFhxZKUFHL/vGcIW9r0hsLy7yE
Axz3Z0FBwi8U26MxTVmnz1VHRbwmIlQPcMbvtzeSBJXZbqgz+gngmYF5dz3jtSmN0CIyN8UFdZmd
YzvrF4Ju12344KceoIhTzIvqllttsv1hhFmjv0+9t/4GHJ1yxA6hgEFD4TeXDo06CvopcafR5QzW
T5PrzGOlcPUjJjvfQgc1ch54IbY1pyDubMM5dSggZj+nJdgYQHreWd8X5tRfrFQeLWZQJuNoWs34
BhWRq8oSQBBgrKiaRdyxdqQyp2+TGE5uPLJo/bQ5tP8d3MLVs3RrLIM5ndybien14BedCsVueeVM
mIaHK+YIytEQQMYGLpzjenQFDYmgtAZCfU0cnziEaxOod1RTybD64txbLII3HxUhsbh+dqO2ca69
xXSLrfEMoZoSXgNkpiQbmWmRpX0N2XS+MEehLQay6fejxN5sFWibI++KhzwIJJ/yHkuW6UX1b/f2
oHGQNkhLG/EYWX7aNmDeLC5Fzdxxgazaj6QrbRWzXYvdypr1G2/POSiy7SNUXI16iniwtCKtW+Pv
2kbQeroEtexgpJrZX3IJDhOb68nWVI2rqSsR3DrWxwrdzAiqQ/V0OZrwhUC+dKPp3kPNCSK9xDZx
b7tt6ZjuGCTXSLNvUQbbHkHR2k+WtZPIWTRp8C9qghjNoIQF7fgfGtB+hKCVqtlFULJioneE+jbX
mUWZhphVgrZ2+a903QrQn4v2ySqlxgHOUFTQ4zohjF1nG7rjti7qdv6eSp7JLvIKLhkhV6743HMw
KvwE9C19IHwMTz7ApEasTsQwq81UMhtIzQNI+gSPcT1Jk8bmO9urpylPKPfwC55fhobGJm5h8xnU
GdCYAMytOTiOWeNyRRglKJk7O/8joXQB3xWtR8EdvYDnod4IyKla7mDkpSRuaHRRBGpO6JJwg+go
ZFXitASw0W5nLAUuqGqxh9Jjjad2sujgvjbw9L+sLCjnKp5qaJquOQg8N8Eak7sa3Z+UyO8VWn1T
5U/bC8QWaUQZ1icWZdSD43mE6KMGjy1wImkctuh8YcqFOY5sUR2UXyBVFu/KNi3QyKYE5Gj6I+TB
VCRkTjZ/swoRSUaqzOk5PDvOZz9UHW2ZbRGCCxNQitTopiv4TPlSkPXXkvCwS1x5FmzGGQ++YBDK
aIJjJwNQ1AGmz8xzjHVzDGi19kYOA0WuMvg5p6vhD9ah9zWlnWKQIvAIMLYzvbDsXpzEDq+YSbQ/
GYMeSqPZGZGLHPYXJEbw51Yy/+vw1CZ+0BeUBLQUb2MIMLrt+c7q5Z63xxSDTwY/SoVp5LHmryq2
ILwHxSBy41evCHVdAsK71bs2zeBMT69sLV6ngWtAtGnkrp79hFXxeDcyQEoPfvlXcq1jJRSJvO4R
iehnCktAhjw4DpWXC2pooJ3xbwagrx8CB/KKCk1vkNZgDdjIa2guJzV8SO6TirZXzdY3OGek1/kq
Q+6DrEiiT/V06VWcWdZHMJSe1ixztioPdjHrVdpjkp6l8DIGMi+3LKKnUT9RbqEhAGhdoxNEOGOl
om7UnysxMfgcyLSeeEGS2GHtWcE3YXbgTUICwJzUcMZFJaeTSvymfWh9hxGIg7vBWkF8rAI90Myi
3pOLSBOkwkOzjd4dnf1cfPjwNhrHqTGkF+ow4O/w6L6y+ayG+0nk3YolocTNgISBOa1rWs96+wCK
5FL4xCt/SaeoQkc32+k2hRJJjQXsftS79SY1dgmXYzhoJH/9eQOAvV+X9z94F8oDHIqUmMsP1xGg
gD/fSyQcyEpiPb1nIRFGVPRzyANAJvsUBAirl/9M0SYAux6JOmDAhuzdJdsc/KoWuhw6vro3QQl8
XOhhukfLQGUN525JSy2kCCP5dhkKZuau3MgQ3mgl9tRtMxu7FBWweJECPyAtia8ATMK6PD4D1BuR
SmNO24yfjaY1rPBF3XCSGzirNB8615cHgre2/K4xn7HzSaDbwKEv2Dc5iUaSVEVyA0VHTt4KXSq1
YnAMfLPjAmRnxYk8EQJMirlLMskXEhHDTbuKO+HWzDNanyham+gz09GfaRL2dbLvbC+UfPgayf5r
/CgDlMBzWc6fMyJI6GmnXxsx3WgdQNG8nmN60aK5dTKhleyqZpM7GsWFvW72969+5P5397GY1Tmj
jreJ0WN33i/bMKaUGxqKzLMkLQEjav29oCkyDHoP4uXDRcJzwZFsjP54Ofh/KHTO70zRpLmljEpc
3PA/qI1ZEHNfrMn9sDPEAsKL9i6yQe2Q8bn9x62BdcpIDBFkNv1liYyMlJX8cX2A0lAbnChv6YQZ
Epgj8GhrAgLqSTxRRvw+QaXdWqMA95AKnWTh4m36Y8CMw8a3j61K4XV35p8rKEUSCOPIPF0P/bdP
C4OHsfI9aI7PDDpRFI3S7bFnCzpveLTCsTsFoZeiOfJZ5x7MHEjcOOtiWvQHKnpo+Chdx7RTGwM1
MyWJKoa+ccxxM1NvJiw9MiFg4ArxVurmE+05tSc2yoFNwlnLosgmvy56nWlOpHifhjHw64/sq8zn
KvoNMMaY8juinsjoRfH5LvDUWO9HhEBYx8I7UZnxYIYGr8csC2VzeCxrFr9gZKjFJ2/W583P/dKz
7MmZO/CKYjxwnBTKmUYUDPxkltOFXJ0l9/Uvu9r1r/oGph4Ec6CXJ6DzmKDA7v7aYhAwC7mMhVJ+
Ekcuk5DQzMbbM4sE+hcf8au2zXdSFGCN+aG89eJbYBOolqgym8ZpuStKfb63V9XztRj0kmK5i7em
sLrVHEev9O5FAxT8wLjK6Kikme7XtL9Pcv9em3cm7coL7+5RhDEfPa6Z62NTfJ6Px5E6klYYoEFS
aGpwGtIrwkFwKcjR921KZCqhTCkyLywTWRMAhD7ZxZIU336TXi6JGxVRif0qnjWiDAb6PpGFMfmu
JcXZxHTK5hNzqPo5zlytkG/03L5bbVUfb+VKF5hhKdHaNTHlJTl12mJehuCRHqSenNGiL+PdQZ1j
SgjDZk4Cnz8QHydq7Its6ZHP7a8/rjul6709JwdtWXtG/wkav+wr0PCX4tnoe99eis1Z4i+fPpDk
+gi2hfKhxOi2IcynaWznxQfO5r0nrQWoWZG57+aF0704Dc0RMbsuNtzO4qRAGUQoXfvso7QroHFc
fYfvxZT8yQtKcdhq+I/PK5sh+jKHjzxk9YmtKgVpuiiaVkqNMQA4TKRn3AGeQsVvDI4Itz3dZLBJ
2Chs8MhISmJOyiqcE+yBlfjZ1Dm895z7uL/zB6kCBavgDWtbr4pZW5qRftlMTDz5rSWPHy0K1mc1
8tIaYFFiX4C7kzDVUN9Qf+wfPpUCYzZlPvTDmpFWc6IJMoiYmcqMOrOZLGMgnD5iQRj62S6Ec36B
FcUi2Gwpcusan7QEL8Ja2D9SkLEs1snk+FRov/TYmX2GBa+X4byPUbyioEeM6WuFqhTPDCx2t6Yo
BgZsKFS8UEb/B598FTk3lErgLwuwGO9c3rvd2VCMffqKVrFTs4O/l496GNdJS7n0LMXnMj3HwNZc
7iVGCRlbt5U5HcpacSr5O0iC3LwWW+HHX6S757NX87TvFGoVAxRzHLcj0eY0m+Ku+uPqQXioQDOv
8/pvK6R1B15JOBOQTJEvBF6eeUU+XCc6upou7de/BV89FB43YRkdfxhjo30uR0WOaYOUrnGBNV9F
lV4kNYnGrYlDGgMeXZdAxZHF9+lmnJB4DxhNN360X9e9aYIRvNpj0pHGxU1tSy1Q/qnBRFStRJhN
QjSBmRjReUkGfc/sMerQh7mWQMGkxbNCu3YwVzMcVSnhGc+k1kbFed1OWqBXfiMIa9FdKvgVqdBE
Xl8laJ6VpNsq4P5sCPNxHnafJxXvowKmr0LkEhtLnzJuYBLeJI4hzE+ZvkwymyM2/iBevr7V7jDi
2WSGoe9VUdJFYf2ALOt7fpEqWyuDWIc3Mt+D3Rh7RfgNBkZYDbjqKP8afOR4aVELJVe9iAMPxNhf
9pSKMhPcJVcgYycnSnaFucwhR1qdYH5L07tr1yHCJyjlkFQqvbxpk//gtbjrOLvNlOAC/3NGP0lR
RtsopfUDfgzz8rfp/Y3xUo7pZ+3r/lAj4+jsaZm18iriOvEizigu7gwo2zCbeRjIJejgm7CdvkUW
KsUG4A6DnASmuwJIXgRI4330P8tpEmWnklyuoXp7rIYMjS6cdu1cM2ILB/mxr3k49AwvabJ30Xbz
ikmfbPbN6kt02IPUXwQzI0JckKEWrKUTfJ47ZAJ0v15CMF+RZlr67fk3WoG5JDz+ezvHn1FZo2UE
E0kqhYY45S52ezTcq1X4eU/XT5VH6E1U7505NlHeXRNfK/k2POSpe4a0jOSaeagTD6FfS4uJ88m1
gOPQIWZC6JmajWGaWI+4eu4t10ZzpOpuMAZyk+fey4KCeM4P0QjQXOrAzHplgtznlyVXGKDwoVbV
xI4PBQnErQF841b3qsarIVhv9dVZVSvxp3TlyXXHlrjlk2rba6VBHA1Fl48mywQib5zOhdH4cHdi
e4jSDDj6/Q+MLhied2WRgPiD1VC6i0eaD3/RxLqD4ahlCvJPwq3kJc+amJQZd6bAdEpqCrUAQA75
yswontAgCJqtAwXCsuA39g6rqvQYh+glW3qQg+p8PyEVNuvbV7xNugne3wp3yJBMnAESuVvvpL41
Qa5Sjkj3fmAM8KjMhJG6+gX+lIrb8erHSKgqzAM8gkxPv8xoLqDKUumaANC0v3zjo/G3W/1Tu7X+
056J6A7nJEavys8TzO7nmDsCldVR1DUmpMAs4I1OSR536fHcrHg/WVkHaEgnlxmm3uaUpZaW8zEC
m0rqWy5IYVPtvna8DUeWL64v49FuKD8px6o1gv50aKA/osx7eVQj2crf6jpTzT8X11ndVKIn49ax
iOB0+m6FyTfqF7SeGCdAc0d72vanV7bojqtVxjS2nKas8W3/jDOQHwzhKjPu26V6QKcRe4zz8bQ/
OzQc11T9EBNPVi2+ZwFxn5xah4E+BUXgAK9i/9lIkG2WHKqkvRqunFlmQ/Ky5VOccwwxWJ1+Zq4X
FkiIWWHmnYZA5GDgpKImS6ddK6/PmG1lSOoHolOi4zq2chIE7+tY9D9s29ysPIadRzMXigdhlxzd
E64YyP7qeC2ztw/65qKgcysGSH3DqJIr6kpKggV88Wq6sIQYEyZ1wNJUddw3wF93Jm7Iobeb0Byz
51YuEYwSHGhUDrO58bx88WEcXQQn4EG846YcNJbNLpODT/gko32bOiDSvLpgMyEjqqPDnRtgZmAR
RH7U7nHIKupJjxErVqIXM35AwOPhOhA4LoB8rVNZQQ8ZSfaOsGFVAtgqk5aUKnl427rfyUW9Lzeo
qRck5Ez3QP0C4lcoZIGbPzKoSZpbkZQ/PS3NRFh459dY/LoxAxV0REqN2CQcy0m04uxM91Bq75hn
InMtUVAim9sqYs9ZuUToSgwTB2VDR4T5+4yflUiiZ3HVxom5lmOfrTuT5w9ClfMsMuBhraT2LPdT
1xVe3vM/e9njOn47YMbFF+m3fYvpmoVuV34hwzPpBo6S729DJtaHaa1M2Bz3TVsZ2Wy7niCSNkjd
LAb7gk0TAGvmeBf8bkUpmHi3fzFHc3DHL5IA8CvJXQ9x9SeX5eHNzGc32shGAcUlZsMH7bmBiR02
ne8MXMZsLxaMyCq3LYq6eLYI4x3dfByhimJlZKzb9RRTK0TGeEnQ5rDEUziNeNGe6giKgW4Oya+o
oAKVj73wtzkcMhFyucvaiUjWxRaQucOj2AV00ZRQY0NKMcC6Maf5nmc6Q9nBKhbOuu+B4yvaeARk
kYVJ5JDBYc+9/gLZ/9xg5+uLa9zbnNbzzlYoIKzVu0BJs9Ua9ixfK12u8hKESyNS1tUbWJDDivjA
02VkmcNE8yNnfbM4zOmeN+5nYmyDQrfGmmiNwzeERGdF+bGL9tIaucR0/ur050K5QPIETKFk7Iov
mxAmyxKkO/88BB04DvvKFTRt4wbpHU+8WmAYRw/8nUruRRohR8nZA+J2PFJdUuta7cZKiUX5hoH6
G4MUFl2nbHnLblk8AmtFYJ+ygrLvDA+cwmnvzh+oZgdBxo+x9o9Af45MJmjbrJ6kR/TOBSr2wILZ
vY+H5pnHqRJ9zfcw74CC1WahYOAUSvlbeA7PgZtqdXesuC8pzWVWAh0I3NVq6SfMDAZR/VoJcrjL
TfdNOfFamlPV4NgL7YlH7Fv7gtP4UYCwpN+xZg5i67JKaCXvZZOp0Tr9Nn3GvzmK4ch96a/psRH2
0p6+H6ZS2WWN9El3xUzm8jukDLd6aTZFZYeGJbStVO0UIANu2hj4BOdM8JdQ8Od2y42AmUieVjte
8NUjMMTMlc9AosX7M/yLwqPTjVfKzK+3467XF+Wm2ohjI8NCxPJv1BM3DI2PDPK2ol1VcxU5swsG
1MG9rmsplpZeNVSh5uUq5KaLlgvcYJ7MhRl5FrOEfrop5P2essB05JiUmnQcsZi4K++QzrX9p7mf
sWJKHG/pTmrZiXWCaLGHgO1kQ4Keq5jFc376zpNk0SiGJvlQiIAnj1fXo0DvFVJCpfSs72oA8ki/
tESmbX9poSH+oyGmX4R8qw8AvQXTo7aoOTuZPmB3IptozDrsJCOIIPgH9+BLMIGwBzq2tONiU7MM
k7uRazraSmlz/ZuSl6hKpekw+jpkmBwhLvDmFfBL+FFSX3FACViKZW5KypbHGpDZfTHGr1fhfOjU
xgWkoBu8Hy4p5jhOR8wADhFl/yvvkB/yZQrR5BaKCMSfmQg4W3pL3jj10qKNvPmurXeH+rUznedF
vfOcRxUsmdwbMp60zdhu+QlrwauaWYYp271beCLp4HgM8VSESnbuG11Hb+PNW0dSKEz1wmUizYr2
wHRTsb9oqZDGLbBsUryMgvy9yqUb3A9W6PA6GWvRI1jzeFxQlM2ZvTHUBm8VMVCK+evYYrYk4ieu
QI+DdQCd4TNTFxMdfhFNfiopLrjRVw0QRBUQyHkR8jysKoqq0R3XA13TYLU8JRZJI+ZGBgBtdIog
dTFdOK2jyG6NBQDpWT8mMXKbcJXfsrQPC+/p/e/QLjRGKOnbNelomal0UvSOoOHsayR5HZvh7dNG
Me0BEKgKJPqefjMPJ09hrbonr9E7yMeNSRzjXZ+ZoSiv/EfG4QC/gUkpf1bzK9Ek4FKW+WRsPsET
B+QBnagL9UlIk2Af6xMLKvZLrpI6IRUlmXS+pZ3ZxPBZhH3B+SBQ9fTvRgy9Rlc+XH4GinptYHMK
5iV2LL0Enq46foKJRodzxAbMGhyAGqOC6zcZENWZEZ6inWkzKR2H8wVJt9BKydxR1DPBRySiGLxE
HWm8p1NCnjC7AYBz2AFc8hXIEaK/D6obrucrJ5gfV0bXVr13DDsuWSU9EROFVCFjoSJtkJ+6WObu
1rImjWXLbdVeYQwadsiXfURyiddbcu5ZsJWorQ83Zj7ig7c3Y/oek29TrK3rbq4QHycfDBCNNt1X
2J4/88F2tNx6CLK27UOrRRgtVvcWhY5+zzg1dAMN4qzO3tsVAJTuxtWVu2t/GJ9sp3MfDwpcNisb
V4sFLkWZ01lPaMv+1fEYDv+TZVT7XGVGjUga3Emk6RMq9BAJyOZoZtfLCShxIVBxiaL+6UbDAmyc
fGjbY7QeO50+iHfjcw0vXS7Oq7qTPXr+4iGEM1+iXXIy44jHGYPSgnu9Blu2veqR6vjWhzoflYTG
fc0qwPp6cWpEaG/Vg7d2DX4+FhwBKmY9N3NgAYTrzraRDt0UGnwLW99wUCUhaydPLCoRXgrEs0P9
RkWTC1UA0TzfEEurX1JDqpvBmoT9n+P7ujeDHAKwHB9wq2b2lBw7GAyj41EV99CSc2BkFnmIOsXy
/aRC/xWLKLLLlFizlWe3+gofAKWFzOgP1k2bt0vx4HkwCABRMsaJ1CoUTNjFIFL/w6eFUqI9PdTt
bbfHuPUFjHDh9361AGeKm3a3oNoGCtujZ1X7vObMXi5Uh8iAcfwvM6dGeJ8+Vwx6mgoCi9riAxU9
tpiDuIGUtb2HEZ14kwA1G2fEC+iijor0bmVuYzg9AdGvh8e1MdutPLasFb/g9dB6kDKwD9m44JCr
+NfIUMQQXrLg5YU/0EKLQeyjrJGuyaQ4r+CqRCVUgSNKDac8Vg9AqHG7gvg93QEf5oMc9PqbhQzb
tW84EcqrBfAP639LIf0rZ2702g8ze+G8iVIr3uAAlYOZC43cGyIeACAh9TfUlQwRvloBeD18CsXE
RX6dTXqX2cOhOgQ5bsJ2iBv7wec6bhnFJZTVUVBjq+sRNXTshFF1BBgULmcPIKtC3mu0X+7+ROc/
QNPvTWSOsh6NbK4Zc+1R59MqLGiIpnMEBKaHxDUjNxB2RDflhbr9KTDK+byfqI+0tRvSGvKsHp6E
PQ10UhdD8P/Msvmj7QBc+TijNYt8wUAv2+Eq80efu+2JtLmanRwu/NYEXTyU8TblOzoEb8tlPIn6
haFbP1xLOUAP3ccZZZtOTTrdOpm77bwx7xb//QERdRIXbB+xV4RP1q92mW4nJX2u2ENwqjaBu+Y4
Vn88LT9QBRCWDpQhwRxvOXvyASVPshXHvoCEmHTPUesjjPdqcXDJB1B98ydFlJpnUhyPFq+LhLfG
shf0eOcBVonaFUSgMFPLs88D5F8OkcoVjM+o52k6qNNRtS1RcUGLvgcCn9h0WMuH9bJl6tcSCr1/
655fXL/VPGVwgj9hZH5mAhzrYb1UxUSHY4fSEl/XKtjvsQ+zkY6+TDIS2SZ6qf5kWr1jJfu4+9TC
MsXlVkVLnUVD6OE6uqkhT0Umd2ddHLqZYFnTtTiFKQ51awK6FjRBsbc6Fg/dtTqgW+86A8vZJhk/
Jc7Jxmko18SwtCuaYEnpnsPc0DHidURtXFT7WvSir/DXy0c6S5OQBpf60wKmNk630C/5kDKq4JWb
DkBbD+m0nu/FRG6rO7v0sh6OlNBSWTnFfM2sXgzWoPmecIh8+cZcwNwVkyy+JzADpfPYBwNaCMgJ
DGktem9bm0mWPkt5Px9q1ToqOsYTvGJI7ktsM2Uyb2zvY0hxI5at6PHiyFnMl5lD455K8KChpBsm
+eqGuWZjbMGGzUs+aJkiA7NWu6R8LAvXIBKt5RZOSXrjLJWcWGpueNZpImYrurWuU8q3LdSjbLHM
lu6yZT7Ji7/1/nb9H83Jlv7cgMk+8xwOBfMexgmNJhBbR+rTA4EdgxL92rfPbxBmMbWBjVf/6QFP
tGyPmDfzFqa1SHyJFiLptxRKMosYZDSJ6PkzBacegosK3xB2055jpNF/F/lN0SXYKO3TjxIn2bPJ
rC6HAblmGS9CWhJ8ljqSR13Qu9QratXf0s38AZZ437soSk69JP9h2YJO4V8j8D3EX/qgDBToQ9rK
vSE5K6/lVVUAXsD/m44fiUFyraiY0sCoslabsplaXfPEqpPKY2UU+Nu0CgWTOx6d05chrxCM2bzv
rNJWyuWmMfFYzn6XrSxIS+B8Cr3OCOqr6S1K3WMcSpzzHNPuujwqWo9FntnGWAP8L8ApqIcR/HBN
uZiB/4eprJWb2HkVgqCvxba0fzzF37OmqGmDozPGzFocjwKyUxqwT9bZg+WB7r1eVioijImesv53
VrL4pzZE2eGYuyd4zpn1KasAIDfEsp7HW7hkNwintU13UA7dsJPbj5g34m1/1gaKnOlxNdy+SKjw
WAH7a36rveYQXQCadMaPFMgDeANe6OhfV4xdtmtALDktRdrFCEgppH+egxoNqWftExV39a6lIL/L
Q+Y8kSgXwPNKznXc6wdFdonBtngrpAZSGz4IStHoE7nBp+U6AP6MqrmSrQXyT+S4thEn9OouQGrM
j+W5QuLGoxiwqdqA6wJC/txfcYa2+fqokpejUuowKueahX1iY5Wr63jDCBDlFS4xrYf5LvghFFPz
y7zPuuP2ESK4dTboXieF+GCS1iJblbMxl1yclDUN7Vs9wO1IymMKmdtKv9ZKaag+lYvSUZJsVdDt
JwCStW7yj2SjTfX0U5+LGLWH3u487ahUZXBBEpNtjs//CtsHvQeFYK/3JD7Z+/xqYBJ87d6otA0W
dfgYabxnJj9ItTd6uPGE1gTA05Mnjsis30wKpbG23nO75h6uK+USf2hxZTtQrTe23TOxXmAr04l9
ChW22pvWpmBDxnLAYRljU2tqkCGrLNIttUPZkjXTrsARgjfN6gU0+tLGyCk3P3jvXZTdAtALAqTW
lTfgFuF7BdVd9oiLPbBZ+Ps7jkgjDhYfRMIjs/EaOa/Ek5feGadllIWD+BU/NQfl8/oj2Prf09C6
sIv53IKdSd8QlbLCAbzYknyxkdZMBufuId3XV/Xk3N+xnHih9sS0G9OQaxHZdziGRLQHn0JSyujW
k2LiFmrWqa6uT61h7+ZHMRUzvWkV22PIIdc3LlSUZpCZi4hQrq8iWtlrTsiZDSPxAQBJzf/u2G40
OYK6iCIlYqKBQmuSWe+JZ4vxHGE2FG+2E2lzm4oZlWClXbJR/eUIoW/8rGTD7cVSRJSaOIpvC56+
Wnx/XBBCyTfE7yxAUKcgQdHAVF7YLq3Rg8Jj9qoYG6HrHjq3aA4/N2wfQxVVwpJ64eZhySZrgQa0
3e0/bcUWMF3m9qCElkmdiqHU622SvoL/OOoFhLe2IHJEIZHrILviecE7mEMdGR1QcFkPRIqdy8qM
KI5jJNR6Iz5Rhz3Z0Y7ylaPLN1UVbwBBFXvWy9C9WFCbBg7kPHRe41QWtd1neScqeD+yfeTBw+Ax
TnbgZG/V+CNngEMNFwpYCRhqskd0gFmzagYvn8iHkJk5qWd3dRF62KpmzBK5m0WmXu5kYtgri2qT
Dwvql+suf49vxr5PBtqxIW2ioBNYyQ1vPpHGOk0w2KJJ/H1/nX5ySf1JZFfFfTHbJT63qDFkXE5o
30uobNcyzbgvPYER51IM3ohHwA3j8GJJtX9Vb+8Xn9gpL2oJlz4zj/batKbDS2WCH+6R7h2c/XEl
ou7MIiK3qcEUzqb434D4NYxuN+pmthrOC6cqo3a7PRt3rN1G4SwpW0/XGV/WngodGcO50Z3a1S4S
QFerhfthNOk4qSFdYOmq0Vu/+74jttyaoOI1BUKFGxo1p3NGlrVGDLJ3wq7HZ9T7OXJZCL5o8xC5
XBkmBAqJdmZu8zfaF0Aq6uT5J56+W6PnFIE5eYvfPlig7x01xIXJPPoDxdoeyjO7GMHKT8zO9g5V
/JXoXvCC4iw98Dx0TnUJBjPnvck9uV8Xlif46pAdLRFF7OgP27Zzw6r3vcbTdRD3T7Mz03pt45nL
aKme3LeMXz0jaKGdjuQ0mmZqsWRa2hmfC16+2hq4qlAIbi1ZF6RND764+V9sfleyGxJ3M/JE0+RA
c3Hy+LOomrviJ8hZQ2+Qnj1XmVBdPpYIoL59hN9lMtemfLYmglVZXUizKJy4LAk6SYGaZY0Ea8A/
mC2RPJHzajFM0ZcOwQ6gjqAJ3YGtG32Kf5b0tNYLvK8OXzVpO2nOWinxJs4Y6Joqx4MAXGUakDF8
STat1uRPeaJkykCBD4yHuuAUvhNWLx2oxcpkClJ99lCHg+iBmGkTuNXD2qVPluJXUb+H//sSw29P
jfk/66fjimysaPHx0/sPio1YKfNdjMvZuy3WygGb0Ih/h6RePAodNsTBu5c6LU+pwRp4DTqHat7r
7k3NferhwrzJDS1XM9Rikkz/JBBm+rhfIxIMRBsFaAA3vMDHtIocpJNAhXtI3nckyfVjZPs23Lxt
MS7dt2md0WSoFKa21Y+7hXFNnlM3ekbkUkI3c6OZZ5+k1KqpyncnFd9Om8Qn6e/Y3+dcr/sxE4S9
3xrzGf5whol370HgWW2cqdNNXrc4yQX7dIZ/t2ZmCuNKG+IFti7Mwga8Z1c+5ckOUi0dkDUxCXus
rI+YRuTFRn68porT5lcMkHxcEpdsugBCYARTDY8YIWd4n39aNtFNSHzW8R/iYUz1PZ28VQdVk98X
ihREVyek3XWCtw2/sKBGk8d8wRDrvDzKULUcDWwVtzVLBxIR5ASfXTj/koLCgXtCWhj7F+gFsf83
bRHhLb77sjuV9L8plqFkHmOmK8Ahz4AAH2ZL8+L6l14FkbDptJYvjTzwe84nd9Y3ldm5nz7L1UGV
ZYLmZTyGYHn8ENdj7S1FbFXj5ueVJoW/Zk8D/uUCPS5cuKtm4S6Ri2cxexz//bjBNw54H8scueoB
puK0F7MI01mJDGWye6riBxVACoeSiilk9acyX4HlAZEAFa+D77rrlToRCzZuK382T1UhDkWXa98k
NL6DJ04LoVl7PR+p89H+F8DU0SNs7/iCpBSxeeUBmtAABcWrbyju0ixoyIehDUpcC9uXN0GE2k62
gJG1kZZxhh+3QZq+JxzTUVCCm7654vY4fyGyKmX0vmreGthlaRpRLSopu/bs1hSCQBp1PgiQd9rO
sT0DIUHnv4nQJ1Aik9agh/F0NuepGVtLCYdhv6gDFOaaDhn98BV6pMu9W7cZUz6E2LjerZg+RUqy
a7dZm5JP/YXXLYa0KBwepAIvAzftm7vKGjD9UOnsAh3vZ3ljnvhIVhzwfwnzVx7e4y0V3ddF8JSw
70RgKqPfVLsIhvJDAbr+IAtB/cCijIyWJ5PojSXooq6MGi/lE95rIFA90isbqyUB2Gaz1vPUiXnA
SWHEolZsxSbHJawUprLY9Dq9Wjb5qe2j7Zfagqo25Y7LhtTWs7GWWNNyBeimkU45P/Dh5GvoYpZI
1T9z4lRlcs1KKjn7vAnppM/48d28zMWa+35VrYIxEWUkr2jXXF6UK0XNJIzsR1lpPJe6Td8m9GA3
9vvW/NjELmlKC6c8zD+kym90hr4pMdoF0QxWsn/FhlKMK+TOxYVI0/BJhllUHn0X+zEb17+g2p9q
xQKknehO3juOijC/uJln5HiiJREz54iXATfqRpUGtMkYQzI1S3+uFubiHFqBbRiqHNeQltq2kvsZ
3xv4w2Z9qeQbMM16y3idslaCXu0Zdt8Cz70CTM2MBH2bzmK+b6dPStfQs9espDzAMzgmu7FqHR1t
8WKJ7fE9rOscjbBWTAK1LWcOUDqVREzRD5t7gonixHWf+SlCPo6NtbjW2xoxjBGxQWElD3/e26cd
y1F9FC5p1KZZXCiTULsCRqnyevOyggT3WhsPgszOc17E1+2Na7I+Xq/tmsdgtbrHbCHZMzfboUJR
ddep4SUK//LfcHW8gkEPWf0CpJqZLKWPKFkotvx9wWusnsogAlUtDEMvYyQhvxTpyd7kESXPlrm3
sEBxx0doyRc2tRkSkBbOK23qK1fzFNblo//XrpZ801V/49/rGOdoy99uHfxfkJuPIHn3SJcym6GR
mhxWS9My248TTN1s0DGOgz2bHzSSLX13t7LNw08e69GP7Vb2z6LvcW6xcwOJr8QSLnodAWUdSJCi
oxgaWQfsZlDxWYLM/pMW4UfY14alzqpf9i/Pto4OPMnav1TJ61EJTseuPxlQNvmr/vpCjn38qNu8
9eU5j1TYUutrZYI4AncXWsOLW4oG1m81VpTGh/0znZIoiYhtrOQwUGWeFpfdKbc+Sb+EMsoxAjiG
V1+CfINvXCSOBrEb4r843TS283G37KbeAMztZRiTUGNWAIP8aBuTiXrLkbv0TsBpbvl1DGrnZRs9
lrDzBLVvrIufveAQVtdTJXl45uxhhfM7EFagENvHl+y29Xh/WalE/aYhlH7pBi+KvW6/SgqeEsgv
+NjfjprxonDk1dC6R+GupJumZKOFfHSTUNL1TtVCi0f1xaSjo5uPMaojyCbu753096tXrSDf9d7U
9xcQowZ8GTLwOq3C4VrXpcKKxhWW3Vcl7emnglKy1KWuBewUEzI4FlEi7r1Kk5AOZw1VAU9OUxVw
YbVZMzsER9hzyH/aqoe9iOW5uIBUy0ehw56EOap/AeeAD6CJ4k5XVi4mP6hAFAC8XFQnUiQ1j22w
i6EbdDuBc3n9hNgM07WnmPp7FPTPzGaQZ2+RAzI5xWzIzIqBU+BUWXxf7y5Y5eIegPurGA4mhZoB
/QwR3UNsMIW/foTsfeF3Axs54n1FwwIBoVWrVRD/uQriBgQT8YCRAPVuJm3kS9i21l85ub936umm
kCe/8JdnZkdEy+ZGKNC/5jdMeugNpSKScteZHX3MQMD0cPmaYWJfcd3E3QqvPyUeS9owA5w29pXL
k3omQBLe76+4PUs3TsvXg43Jt5KfNbTnwVK/PNQ3ZV3ZvsLzF/HCWAO+vhcIKENTlmo/tTgZEb0x
t/59A+ad7z5rUp2XM+tU7W4q0SAd0rj97FYYxUIyBc/FStKwnhsNCEqy2f32NKi+RKav5uURCRFJ
4u5u+lG3Tsk2JVOvF2OeBOGyF5V0YoBLl09v8T6ideeeGMUyxyWicyk9zNXaAxMnRMmQ0FSotRZR
H8NqhnjqICT81kk173HUdtNMkeSqifGzOoSf7RjtkDJfgFfiLoW30FanMdkX5yQ4vb4ZGtytTDeh
93EnnO0E/lTabr03R3ygqGFPAqWg3VpbEtJ7X3BLlUlUwXHoBpGGa99ntT0zaTTxhUmi4UXKblCL
MOvpBJFPAXuztpNy1gP+WN6oe+8wrUB+dRHbAUba0JLVY50rtbMeFptxzTwyIRl45Z3ADesrGauc
uIxW2g1DVNunn84Npw3qLsbENRbsFTe9pp/DWIEMezY37Q6bIhyfF7UNuXRvnYJ+gyZt2UqJ09mF
9w9SxPj0I/125DyZOLE6gfHTl/PHNNS2Y12jLQ9tm+xSuY834h8fvO3IP3BriyLQOCfqQTfhs7Ur
3Oe+RvOYUZU5W39aGRe2g7xhouSsTmxQQDL13ItnYWDiA1EMze/uz7RjFk4uRhZqhTvyPHM8fcOO
9tegWPoEFt6hX5L11EKkyoBURkIJQFlKgc6qwsB3i/aG8dIpHadxkPUrkY4yGhCiYFiZDhyLcKgd
COtFgXGuCSF58J2mLITc2sbhL6BPdxVf7MQJyFmdSA02RLdhKH4wjmEse20o4ZJD+pkPc9hoinLU
aH4FdYY2sMDVtXSDaXmBQpcJoDpu6kTzHp8mKrGCo6W6jQfyL0cA/cJPAeIjLemFGhNP4ZtHbmk2
cN1Uumcd2CChJl7gA0r8I+Tu3J6CuHP+b/7dikOM3842j+AfM1yMVjUoF+WeDC+oRoEq2LqhXYKh
ZBjNyLt9Ci2/wDw17FXYkR5w5F0SEqzfRVqsAIJ9cnQCpo30KwrBAlVeVJOxfuvSG9yVT0GCl4s3
ICdZidYDqOrQTbGVSbkIlNvOmBk7aul4iRhmXEhTa5aGmksnRx3mBhRInGyMDYDeXSwZVoZSBVBL
bgds1lV81icRNzlnHokX1p7wFs0uv9GwubiuG937sGRDsMhZaWV5ZsXS1LR2tJSIV7x7UgdTtNLq
jGYWJ1B9CzRmsQnOJCGdpn9SjAculSivrtGTDhQLnXRclAY8/tETusHw99gb9hiNL2wT2aKTgFDX
CiGRBsYp5kVaGJ2zFLV5YwvHCjNXfWJ3jIDbleLbMpdrw/Ci5ssh3LqUAT2cKF9LYKlm2/xlLcoJ
M6nEldDQzMbyyACG3aUA10XjgSDw0TO6WMY2MuY0i0V5l8ixWthKvTG2Qc+TaB540Gw6aiqDZ+Px
1ONeea+uYbsR/vRaNSIZHj8Dq9ze4ArLvo4p+LhXJdqySrQPAFWZ2qx6qXOQkaMqSRPJSeq52oSL
//iPXa5VDzxJo/kf4Ydv6b+57oGBJoVsQubf6MfTJo+uTDHd2Oza9wE1oTx2vLI9sDnAFB8IL2fQ
dQWQzb42S55cEXYiuOaVVV0HY65TVsSbXFtS7xvlx+wxSgYGUm7z8O8P4wulaibmsudBhNBL+/xM
g8K6Sw2RWgACLFy1rz/eV9IfEVUSAzlEL7nU7Ci8wH5C5IctpfKTBg3dWcWsHMUUnkRltHr154Iq
Ptx33jQ3mNKth3sXV1Pz0hd8ObAZoU6ddyZX+iaHufAfTUpYjTrYuT0+svwm0+zxq07yqiJrvgql
E/Ex0IBKuvSXyYYas21I8KLVf4esqLy1qLbvMAnDKnhpAcunE0/XOKm5x+TI7RCo+IvohzXVkCN4
/0avSme0wVT01+D3wbaiRCXvHTOkq48q0KAm2+OBReMQHzBtmwEBvOfL/cDi6uIW1v0JTRhswKD0
eBqFO05odfeUG63ED29GoKPplvdXIAshqOsdG/vQH1wY126HPEiUHFzT/L8NdxpISKCU67XWONM5
+3ie3DNu3vrdDCnJLmlvRfqCkf8oipXFdwOW0EkVAE9eh8yiQN1sBRA9mWqTk118H7db4Qh9/fC0
ZPrhnjNOufBI/IFGBM+nVq9qPuUv6D3fEDEqzuVvzjYa7ZuhKQ9pONsXhKTD9flfrEQrpfSnOEUK
QJ98i4rI2OfDfvzB5d9aRK6ngVOQ3R5nDN2XCNDtXvzKhkulDXsMignMPOqHEMMP/Cvn0R0DTJTN
lGachvKVETaIrYDFyWAgWYyFeE6G0wNxvcblo31gylOjU4aWHW99q+Fjw+RyPNc8dFXb6PVybMif
0WbK/ELgR8B4E+H4SM3KdVHgXRfL/h1BvRf9rl4boMdf7nyO4fcp05Dq8FJ0pBo43Tva/KNkteNP
MKnVrQQ4X5iVZ17vPEe6D363vU2C5Nv3mBs2foo+lVw25JbRfwFMLr5G7sgumkAWSXziP7N0tXH2
Gn45yW9K29gC6evhW0KX6dFhVADraaSbFhOD77aKEmWabmNzL0k1rL7c6yrTR3K6bEKj3omPgs+Y
oVLU4XM3N7KRbgsoJpUBUVZX0YMGuY11XV8KG+av4qeVnpR5u52pUfMynZn2blOOlyeDihYAjPB6
QMz+ktByPtmYuXS5q53zQDtSNHIFj3rZ81tgOSY4uj+K8xfo0xzLz2uQJ1fjk3/qyw6Y5ukO3k/V
1yGJh/T96EZYR4x/9tBWTHPu5p5NoM4pGLkqReMBES+aJmiGTUJ7PZgrFZiSmpaHxmq/KD7zeFJm
lZjGmKIU03YboWhIShIkQRrIzDwb2123KeTRu5+mkfxMKH0LFAdLYMUaHbZEAqEFWdfyQRlPsg1P
zlU5TiCDC8F0TdaQoiLEqLvcIiDS3zjGcaSq57pOg4JXyVpjg79OUU3m+Rv7H852PJPRv0HW3eTh
IQc1N22r9A99eoVytkwKHPDtMvCYc9Ja4pMysxmz7KycLLvg7AsG8b4gG3tDV948LRDd79De8Td1
Saj18DkB9xvGlI6k/K1DFiDaZR5tR6smGF8AZWG+df3ba9uMpE0k0gTxfYxERENGRLBNeoCkE78b
xb9lE0MuqSb+IhVz18+cNEkdh0fcDRBbAXALAn9bfm5/E3/1iMn6o7G8yDfOfqHDHAECQm/+ZyHy
M8i17+rbdfOApU9BRNutR/oHMw+QIazgMgGw577dB92W455GBCQp8xmtKddXvGtmUIEuvRNof0NC
YASg8WL1vr/yMcCG9Y4QPirP9quD52bSs5/qVrloqFAOybW/+0n3PAWLi2VnlbWEsJHchp15BMNs
jAxFnCDPs2o3GsoXkYjpWbjNDBmQJ0M18Z2Tha+N0aWfNNhM5ec2OUeyZr2zvgQ+5N9RDAzi6I6s
HMkxEaa67GQlVJ9yl/qKM6cIQGGa/n3AtzcRYyFvmMMv+medQShMM0Pem6UKSk7ls+478gxIpLJL
dnwfARZMJErjiqYOapj+bpzUfasy2AUg5d0OtLaH1FFKQbSShJHqby7WgVkrNC0XkX08Mh7l/68t
PwZIws/13NkoFn5KBarl2sS8nauPbbFOTUDvNNKi65DiKwyw6G16skvc5HN8XAakumcQV11eOQoR
xn8EnW0bRkkQcAObxSonF+znMSIdbqC3EGf/pblHM/dsJgD2bsDpz349LBcwihYRbwSAa1+EcRAl
2U4MZYfFTNWBb8Lxm010/H/NVTBxNNUe6g76OEAGyl8/K1RzOlFEpPGOCzvmgSjtGuhczw41cCiG
cCNxfYEeA+ZykQ9S/rWn8eCcCiadCnVpnN/v1mgLAEJrhG1rKEi8R2xSARnEkqN9cnCYBAAm4mIL
FYjGSd4bO4ufdDXzXW9yKJdC6/lRDWlc+mKWVJ/QeQaaOePBr9NWZp2PNFdqCMnNZdWuqApV8Pq8
fUnQ9o4bmMR7rOCMORCNqNwiayIc7N30f21BTORePuRpd7AbKMquBA95Lj1QCoO+hx1LKtkMAjhv
CV6XAei6NjAG4uJOnv0m7t6ZpPdGwJr3aTtextICetuoWHrCtuf6aLE/O4eoylPRucld5cv0MUV+
hXW9Jtpbe6dEjwJ4pl82X3oh0Eiy1bvj5QweW9KoeFzxfWKLjyp6y05utNPtqkANK4RueNvhEbwg
vu8E3Jk0X0WkR5ZsP/BIWezHYJejj9UbMqY++g1Tm7fJ6E93PP57NrogWvgy1atJbjl74z42QK8Q
TT2o6lZ6qhASx3bFC0+MZNtRUN1uILCoF1R3bTAbddsERqjufa+JANHpAdqvj/6A/DeUOzoIk9kf
NaeRbmKK705Qba9P19vT0LRMQN4W1VdzEu1fkvu9eoM8rRdkpIpBeCwhnITNdVktjLlpQuzCxujK
ilS6epCcKqQycABzYQu7qYa8tgcyHic063khLaXlduVMNBhVL5yGb9x2vWh17UwBlqpl4l6UMly/
Sk7DsQMfURwhtVLMmx5FCn+pm++mU/EPnR3QxxBc+6X7XUTGV/+abkSQjZaaO3HibcZ/TPldZwlX
wSAjnW3V8TKHqQVBWVJsBHfK7T4cWIUivjNew3whpSCSQAjsHk3p2cvRxVv6tTzWkGmvpM/QY/r8
WJ+gUyw1QO5wFLUWQTFQSRMwBcjlVzDM2JwkMNfeuITEYL2gsp3LQAKQetVvACE2gXHQIswmU4Vp
Fbds8xVDhqOSHKhCWUgjgXDd8vhhFXUzHQqsTiJxq9KaAJZwjXn7zdCLrOGr7WTyFsVrPsz4z6o9
zZVgTv/TnBu84WrueZfjQ8I48yOx3py9n9in9YvdKuSUY/Bk2ihtszkwspGS1yqSlR5H2YA5MlC+
tA2vs8qgUbxaTDMrZW20Cc42vmPaJy5D3L0Wl+mhE9y8X6jI3wFuYrbdBJqaUETAFO+Ef39yY8rC
pHaicjSuxgYrkvcBDtCNVGvM1xlwfLAtx6aS/FhVpwRhE2oxMpPSXIvcko4+cri3ZtZg0sdzusUV
d45oWmWHEDkWw/JCCHyqwiLU39qQWNJ1kVdlGsQv8bZxH/WguITzKPkE4X/KBKUPqCttmdV7j/xi
QR2yR/Nlxrs2VOr7ONtG6pnEwlZunbhF0aPMGliQhM+VISCWT0BcVcvUwgWuV7rPigN62uuGWrAh
rtnimShyE8vXqIFQF1CgVsoDfN+VVWkr7PRY4ohNCWSj0VXTB70xtl+k9zEjO4aTJjeJNd8VWXA3
mG98pzNCFHOvivc7Ojv/bNraXXJ3FsJHnc2gCg/HfnxxcMUvwu/8oWj/LVrNbvk6coWDE5cl1nA7
UNltt6ROT6dwPamfb7EcXMMOADCIXcCV9yrN9IJIvJdn+8l9AMdkGXUOK+ZrkF42FH9LG+C/6gcG
iF15r9KmRyDn14Y4h/A5stB9D0QOcV0Z9u9JLKZDiLgnA0kTk1Plo3GuYuE9XrHGn9nSFlB7uj2W
/RAB+Jq6f0Uf2C7oM13kiOiG9NDYYY6nPb01SHizWI5DeVoapi1ds+/5Byxplq1u8sJ2GE6Cr8GR
8QChFEBkWxrIebiD2hIIpB5eH+nyYyE9Dbar1FakiPBcvdJycrhguBEjTCxArNV1EreAE4xmKP5v
otGXbRIJ2CLOeXfOcroIeVIu1TEdOYbWiaEfmGKFkXpkvBomkL8FdF5Aerz70YCDN/icib1UVtxX
TAPcPH9prVY9VZzrYV+NdV4tlcsfoG2QpFq9NS+n5lYE/V58a6uG6eB7AM9ZUugxCNgN6Mif7ZmJ
O59ZrH9c3s50Gl+5UR9bNf5JNUXopt2YMnIliFCS+vpwRiZ59YrSKOGUUiUSNiJkmlE8VPy3Ie9s
+f/RxJKdagU6CaAd+VrF+aVbeXGryCiCQG9pfm4u1HWCIGHs1IqlDvALxgtrbrdKHzLiPv7lJb6J
aIo99uoT0ioowGnqe6P+XHa+hCsjv3AmsSPwSw4CqF4WAd1/n3UQBQXxlPsTuBq1dNGPkifeOnub
4EWf7YlRqJbdXnwgnr2YwCYgvDwxNPEBwiTzzBYLMIznTHhHbdZMkh0dZ0E24rF628+hqBXI/LHW
FIUcq10s53FzT7PocV1DCff8paILHnkvVXD3YHPHHAAm5avI69Qwy/E1WX/4CHlUAn4YwA8L6VtB
cOK8VoY5XELHyo30eDs5Pk/UMTAGIy2z4jMBr1Y4mk/Mlkpbhs9EUNZi0delZb54DUcqAL5DnXKk
hsyHy400uUl6qw1O/3EKVUvhYW2O/AxlnOh5bdgA1Cd0xUtmdW5Rhw51rF4nRQSbdEAh38G7je6b
B8zNlRb37fITm5acFYOUVUOYP4ILV9XH4Op8NPn0oA46KP8I329WszzA+hIbkIPU0hZdiBR6qztw
/sq0rUqAUHL2WwfQBgAKrNbqLuCDpkTe4n43fYHTbW/3FXDD9xZQxHfyB5f/GMk2GJcDZt2aiC7K
fGrp2EFf8OQx7B1t/OIuTYYQ+bINiqJHrt3AdU9myrdiMebToZ6EoV3VU+8G6OJPJUTJfeUTXQZ7
W/or5M7eleW0SJcFZ88V0VcR76L73iZv+0iuqdUiJKfLRTnIJC+oR/rLA0nI1d4I8UQW3upgKBk2
pLiraMShHPdOiXhanwSLO3J0P/kkKFg84V4huclukquLmTLjF/8Ejp7bGJwszIYf2LzF0mfSu2+F
va2rFpyqvBf8Lrn4WTvpXoUdVMgixHYkbM9KtXUToM7gQ0QgF8QFQh47JrwZwLqG2IHWtLCOim/W
afyl7kvVdZ42a10XvNKGlT5FnUKy6tbqebTMEE+i9vRNr0n10LBXLmKV3Qgt/ZiCSqh3SR8YLxY/
s2Wes4+dnWvRHoN6QTc8cOOzBrhYNNh5EACqqB0YA2eF+zleoFfhHpO3MONzPMrSnoFDoZZ/1vzy
IdbPt5i02ChrTchkQ/yZuKDhpSugcatY+Wy0YA+t015CHnMdKjZ1HlRqHr7ki5AjhKJ6Ud4t1Ugm
NdarYGLHqYZMcd8fwPpMlovVAiK4rl3xOKkjLoyC5h5naAIr9sV1tTmAb2g4m52zklNC7hV+tCK0
I0BpcD8La0wS9KGcrHx3/ry1YP6KbZnXt+F2O8WKoHJYUTCD37SzhV8ngMIo9bqB7DFy6Gs1x4/f
lW+nzs0BXivxetjfIQ+rqxMZ90kE7gKVZ1Pw5Qbs25EBh4C76hPFtSQqJC1NtaZWLQduslwfIec/
JOoBeuDicFXB0UMXPHAZcTG3kXe5sNAMaICaspaaOJxPhJgy7M+szDBOQ3eUlGamCMPrT08UoSN7
WG7yn+4+0xibCZoY+A5cTWzqe0lAjym/qM5lAsYwQDmRsUh4azkUi2199+F+/Ew0PRQgTm7NpmYv
avRcrKw1pAZTXcKs6ReO7xg9tqExWDX9vaQrSS639ibqCSadcCftjsV0dCSgB2Zd48MSYX7QlEcv
YG49GxrH1PpzFKWjhZMrWRWILTBN3eYbVouJkm4xBEaaseqy1xjU7AkFcqUNrWDz9ncnftmdRif4
07OGUjtX/rc0G1kTiD4iVdfEwcyMhKffkNm1fBAfBD8j7OIdRMVUYBRkPl1kSSplM7fBi37YsSgu
CawKsqnJzJ3Wm7fzYWGCRT65+cUzJsC465QsDqsN537Q306ECJDTpkB0SiasdWmPGmtgytug0TbE
hNQ51YvLvDE0/FWbwBFTSnXmN95bDjlzHU6UHgRL+pv/pjdtkcmo29qpKpCqpSLNDTQHAdX75Lvr
SM3i9N4crdRb+SXQ7eHzbGoKMuXBcCmoL781OglnNf3ehQd6VBuv2rwOfTZ/fPtfBqRrKEItnNt8
Ab1awFNY0Am73myHIyxrZ79QXVQKcb5YJLSjcR/QjhL4HaoPHLuk50naYNqh011kQuvrsLDX4maA
D1vBa25HyNaUMQ6vnPoxlF7SZx7hf+XoyKHm4YqkrDXT4DAK5nVAelz23W2/jbi06L0QwXpQvuwy
Wv+QCefqly03Ym6980d+x6dRuuhxigqIe9YIysU26RmznVdyLuVsHUyPOJ78T9r0YTHWZ/+a9iq6
ae0zh/XXE18dMM8TEJwDb47D5qIeiHmxRmi4FDNxtXicYjHTwhRjcDB8pc1VwtIR1cVEAK3dHrwh
rh5EWeOvN5tEnrVGBRZSFcybxYYbQoSWtWa9ATkJ9xFgIHFlzx1neRWXR93bfH42JDIynqACWNbe
ZWXMRoUhVK9EorDfMnJmYFlJizjOtls6RWhcKodO9I+aq6JmVcokIOaYkD2EP7ROrVA0M5VsISHm
UaeCBsJyfxhrUe6Qu+ftNMthDBZZ8KennTmZ/K1Cm2SqTAB0Ghyy2gti8k2tvKCh5C+FXG/sWgOX
goUi6Cz9RYZDOr+Ff6nqFlLHkNTZLB0bUrk+vLZ0j+lpVouvP7pcMJMuwENRXHZi5UEQk99ZPYpS
SFIEOUqtIK9ICdWBydIixXBaOVIDDC+mk0bdBZ5c+I97NXNPaDG7U/Ttmtc1RRPbgvwF8TnhRE0/
sXqxxrxNur6mynq17jIen/Gj59cjJly8ZoxuOecJN7rFgwMGMK5IBx82Gur/srV/cjHJxpfErGr2
/3p52kny4ge3vloJogAErE++Grj/KRmJL4K0tW4Qx/GcxW6jdh0K8CV+6jojIule5KzAW4krhmkj
OKzf5KS5lphfxoCFnjsWO+Y45cjfMCi36rFZFvxtsDBLu95MmXwtne5JkiYgJb9OVkNRbMiLneee
JhwJybIQ3NVcQZcdmNlt+BMKyYZw621f09N2o44+4+bcpM0EMRzOt+um/hllyH403x7zCS9MQOto
tILEOqG7W6wDzCfns2LI7KvNflhOsLtrm+Wp7Wtj7drATc51+eKQZGBMe5xrCayeNuwfizVEvMAy
3djfvEatWyPWCSbCdKJQTYMMxKZJ8Yj42hzyb702MTA1hMTFUqeQgKhYlXwjMwz1CfY5aUhRxcNi
lXve5kJ3KOyPkQDVUjqXVJ96flpRkYbIUVSYYqGDn5X347Qzsa0yfNCmiyQzUfhVC3xVJO2B8Was
vWqLbxziN+1fhJRAaJpt0OEpjeewPBXdLC+TEGQjaoTGvIf7e+MvdHEeszdFpSvU39PgHKNby0/v
WF9J3PXE+U7Lx5aQxFlDMDsspSYk+KxSy4uoaFlOxLZ9Kzc/9SInhFjrLRZKb5wtz/A0bbX7lETi
9bDnf7vTb2pt+trrmfyLb+3gu+CDxc9CGH5y4Bke94PHto/AVvMmTHSSKkARcjP+wXxu3jkYnP7+
k+c0iOwqblYSYYWWmZq40GHdCbjuqQx1AP4lDsadcfkk+qb7cpG8BShrTMKF+wOILOAwBnvtyz6H
t632CyhkHwnO5ACVkFeoVcaC1ygQ9AFz4nlvkFP3iIB4GzlMrJNHfEYibLIf/n82DrlGtQnqpKug
C86c5RNNB/TAgqCpY++VSs1ItB8oNkPln3R1CltnkSP8GpsBLsiVPpIHXGXoEiuVFm9Wgn1Egqzk
uV3S5mLeuV1YE56nrHQKuOd3euCFzX+2vO0N/mRzGOFG1o9YUpsIGrk4gHO+qH4U5Ph1Oo4M+FPJ
hDSPLYQmVTSrRC7MzqDXHyp2vNuPYYnncWAGx9gaMyTrLmpkq/qWdryN7PYp2lSH4PEWbXz4TscV
oPWGzNoGrA3g80GrtG5Vh+DqHGctEO82fT77D9BkbHdgMGhbmKu+RdzvjY+vyzyS1QD2skG/kPx5
w0HT2t/SRrSog2eWq9VdO1NWI001C0wpzcVgk+7I3chA15pYQN+HbGHZE/I81DJ41F14GsFyt38a
fEI60Pa+09HnhEbU1iJ1YyD0YXWhB7AUvUOVeSoctJ8tFhR7qW8seLZs8Xnx+Xp+d/kzpkJIcjZH
i389vKRIKPfWvn4Ldn0EGUqCQWAOtJ6AirVfGDlC72NyDWsdzKK737zrUs6XmDgWM3hO3EJeZZ3h
fkMNCXQiXMgqUTKgb5NsYh6uQjJXXPegFyOrTUY82Rxg8dW10PwMvv4ie1V39GoTUX6r9QCjDBu2
8ghFlqrIlS8VFacoozd1kMVvq9SiWujonQIh1zyRd//u+hT2vMyQT99pF5CCbp3LVCnrumoNtDOX
xnMqj7UnfXbmw/dV4cw4AFiHwp7tV3hmj7DSHEN8ur2pJmrE6FvUlweTS6vYxLn8cEl5KvZD9qC6
cKPbd8FMVKJ82LmvglWZl7HF3BRfAUlWJyHRTMCdv1yfizfLigIZ9EEDc52CZOqWc+8JSXnkr0O0
fl+Qp4KJqRWIucKKUQwVEIwHL/CpghFovZXybvV4XWgN9MHPyhjoo9kIImQrcS7kkO5NWvLr8N97
J/9fTnjKTJmv5c38X6F7+oMOuiFhOYledRCBt/BilZ++1Eqo0APfYDwoBQoKOr9Dv/CPmMjL4yi/
Cbq8AJSCknJ17f2dO9shno9+NxKvvjNoK+f7ImKs3rjMguRpgOw71vGjwdwtQgubRlY5RuzqNoTI
SIEquslJttfduF3iu72IyVX1a8Bys1C6vC8CetFKrDX7ysDFV3B/QJngxQH3vEmdj9ewmTpMAzqy
1XQKdNJqeKW/EUj5OtyDuV7fSjHmDn/Pi6G1T4MjjGdugs+4jVIkcbocOcfhrg11151XI0vuiGes
z5aP/xhMwiU7nucQsdB23T5i1GMAmGL3c3vOsNNU/3QtRk5fKPjRtuUVgw07Htpmw1gWlTtZ8YHV
EL6riQlUjxP66XMs4ck3quM+WUmc2hgEYZqjH/H5LgkKJOWM7gG8/pyDpBueHp2nFkg8Uyv5WlZ+
FoRt203Qii6IH/WVMU01DYEk4BskCmWh25XHtv6VPVrSwJoHUbVA3YsA2+PRTFujtQjvomOW7u/f
iakfHYamPx4NHQq9yFu4us7m7oltYIO0kwqSFcrNmKy5AsZ+wlYq+4wesPmBIfs0qKpSYrmLtGxe
j/uoAQFaxHLGCPJ/z/IUxglFf+x+kBvy9c65DDpd962hMA8p3j4xtAgG0pp2pgHRc/s9pgYlED73
buhYsgu6uMy1cwRMzFUB41vRdi9TFmz1ulJNwRCZIcKvXoQJnePqo++cSfoZv6X2ULM418IzY+qo
J2A10fs3vfQJ6akmoFNkvMIy+/DCd/Bb3YJTX0zj1KKiMsWTUdWqM9uVO8MlayVPzT152k2zuHRK
MZzqQjAC9yKRKu9bX3FO+sSNw09MXoCTAvnKY7XGfVuTNgx13hBFCyUtDgs1fDHg6Kyarlk8pX9I
HKUTM21hqn3LN7dC+0Ha6aRkYw1/iUIB/UZGcIyEdauewPYiUd+jOye9i0grPiVwXUoGaklPN5xz
UwrKQVkOOA1/PNbleuYEaq4XUlHutdPvj/PzwOveTMQXskmU4blTWIBrApy1bdmzJ4NlYbXykiua
U85ZOdFS8loolTdndts8GgYLhW1OXBGXfa03ksV1oyZ7jfFwaKXv/CTdhNuuCIHfu2EJzroNMlV2
5lKKVmYt99QGQAfMXvi6nUJC5Z/OD+ePwsADGb1VHp6EVjHTVwEdPsB18CLn2Z8K5SR4XolgjSbC
nVc4VuguLiJCvJGNyf7dUTMCOdqMI/ErJ6usF9SIb3UUICtcICw2WojQbkHIkiK1ybDvG/mlrTIE
/kRvtn99f+DS1U64CmFxy2E9fx3gvGYssMY9A12ar0o/0kx8ooA/6SUZaKzfvi2cH4eR1YyAVM92
d79q+vFehGhoKVAIE56cqzm0zt0vcMgtupkKSfAf5FqsQmhZDLCF2YgRAQDFILAZeBYds1XoqWdN
eoC41wQbYxBQcsoVqPFwQSnl+FRUbuNEyelySoyfgdGSQV4nXF7EFwiUcG0XTFfL1+vdLdHIa8HJ
vtLpslNysQLUPz1+XFXixPFbQ6I4BzxL6KQ9VVLvfatwpYr9jyglQy8S5HLbezrH7MPbNwvn2O95
HQwuXYzLQeDEjcI3GlNDDWR4Mb/US7IAWX+KrP+ywCCT2NPXkKKnGsHS3DNrWUjilv6CE8HFVVba
pv2HxAo2Kmzj2aBBdoRZ8G490GlmdwvOTwt0BJcoHS9S3HaxH5dm9C3k2CIbi9JH9PERk2m9e6QK
ZDZjbGqAn0634p/9NKtBE9MtOd5Mga6/+wHgvMpB4jn8Vm2xZvhpKNd+TKM2y00+3ewDu9rkd/Uy
pd0G9laPRdtlzhl2sE/OfohvasRQC9WWFJczcnh196c1eIDwm1w0UWcm85pZBUQZJ7SPDCjJ+oFg
XRr8vcgOQV76v/ffRmE8FwcCJj1giNGPfPHiKqOA9Q5l+a1iEHSzBjjWikvmUHuKRj6ZoBthF1bc
TljBSRscSxa3JtRamb7I8VV+jq3umeQ58VtsEBPYpYFSGkpN8cI1kaHGlDZbZQR5QGunuF82SOMO
rmmJn8FTfLgmkNdpi1JeFW2ZIVuojmVepJYfc9tKxdEiQj5u3yjx2MV8E05n0nYWeBoLOTpPRdJw
47Gomop+z23jKmpy/Md0UARDe2+6c97sbuNjbDyyct1SiBUiEPmf22CTr7KviHjG5B5iiuBXtgTd
JdzU/dGWv1eErUPvFT4DiYSbFePmKv+2/Khk4BQIAqmEzvK7Le3nkF8cT6ZnCa+jTabuudLJ9+Xo
uNtOmDmfEoltQsBVZNJSir+V0dj5zW6TRcDXvYYQ4L4UtrSOG3kpJ5FlkuWpsr82keDIUNa6jDOL
wOc8iS2pZk5p7QoViW/k07tuVf1PLz4sg8WijFcYotm85KmKQ8nXev6j7ax6fzr8DbpZ2i6xbDf8
uAV5RoQZhzCF0UHzBIX+0LD1xwWhDnhu+pjQDgdUEpGCzYEC5tIFXeFh7Fm3CKS4F35BixIDmlgv
MTmXSygOl+ald04u6b1nHB1D9keMyxHsg+wwcar1b2A3hnDTRc1KHhFMOsv+mjDVFkX0Vm0oY91a
CJuvZY38HtsmnD5qdztZ7PgdJZhlqnWe9P5XdIK9szW8RkHjXbpDAWs7HrZc3vrFIaJ4tByGXWwn
KFPpP8HCxlGIQaP1zzqQ3j2OarzulaVRFOXxMws6sEhAygYTIxySRBkdW5BzN7j/DQIj6z5m9ix8
6AyaVhkFVgIpwNk2A6C+N7IsZo7q1n4IXljSuspQrnOfdeKyo4iDs7a9L4FFpXZGUTJk+Gd1DYvk
hWhtnJlgemTMrlmCslIIr/kFnjvE9bQiu4MB6erTXFLUQ0cFGX1wY1zRpJcWwKM3QMhwPls+C8n0
6YKahOajYffzhdULViky5GLQvzxsCBwCB2ik+iBhWHhPhVu5jToIam+7ot4F1LcQ6TW4j9FnuoGu
aWI/NDlaWyZRjZ23w8oPnZ+mpirI6n2wy/o+Ya/7jTzuHLhgCWpqmVwz9KblPhDcJLJT4T+rxePH
RDAmQ/8xEDwfd3uEwTXUDt606J4IUxvzVPlqG6QL1gG9FvklBuWjzW90B69frTBX9hB6wZdpi1U8
KznGfbks1V3HYKIHXPbhFYROHUsA0B4bgLpO3kNY0jG6nrRnLVUiLBl3cgtpwn2rS2AZO18FsqgM
1p1l/IEdCdgvMbA5YX1Gz4hXniSFaQvuu4MXdnYWEsXhR61W/NOXBhF1w4uaRZ8E2i1+0wwboZGD
NVZWCFFMQU6PMAAfs8muAqWie9/laBui/j32pCozgZ9MmqUTYL90h74AdXSGkmOgZ2VibLWqjwsI
h1qKramQ8Ypiji2Up3iAmnQNbyiWxshc3YMql5zQUFPA0eXhuNTkMllb0D62FwHPte9LZUmJLrTV
HPQ8IO7oJqSSMNG3FyylDNoPj3zN+VqT+YpswqFjoP0sU9eI6pKdkPz+D/ZV58P/DolRZXI2IepK
7gjwhkHZ15i47bsyo5UbbP+VvJyoqFs2rn+p7sDn/rUN3wy37ncqzVOkMhmfq4tMDsWIA0cl17Kg
nHZKQo5iXX2/ZSOnGfHuv7krakfnfPpo4fTx9JzNUZV4wOn8IPJQDVTEFoDgkRxyIJkQGd28uOlg
aY74oFph6aH8Z88CyIG8PKlhYAvZyr3mPm3ylBIsdEI+RWpJTtI9EchtSOdIWvBXt3qBv+WHBNQv
dPgWjDTchJ9szoLB8EE3AqRQjAzsqYbEUkKUCW4qD3ltO/YEWiPvy4er69a7/lA8dJJGFdMDC5uR
zxngfJDvQeCZRFeuDTo/L3dpwdpXHRRk+CIrGmWVf3GgTkSUIaM3RSwb3RBeJ8iEaeOEC1K9N+Wb
B9XR1P5GrHdxEHVJDFR6Hu16LHjk0XJzhmdiO6JJUD8iZ8FizLxLsWuEvIOdOIT5ixkM/z89KtcN
ekjqYPpw5abWHxlGZ0USCcOnFG8rT0u7fgxXSfpYmuU2C4+/JjOlSazmUdXqCjP+GFuShsT6l+pa
4ONNc4Sg9FGwcvVVUSiVdlwA8UTCzjz+73AoiV2CUrqOABUPVnXA2nCwXBjPxpZ44xG+zhXtG5gN
jRkLm+y11tYjE8O39S8sUrZa1+kwCATY+hO3l8SAgCVn2XH5iIBiPfNhz1EbhJ9pgJLRvhYDCvef
lBQW0GlgJ4hiaqhFTfvJfT1gPmz+czcxixBSlLTCZnKKR9eqWj3hTyUdNhaHFwh56CEljFgxN5Yd
nxcjBScZHPFmOY3NymsPco14Z0HhXLjrLergnHHCqK4HWuZ6fQSKUEMZi6lpkppv+1ZmSJfLZhBR
PuMHEnlNGHUcOtCTpP8baVjkKEC6xswF8hqC5c1OI+JvidzXdbn4DHgzmUlMLW1HWrbTZh4g+naK
ie/I5NHSSzZj5nVSMBLJ7DICBvRRcfAYJICMMIBXLG1IEUPrjCqOl8Q9thYqUh9DVlqv9ZuHZcZL
iiHx0+4yddM0MY2FjyKYfJ1WC+rRChoS6Ar+3ELmjoTtzA4qmATC/hTAP+bbacbmxZSZDoaJ/jrD
MtqszBrdmfiy6PmcGTTi+F8j9zCjacyPuE0YXWO1npu4Ay7l5WivGSE+wRvFonaIpek8b/mSS1Ir
u6CiOooJ2INeC7dorwTQKm3um1hfgqGUvfOTqC/yxzq+svbElSZfpUFFGDceXO9c30SnuWRTw8J8
gb0/bGDh+noQfTql+ZNjnJd3sT40olqnPNyXtpx0OudWix4Z9MtbNY5HTZMITPxdowR8K5oRA9OT
QNoiPMykpWop8QDhCeImkJxFwskAC3pJINeykCGlinPKPW0m28yGnutAaZQGIkq+MX67qg+1U8MP
MXS8LNjzWWE7f3pvwQcxpKzdBtv56jZTCPxqasNfIbeRLltu/XG2FDTB78Wa3cm4ACc3aJKfYbgx
rPoMqKcVwYERrfJZlMmWh/MUEBYnnH8JwCapwo2xxRNR9f+hXx4SzbUyX7OpZWFoMwVpK3Ju7uVC
Cp2/1IG23Bf0m49uyH6leB+ct5bTaXQmLEO5ruO7JKo12kruHV7qIZ2zGvU+iLzXjx6Q5MYde50b
iLMp57WdCjT7voxEBsQP2OtzdRwrjIxkE+/XCAfbBhGh9fFi7cL9LWknoMrLpTrDaW4HmcQnWBvX
RNPozIowcGDBJs36+9wD54iydNFDW5qLcPG3RgpYNuhuSEV31bGV+4ho83s0nagxFfiKEihfb5Of
/bDaYwOgTh7CkA+OM2oc+ETJIyIo5oqGzpiNvdBbJKWq7Jz7ezAl1qhUf1ePxFzlK1niWfzM1JpU
f4O2xGHoKC1u+SAG/NEViQ/GRFWO7mODvAafztBcq549Q2fpG4xXsAoIt3qGkqEEQgh5H520ocJ5
P0gTaXPgc9/5WkVSPWAgy6gM11TRnEFfYzplrqJCttqUdrEwXA1Yh3LFkZpaN5yEblcQ4L2dzmsM
in4dC7Vcy2+gGGhh9L5Km1So2OMin/SMvdBGi3G/vN9ihBpdZHBBLz+2cZgtx4amwdZRfFmskQ+O
X2JG6FpwX/Oss5Np5q4Aetx+hzp64tB/jQZtbXfg020LPVedTN1fHkmZdfl06hJC/38fXPMDd4ws
CsI2XEkne08yzTAWJiEwWG3YFvROyw+iYcocxYe+N+TnSHmZFvT1Lu4VQ0MkU9A/RpoenZOifckS
x8uzPg4zY/se5c8qmNCEoEPhrdxjY8Hd57NC3GO3pC3hN9b8wEuYTjgCzrPtQ+F1vt6W5z8D5Nmi
KgQT/W3T+9PAs1pOI1H9UfbxZs+7FfVR9AEjA4ZX9dEJO3Ld2xhpIMaJSJBdK/UEeZ49tDh9jpst
fcKXNeLHin0+q/EUUemuzqlO2yt1+6lndY5PZB4/o+ViZ4GTRvHwsBeIYxu2e9eS6Z9sDG6Wg6nR
o9KZd1qHPA9fYmJs/WkL4SMrQKb2RVS0RY1SEgW21giAwqtmTIzmQ3yut97yRUwydUnxkKT1VNMY
3ql+/0qH/PWJtLRj6R6J/8lsUvvun+QCP8fy+YAVZXFSEJazugZbj7ZiHhj/li7c2rpFK22Rurjt
KraoFWClwQw6VRDmeNZEaqT4Q+HA+DpHmt4UKYHL+NQIoI86sM44Uw5AJUFnVzxGliIF/sKSa3mC
QTEeq+VuCLPQWAlwfReYCWI9bGHuJ01kTjBBoTzrCD4mBLI39r5oosRouwmqaU9/eQwjVYCyBiC6
RaqTKVlrvCoKxB/139+ultxfnCvYghxdfLnY7MfpQeAdhlddxTZ1Ilt/pYZI4GYXjBKOfg5MfxY7
WyNVegpcLgIyzq4s2DHnn+j/dYQOZmfI5cTOMI+raqlnHhVB1Ef9/edhO52TSoswTuNMHtM/PaiU
+gAoU/bpdn0eH0UrzCqwqfTbIqp4eBSf3J4gLUkkxqygano9OM1aM2H2x1XyeqF+EvFjizLp+VgU
9G4TZ/89maXU028u3Sn1EjB2h33kkh8AwUzvh3JBrdZmil0teRCY60+hcCG+zmmkYBhLWByhLSfq
ftJU45fniVmUSbcrOsmPz2kv/bWlpkgngLwGUCNmn6MxSkAkXibXjt8TlF/ZcLYlJvg+3nnQjglr
jRTcUXwHXdXItPKCmnfDxntjWl8eCQEcXXGzGWDptDa8KD1enZQcPGhY5an9XZ7c70iMskqcNyaz
LPRoWFsGpEhM/6Qj1j86Yq7ql4KQmwivDzw3ZwZwXkMcuj8eHD766ehBrcEe2JpAWTk+FP/WhHUw
FHtmJ9IieaDkL0DLaVnlHBuV0AJZcne7eGpoG2U42VsazcHioDtriB9EjQnldAFzqw3K0iiY2Byo
vhyCxiSEbIt5zyo/EI4nOryklFo34G3jyAzjryAInCKIH8PrGGPWJ17bqlMI+M8txKf8pXzEIgZK
utZevJ1QSYYdTg7rOM4YmrsR5UCssfQdgay0G0NoaZaVUPzBTnPaxwsdzFxqMkL3sHYyYG6aCGaq
mY+QYcw4xT50mCHKJiN7BLRjRgt8l+bYCe8yhN1KyG2vIG7z31ecJYQiCPql7ZIOVh+NaqhSaWB9
ETIntPjeDBsZgpqlC1FjAyuErw9QEzmyuPpPLEHMkscObJNzDzP+LKQFFm8IYRWObSJpD++uFjfs
AtoKBBmFrcuOMvJEXef+Uk1fFLIP1SHH3L5S+kCeU8Sah6g4YJ0OgzavVzoGCPT7qT1Qt2krFLpb
iBuZUW+E9MtWaicQnXB49PXID17SUubkpr9K+vPFyRCcvnB4OUDXmNLCSJe5QZexuGWL6/+fJP4u
eI5xl4xtwxGSTmHcXas7Ge++SLnOhbAl0QFlfsxQ/8RXxeA2pM/Enwbl32aUNUVu1w22wccSHf/E
8ZOSMkipFGl8RbgGCROiB+6iJdTOhwMqXtRDqFkRHsDSniRo3fFSZdLoMmRpsvUGvobSA/1AOvxn
Ud42cYcwMc0qP6wbEFbzpR1iLzBK8GK9mFbTjd3cvgPrNj5mg1/5apNi8LYTazRf2emMtlsUWtg3
lepGUYb5XbnZ9ptkhIGFkMEvkxPqXR69YuLmX7hxOzdpOv4rt1V8H9a8QueO/oGfQMytq54H2gib
ArQzRw++CcJAA6yHqX40xWAR0yxQnCup5t2zRXRl6O+njY3Mf1i/SxY0MmwW+3YP6LyyWoMTOjKF
OrG/B9w6iXw6BLU7AMamLqc7OKWrpXmdHNvPOLZvUOnKp8OowXXbZ8n6SZd/WuLiI85y3BdhT7s9
vbEMoqtnjCldyBTbO/9gWTHymwfGPzlXuBXiPpwMdGKBt/mXRz002Cf5ka+z3fVUf3YFubBRTRtg
bwy/AqFeLQ6m7A0IKZOj4L0hNeHdf+SmOiccl4g0n757T8zy4AE13zVYFePMXYVMYWIA+pv0LpeL
p6Ievf2P59dm4kUs3MYXG/vxdKJdEbZvl1nhgWqhB2DwIm/V8w6oo9pzYRnxEbWPJpVQQDs1Ddzf
jz5ih952mOK4ogiPZKZdXcnIBdidOmbnOdHYG3zzEA56gNtdyNzGbY5BZcok7fhyTmR0rgfQ0eLe
96DnYjAMjoLLVDdQJieWFq/UOnmQ+mdTgZm6SDbw1mnWhR5A63F4ZkDTzPpKLX8KiYiOFu9PQFss
3Fk/hdDgieR3L8leN7NqD+Zi4snJ+M8sFuWS6qMTHsfWasTR1DxxIMIGamveNo2tWfRQQRcGfR6s
OAoRmP3UAsElGnIyxG6sukntx/UnDcKmQ35a4i07VoVxvZAS6LGmzwlemG9DCuzeEvlFdXtjdwV0
t8FuuJMPhapiDe1e1NpJ0JNbFfz0QbnpLj3JRdUWMN2RBOzDh3JmeeujLSNnm1hTL2HE+IAbi4r8
c5A+Rh0JEZrT7LPQnA5T3wwxXqRMgISScUCKJUqtbJFyJpj4vjTPh0WQZHcdd6Op3nQ4xb4AkDyc
wQQA96F6ut4PG5/XxOmRz5YPbwNW59bsApkkrQuddN2SUtek0Idm8YSvS+xITZ/FizkWV73YQIGz
KOe1Pif+0lVCiU09ljcfbS1jozntH6vAAlDuDzeIjaY1z9FjDb0KCQjRPYiA0J+F62ZsG5Qw2+S4
qNEvSAg9v8oZ21zRDknPPPYqZ0pH9miwOHCOn8ZEO9M5T6uPGRw3bRPsIsNYb+kNrB4yJQjwTZu1
RPxT6IbTkRRSMImgkd+ERcg0jvmtwJYPs49YmNtonZv+3v98T9UtaIATXwP435TRe+8rxKn4Ki0a
JP9EqKV5Ne+nr3psUQRzBDmcZSLBWBDovWb2WfAqaNz39R/VgP7PXN0/kF+seWKZue2K7BQxgngh
k0fhM5XjZ9qCCEIuiADeN/eey71mullYazS/CdusuVLFvyCt04NpuzqfR/eP0E3/8s88ROFjTgr4
tyeiIVzOvwDI1B10rCBXHuR+GF+1p7sIS4jO9jrn+v0BrbwnsSaaSplP8kMiE529x+jNuRt38Sx1
iS6+WSJ+VUQSkX13cu19EZp5UKmalDprZjIQpM2fFSGWqCm9pAWVUrxo11Ebs2vUk5R5J/ar5PXS
bg3qhHttPlCV5LGnU6w0lKRBVrM3KGpIDIZsYCizIwoCLGEb4yFWX88pmP6b7QRRSxfhop/Fuq2O
gySoIfQClUVeP6lY31E2rE5Xv659sf9OHgXVXqsWL476PN7FqS1g/tsy0Q7hBBGli8HVxfizJKzv
7uoK+I67yoHbggFOC12VOKCRO8F2rp3w8C5/mYtOQ33T+L3c9+AiDhjMroRzOLqYs5l/4h+A+qK4
jnmVtjZZUSjZwS6ymDFlfALnCkG3eBi92VO43HsDlm2f0V5MUWJb9USuLiTN6Z8eriHyLJPd5dJz
WH7XeY7JMf8nROlUm1s/AGfnWdC19NVM2c/ChuNLsj81mTB1EtqYuNqKvrYh20aapUCRDks+tRSj
QJ/ecgccPDtkG9MxSiqKDMKv2l95pZzXVW/ze092fqUjmjyOSlChd8Thn4IQo3EVfRhv3g2XGmhR
SsbM6ue3YKsWdo+9AYT/xIOSNY+8yQHnDu7xpmZQkqw1dApTRh33uazi5wfV+4SEHWD2IxS8L4My
mkijYMM/QOpo+/QX4SoFt6v9F9t2PkDRSYdzTAu1klgx9J+yVWU25iucsvwjqsHDPHI4ap8bdLya
JDW8Nxtzkzj4h9RnARpJFWBm1OwPWCavHpx8z0LRv8mMeEMdckWqZ+LZWW6SNelXJdKlIm0R63MJ
L9xyq2Wco3Zw94ts9UG+XSQ2Y5JEwjGaFat4/kjs3sw9SJsvQ0/l3e7kMEO0dBKGEUmIlLvjvgpA
sFrvODPOFCDTm5/r8wFelYqTzP11uQzdrW36loAE0rP7/USieq+1JieOamEU0zPdcNuMmeJPBXP4
2Dh3mXWel4kZrnNs5+mjq5YPdDA6ITcw9X3755Og1AiejRj8ozkE+Pt6VNwBNAEpK/lRao69lFwN
CWEUgPo+mTA4RpSAflNBwHyErvKFVlUgG8ThLEVURa2NUFWWqMhb+UsMFZ9Aj+Y4ASlWefnmVeJ0
c14/nkMw5abL8CjGUQWyDnxd+BO6sXljfXErDn7pEyLn9WSwaGD3+3z0ohUq+gX75VFf9GyQx/Rw
ql/nkCJvFAP1FFLwKIcScaZuDsdraCK5inXVTO2tD4uKnJoaFT8b5FFJ0KPd1JuNap+tPAxd+SdQ
CNV87BjdKhnH0GJbjW1xDxdnUZOJrb4Og7Mm6ZTvHWcpimdJdRLBP5F5HL/r1Fq1a7CjZqNSSky+
ZRN8/8rTCzpza8SgMS9YnddZT/Yq7h26l9+0mohT2AJYh0uCUAA4t5JK/L6IewUHA6UMN0tes6HE
0s0tuSwiRzgi0sVluzIVLzQ//XxD6oz/GwbLqgJft03fVKu5swR7Dpxf1vobohtSWH7vPeb4WYWW
fCxAlrHP4RNMztm4CJUJ0EgKHtwecmV/UoYZ4DSv69CfI8tTyN0MXth8mm36BPTCMc5fmR1SFDjq
1JrMLUrasUNQzHy5kZwsSMqQ3PlhNsipxOCakOmbVqqSFlbVkzcJ0JRIlyuwt8c7hWH/QlAg8Z1B
UAt4wf0IQsmjxlW/4MizMAThmmew5r6MUCLHOWi+PksJyZWFEvvuXbSUyrmoEldpusipeutXu2kp
738URUqFdBed/vOnIz7Le93b+uztEEn3AkJttOmb8uMkrN3MA6m4oR6GFtoY7pE7Tdp0tW2moT+G
Rsm2XnC6ybjTfgkrmjx76/MjYw9eiH/74UlvoriEK4bfnEGL/yYBMh2Fn/BPEBOofk+EOgwNlpU1
0DCAWesgwfq9gMlODot2AubT9Uopv6u4ROoJXLT5Z90pZuD+UcRY4EoKwCQ0A/4jX8ongHz+nDiC
15QywDjUxpkctQZkHNGm9WtwyhqICGglUtlGVeSlhtj4kqoIAjDSS4Mf1h4yju0z37RlO36/8ImC
7q+actKZGuTn4csWRaV1Hyk2PNrFcLJiMqZIu9hs0NawkIbLOYaAmw61MLgmwGU6xlFyptWERNvn
dER7ChXLD+rPLBL/BKHCCgi1CUuBUZEJGwFHxDxtTBWrglKFN2PDy9HxfwzTHZtdarAPSelMxM24
ZxQ1Uetm+nBsYXIksT60oM1+W9xpWLtSE25emD5f2mLH+iDA/lY8M/CxonUSd8fdDn4ANiUpF5X9
msrY+xJ9X0EZ01YSmFdGfMZJWxeXUQ2VSZdqiWZ9fKJ+c10JZxN+zCajTRiLK/V9qFCk9O5U16Hq
5IAwmqKvwsXJdKEfTnmkabdDWyUszmVnZ0to6i7w33u9U1UYFVXM8eEMyLmXvxaBj++ydgfS6hNB
HJw+wiZmpPbEpyDLIMuvLKcGgqyzESi2oT00jfhzr6olklNpQ8nFbf4TzOv0nJY87BqTLwF2Diw4
nJZIsf9oVuhbYjxzRLWVIs2Ttgbg6cLGYCtofXcXnO5G0AKQM1ZTTOFcdqXiODHTwWj7s9Y7oGPZ
0ZopRUBpmP62fw+2VzpOGp09mtDApsuIq2FdByak154gR5P4dV+KGhNtegDSqsmTH8Cmq0SY/hjF
NCkDJPoNjmgbR8vx7+jWihP9G4wJeeMCrossgt4ayCY/2zKewfTs1m8BQyQQaJJSr+Q5bBJ4/4cx
NqxUT+I0bxJsZwqXqNv8Fdvf/hO5KVd0b97p9GkbaXmYaKp/wJtVq/u+e29LVC06HuMoJIjD6Aq/
Jt5LshWJLiFXE4GXpGNYmAaeg0OoaXmZxihdjH6gz/wRUeoLZpz8ryaYTFyv4mSLj7vFhYmUpkyp
YJaiCd0Xrn5IfQz2ZtiW6xns/6g8qa2J56Mvv4H27GO4F+Plcfuq9crVWyW8XrpD7TspbjdmDnOc
3zDVNSlze17g+m9CGEl62dosPRCm017/c85+f4V4fEgybAO014R7zSntvELdGSGWI1dQJLrR2SIi
oYxfzLgk6fEzEV4GY/d4pPreuu9rKfcCq2hxMbdvwUEGTHWljRhjDT8ccD7Hl6G67hqQPB/J0mx9
1jSde195NydhJGzf3sXiQtN0/Cn7CQDl7TkyqWWsdtR2/PiqmOH6+wRywiDO45RXsKA4EmNRXkat
AjQWr2Td12JiMrWvAo4mz7BKFfME373B4tl5WYe2uRt20kx4jGP5tkU5xeBK55xlVFCU/cW18fnb
Pz7FD9foGZdbB+9esJmQs+kBhGc7X4+T04cUxJsby+o6vtRnAEWgf0pvlu9E3ibKF7C3T4ddC3mG
6KIFtD6xnWwP32I49vC5NNNGw4PON7FeBFhM7+ySAchzS7qB3M+D3lc/LOWNrCu2ujvp9Eef9sMV
akPTZDcDj/VF5lir6ehtG3iICseTjpN9h25Ots6rlOqQ1et39By/+MaNn+iA/uegrjWb6w7zzI+q
W9U2xkh2lRdvPQe57u95MeY43tbA6h6WMOpXu+bFxbAwG4V/p1Ie38lkTq0YdTWAXlHy7wFAL2a1
30lbLqN68vvt3YeMwuACYX0wDiJ1HxAh7pnitX/h1jSDstmdNOm6+YM43s3Ybtkwh7ckTQJYLAd2
lBol4lBthTt0aMa1LKqGNoKsJVgAAT55RffvGaiRzef4brkoNIiQohytmLwjtaLunQU/kCAfkzdl
csj4968VOnvlNIw68pcK1TcJjjT/fQV60gv08jWTS3yxwhP46F4XA1K+hWmqdN2rd3CtmOT9a32b
962cHpPMTx+ZhFeRsSvFT8F8GZyPinGx6RQzegqR8/DkEPT1vGNVgZ1GoDw666qG09s5hmXwl3tT
+K7EcZs2r6m3H8lMsyrgUhyuK+2tyB3IRHSRbTtHlvdG08Bn8TZeWqoLay7xb4uyVfhWIJX2kA+I
Le9j7ulV9jj6IfEgyRTTVWyzBR8msZU118IQT4+lAj8R/X6eUmfoy46f5yKIvnlvCO0zkqMxzaqc
mv9Jzg5lbPGMkFXecKWVKud3lL+i0uNmp6HVgPQu7CMD4SQtQbdM+/wPEGWVMrNHMBtfwC7FMVO/
eZfPJ454t1YxKI+PmMqGeaoKU9hd+ISuH2DB3fXxL+K07RuV9ZVGqCGzsYbH/VLJcMSHVDR8Vo12
1G7hp6eUifvpT6jTNDMwufkqVqCSPChxezED1w+08vc0px69s2g/yOwsIljx0mV7Pr2ZNKiw8etb
Mfg6etsYR16O2FJX5P1+cP6rU8QogJ9ULL29+3mZbkxFFJ3lNOy7r96Me3eL6eWH1LD2Dw0VMsVk
eNg+nQ2vH5w7sSWvpHoBYh3ctQpyOtGDB4CKBk/gKjDd4hHKSvUMClF8F/Dd97eYqvd3Ari7P7yB
sLI/bBHhtrPuaMUrqAII8WV9qUP6/QTctIlmdhRrEJ/4czLsLsQGqm9Vj3ga26AIrsREtiaT/RYD
m5QEhRp+4bROrdvl8/z1e6wye+eZNkYzt+8OXRGF21u1Sp0bI4y8Sk6cUONUH4fRofexiUqn1UZ4
PSaeGG8BBsJtNdifOhQr/y4MnO95zzOhCdJZ798g8ZGXoezBt9oOtYvu8/iyB+RzjLMOYoXW0iPe
IQZc21b5JblFKy5lxf2YuzgKF13PuL6COghC1ORMfb+e4PpwrWVYiOepAivYlw4+S8bzRHHEf1uT
QS9HXsXS2JMGpA8+DmyGHVCv9jpEPMm9z1WT7fJJOc5M4HyePxuCWEqAJ0wTyKCjwytk+l0XW8v2
Eu5ussLoi0pXuGQu6j6hjStRA3dFCKhd+pEhdNEIh3gbxWmRMFTDNE9NZzLqVDfzsQGRSpDgvL+I
8FV5khHbFC2BR7D/PhMQTzkXocMw4mQMbR7JBUYw6DwqMaRlkb4qHdGjIu+T5lyL7pCQokFhH6xQ
qOeoKfP4+vd7ZI1yhcZIuoOy3q76vLoazpiv0gfF4oYNuhzv5/2hqWFotZ7jr6ZZKMO5rlBqwdem
s2miax+uUEJmSsMD7eZrLRTnCHMKjHBEVDiYyQ08bOhIjsWFnX0h1ifsgshQ8xCBHcLW9XXpy5fJ
+7F8dSa+HL2hRhNXL9aYA5a4rOuMN//DajNajgV3NjhBKW3cuqskHVcz0Lbr5wJbYVWyQHjTuhIK
HxiZ18FMmf9dYc/7Rv+YLsMiSc4k5jSblFzHJi647SvONirX9Fx8/DxcpEw/zcUUDiUkpmnqhzwD
sDUZE47B0byTI/2mRjVthQtihLfTf9iDxj1UdsWxwZIYlQOwgmKAN1W1qDgFsBbjqKXn2UmGYDva
oZAVhspGcND6JSt4qAjxR3dXNnIDK5hVZqQnPA7lpJGmWM/ZeW+jvzUdVV0nWs80S8rQvWJp/eK2
aj6V7X9PjuC8A5KaAozw3xjERwhV5TQDb8AvvxpWKGI1gOkOvhoS/8PEbYGWekeoY0SB2XnH++Dc
kPSgR0KTkXKHj72gG19kvyeTUnaQixwtSEF7b/dcMyOp6RCvW1s+nu0+GrKbJ/alOpUsL6lnbKNX
H371NqHRG7OkhdMpFtpm9H23XcVz71KM85XcQoUsy4B13WaeRO08qocyOOL/bzO24b/BAmOAnTrD
oDgosuYplW4UFvuBwKi24eVmD4uEsmsONNgFUV6c02DSaRKc7BpcVSO8e1+3eQ4A7XushshOWpVc
S2wGfZWgc0LKE21vUTT4lnuA/VekpUn5j5LAxFU9+IRCnCyXb18rkrl/zcgKSzwg7ff1KnC2GPRP
miW7Xlgp1lRPoSkSy3xrKQ2VzVXYca+TenBC4VHyUAZYyzWo+A0zHxmUxZjb7Uo+f6P4KIHVecOK
2EQpKEtoj8cQKiPKEQvy7ZFVYySWlap1oDA4rLWPUm+GI6YZ1xtyyExzU46W2xNvmAGojIMSLHLU
6j61keeXSboaX/CVIwsvlstlKcfBHA29xTml/LePHhqAkMtgWLCa3IWyF2ytUXjIvaxSOE8+JIuN
k6+ZAM67rHjKMv/R+18pm4WAKpV7P/VMAdMuGEhr1K7yftE6iMyg6IOkkgGogWM3McSl1KKw4V4t
1CsJLRqWpd+2+HY95BDUgh3PdNeaUkxDFsCzfBYFQBrEa+qO/3Xp1TNcRDWgU7QQZ2OE3TViVi5a
P16D19NuE4aX2D/s4KCpfIifhlQ/P/m1Bge9AEMXVIrjyGgLjl+vPXHCD2igONFTSzUZvaG21BDv
BD7Z4mi8Szs6SdE/lLUsXoPMg18XMdTaWg3rFw9rbUyjycCaBO/DAwlPpVKh+iKNjaHeA70rkKIE
Mezm5pUf0gkKn0DUS9kLbuVVY50/X71d2Bv5wEJNr53jDxwApO4D4wLlmCi22FWUQ/5j3TADkDq4
3ESGW0MFkgPwiFMOBdH3dpSsrw0emXMQOg4HNK0AprFFd3XLXZfoClhCUBQHZxQLqSLQFckNUVdE
Lc4sPklq5J4/xPbtipdhFmZ5fG2WNbqvj6Cy6/mLcbXrVdNoMRL77ZR2RLPr4omcTeshGoxQKOIY
lTfadx6cmie6Nh8Gs6mPhe8CCQ3/lNmOQR3q/6XaUFREtc5Ta5nqF41P684fb1KpN5jU68+5vE3L
lmzU0n5nU/COZCxo6HM80DTRymHLskEIQgpW5MTFsg187x4KJAJBzaXab6jruALBp0g+/Vgc6Ppt
1r1uMDel6JWwYJclwnsqaAnwPwcjxajeNjXdV4KTBQeHlVXn+pOSEFWJkUWlRhBk8ZKPO8+25vQb
rqNLfTpfChhAkfUgY7BE/dFwft8+b+z20rg0Wb7VGjGJuNCEVAbgB2QX6vT5GRHDGF3cNojBUl64
2yzgSsdybs+UoL1o5RQM4YRuPhDA1KhEBblzuQ8VOMTwhmsxAsvLlmLXeJxiLDCE5ZvOZ158s0kQ
vplntdo8yPvA2K2wfcygreQKd55kHO0Fr5QGIqjGKNSHIAjLNqfuj0MWAVB/j/fzOuizWl0K9ic8
CTgaLLbWMsUpJ5V+obBYAb6/ezZjLM6lufPcd4edu2d8VP0I7urYPqmJvlKwXSaFV/QZ9EW78av2
KB6hwieuvkzTmVfcMMpNK8tUdQuTg3PvOsqPd4EAklWQN/WVjVBe7p2HpxuUN77RvoSKltdnEtxy
jVNSOBaAsCrSK927WZu0+n4/BFV41gnAIKryqMn801Axaqf4IQ7uidi9ME+XxReStOZgBPBrQ05y
jDKxi1kN+0nblt1l0/lHsZ4fQiDnsXbP99Y1G1zNoXjQQElpUb/kmDemjse9dgMAk1z37zLWNjRW
muBPpPg5kaO90mRbGx3iO9Xj7W8/twv2+3DaM51dQpVL2HVYAMOT/sd/tbfeQUhLR0SSVeegZ2Dg
yPjTQ/HxYQ+bHurqcnMJCmRKA8/mmKBFhXIqTOypMJwicQT149JXYqJQGFA54SpYG/wdELxWQxYh
vqtCScO4qly2FWb+mkNXDEny040XsL6ExJVcNpWB2mYY5cauqfNxVOTG+G1yQ5Wi0U47gnwowE2S
q8SOeTU8E+EkMGu/yYgiJZi/pYi3m0j8Czdqk8uk3yhsuqLNiNrfWK22MotibgudPe2dFBkpHO51
l6GOsfh8F2zwJaM3J28BYfxs8hilhSnQv8dDAQ0zkvhNQpeor7VfyCdSgakONwN5etVFSV6bfHGI
NGW1da6pcO05rZR8jhmDo0whjmiaUP5FfXX2KQOQP3dnmM3hJzMCVOWKHKOy/GEC2ql6IuU1RiGn
NhdFTWznqLybIJJkJsArYkPmG2wegxBib/OETbzw6ElcGPfybNX21V5CRen1f3IpkhN3DUL71qKi
HjeKU3iW9nfx6o6s3iHpXK6oo15gP+fd+wFycstRunkBtXC7k9KGioKrCy02KheWWEzuiH1H7T5n
SOyTwncAaO8oUkTjB7AqoDzs1gxU9Fs3IhhGOHVUF0DPUc91uP9i6cWUDRxhE/kBxe51PXWhIXa0
fPGBn43bMHpDAO23urccnuW5ccD/MeAckuv3aVZgAgQuX2fJ9+k02Z/dMjuQ7xoMV0LF+/L34bPT
HfV3tuB6H93qfc/K/yz6/jUOWCq2bxKd5cXT9sa11c4qQRDvOvy/gxp80TaPmkJqTkW1YtiPjvsw
g4Hy7Qk4sG3sYETI3r7iKF9XhQ/Ky56EQCoCGxIrc+WDSSGvcdWvE8xEJFZnWebVRawToUD3uROa
qa2kBY6BNHD45R6rAndnKTMnsQNeR/rtu8aSrT1bFQXKj6LgiC/xKE/T+EO8jgZVpi4vfNreOZPD
jo45RtClBnooheq2ErM3b7G7FCgHsSH/fdCZRynFfqo9GhvjVCKVkXTo4utu1f8H6z47Oxuw1yqX
V2ZZadEJDLQ2I/ZMUw6YqR6xsko0HlvB4vS0Wr6C5J83/s7FfMspztyGNwMxujaLemSeW7YJNomI
YZ6kogUTyn0o4+MYD1IKKbb4jPYOTkqqoMBBgfmyJOd0pgmRNX+hRqLFUfmY5e9uclz4cxbT+6hT
u0mjbr/Tn7IpXV7ckGG+DDmqQGWz6kU05n9TZh67m6bo/bjHCfBGCahm9L7uhdHqtMNP9HqLCcFB
miKvpR1+Ruf9avUFHfbjNTFd1AUWZJHqWvj0LGaPsG+f35h0zXr9zuCpP05EEeWU2Irqj0dF5Pth
u5zHWpk1ZAjw0vt8xXNDAY9VsvYJvXi39113VlLN49zb526rPRbbog/3eU8z/y30Z1q0hDguxxOF
HCaPCSOhhNCSPWZuINBSBeWgq/KXB0lZCnk1tYw3ZJpXiqvqE+VdnjHH7aShBXu6ZO+0+PGidnAT
uuXOzPPwfsJCo+esO/rCmUC0sOyC+3oNxdbtYzGEAUy1Napsf8C5ecl6oyF0LZj41p6qDeO1GnRj
ldhxrM/VPhitQLXa6JMdgSsmzwjqVJAOr65ioH+ZAZooWPU5Z2zpTMtA1b62B9xXwWyaQRfamVwF
P8BJFf7UV4Xl+zzy5KHL9a2tPS2pXA+hpmvZys/h+b/Rh+9sry7D7AM1TYqRwOHQogT6mhwCbOq3
m8ZMv5BIs/qQBmczLQI8DdcmWMS0FBelZKgdr3ehffpo5TM498V6odkAMjK1SEK+k2yxh3wrb3Ti
Kt1TDItlfkNNJZpEv7uOe7jw+A7a2qY26kf4eWXYRkU+kNKCLDa6IoTMT8C8yb1eOP+aZaeWMilI
li2YjltVnrDB1UMWSZ/SVrCn1WuAGLbBTWpJPRXu7O4WHrD0tBSFUHEbCwzQ7D5d495qNnd7gpTM
CsrWDWSpFOWZ8PWY2hhEB6N+OxJNnEvG0PuuIlL+CWaxnV8G0D6zW+SDWxh7tHV/6arnIY+bFD7U
3lhGIxuqP+WFVLUvTR+pznA/8BUa7ahbSXwr6rvVIkN5L8eGlSnyZ1GRYvo61NpgLFLrTWaVBDlI
3YE0CDTgPMhHcI951HUagdPVHE2NA1ywwR57hFPuQZG6j+NUPXuCt1pCMy5oaQJ61agbYkVHOHW1
M1IIXkUNV9rQKIDA281Us8kZ49drBVpzc1/Z2pjWamMqpR4OcWEEYOeHaclY6hKPt+wRvbmRIlW0
vmhXnBtMeatEfCgJ4pgKfLwqtEcsT95qs4t57ZB2H6xqfttnzPBwsuBo6JArrJN4l1F5+2eeIMA9
D1LNyI2Q66wTiYWiMVdkdlbAMbgWBLfPmJj0wGHP9lvbSZAnz+fMnPYznJtskArBSV0Yj57x4gB4
tkt5wZVvgrSF9dq4Wz9o2fHabv9ADzQanxqL0ANDXNE6GxLRz4fa3esmHLWrrgM8+Nz8ebsOwyVa
gt1Ngb2IEj97ePm8JhjlE1qDe4B7AAnxsJ91XkqrUtzWUyn9bd0AkGI9f7j3VVSOErd/z1dsR/Lj
iM1dwZJKWJbYOkd8mMNRISiTWEstoeoztU+km6Uwsj0OShWPfsTzsh/HNQsfJPA+H7ZvVyjArd8v
Ntmyns213uaY9+Lhj2bsdL+y0zpIQn+wQz/2GfciCbnAhzanqbTtJp8b77O2dm32reDIme9yZVe7
pS7lEQJwANES0vfg5R2MGFiD5NgT1g4t3qHkWCJthtNDWodyDZhT/6jlYYjFGc357OoSAj3j1DVB
uRhkQIjYfN9JQEJnQcCCBXLPhdHH6dq7d4UtoTTW5F4ooqGT3uXri+7BjPme/O/oJ9WiYaYJHQAj
4XLpJd3RasPnV+8dPiUXDB4a8Q4xfq+xKTFqolx1FdtNHOgaVVUno0BIjmLMK7q5USw9IoX2rOzA
wJk/UvsSnWOIekDdPj3g1reb+B9NEqQwr31e9nOZ2IvTXjxohMq0rUyo83/9lmzb5IvMuoeIybHi
Qoh8aKBSPQY5SRJjODkto48CrbwVpeqIWbwAbWGyS8LUmcXSQDZe1Wmq/LYD2+MtoZQBA5D/+2fv
EOkOpBkW13XaFzXJ+Jnpg/X1u3HXj9vlF5lzb3KrrRZ5U2YLg0hPvqxYvDPaj7JV+uB636b8gP9x
nUmxnyRfJYZMLu4swlDq6foxmcOSDr+pgFbNKjk+w8Nc0yMO4DoCTAKgv8nq2EVVEuEwcTRG7ylR
cb+loM9AIeeESxEf6ttKfkghL1QkteeQwZLIChTDxoLHUQ/2Cbp5uCVWAKp6OGALtNeJX9xnlxhq
3zqHP5bjhPCC+KCkhLPA+kWa9tzi1YGXmZd4xA7neV2Ahrh8/s3aSRKAivurYTshx8hipZbIlp0u
88H6HOH7ck5FY6yxHJKCRclEeb8CpbShBNs05Q7KSan2kqVSoFw06MSLSUc2yHU4X8Jumw3EuG/u
2O93gbYm0pueVaaI/YIG7QQZn2HqZmA7Qneemk0JXT4xaXAvaN1JN8AhWwYEiRwiPmMqqZSnwxAr
t873JUKQsMI/C4d8tY+hsVf4Lqd7U0L5c1qgPfe9aB4SdebvpwTK+B/tQGhoyrkQLikKr/ByQOSA
nqzFPH3tYradyMAhvu/MMh9/YHoT2S/Dm3hdLQsfrdlLxWGHaU3KpaUMSZGgMYH8IWHCT7RYc04f
ARypBBc40Gjb2j7m0CD3aSxDi/kE0/nSndzB9wQ/zleSlq32X52+3HExiIx3rVgK/QbngoQKlqwk
/L/0eR7vKTCDrnzjrczQb/1uoh0WW3THeRJS1k41MGDay1SzitWzCvnBOenJmhVd+BBoMivM6BUC
U6qSLz5+UPIdrMNSd/+mdji3RPvvuyvgixYxfhuov/HhAp9ypCieZPcJiB3ZxsOX35sfrQvbloHV
fQeHwGMdxvHC9wofq7m9how0JQFUNFwmlWIp2ySAcf38OPzVwHIFIaYURttcsfPoSXkmE7MC56BA
0AknLhNnZ0Q8zj8IEKrR2QXDXNkJ0IjKPfb8mETJSqPvMJd+dc9AN+ILZq+x9sowv8x4uYGOUzEC
BieignzTqhINiBufE2eBXy7C+9XIfBYoz1ITiftdWSXt8bpQb91B/qOyCMR6i3zZ9Ia3bo+6MyJY
IvYL3NAvl3v5UovgQVwaf2QVROHlwRrNlknuju8Fsr4NLrXJhlqtYKpHORbeFGvInsDqjxq0fVrB
kg5kDh3yDduYdQUm/UkEFDP3v2w8QZduUw1gc4xodPGY2c+QdihE6gSkyR9g1HpgCQhlp/7mpykM
UO6af9TqYls/70Pwc1Q8rjslOYPgjoLDzGoOg0d68JaXwbsKDW8dLjzfH7d3j4wG8wfx/UkCY7J+
FgCvL9vxwU/69MgjgiRcgtrcjjVPAlgiJefAjaNdg+Gs2dhw1roY5NXKMXxusACWlXAJXG5g83zc
bybS2XUSqoIOqz2v0714NIeBC/nAhVWTFwtRMazkAb/pIzHTU526kRGj8CLGkRIFoYGvjiklD0FJ
mnR1vOkpPDbldLSwj4Y4CnsqHEQrPL86iwvJB7T+P22/5ARKyZFl7LNh6fmnxDVfC+tQ/S4XVwTm
f9D9fS1qAu2DP7e6G4Y0GpMZnYB0tt6XuWddVxjV2jwJtpdvqpiwOoJp+x6hvhMJCLttCw4E+Zb8
mk3dVZmyBKWXjNmVyttXFDfDg/Z53jCsNMXamKVjDMDDcZFYc5k5Y5+sq83exp2bG3zm+TnatXbJ
DfKzh5opnlnuGUJUNFsRSxOJfLiRqao8IfrCN82+A9z97IPx601J186k4ev8+mN/KeIB9JjbLkcU
AzrrorARVZ90GivMwoXEiJSPLqbfCIRoNjZbEIvJdgAA3/HW0crd7QTWYJmTDH8M3A6NZWSf4VxU
9hAI7PJpXEcO6sq2V5xvVDGq43N9BW/a1Imv3BAtENqxouUQprr8fPI9OF31yHdS1JSFxTCh5z8m
sYje2wdt1O45fvAQQgJ0FU8dRQFrKS0SLD4DrmHr/jQUI8dZRjiUDZk3dItHdisdSiN2QdxyOEpx
7DI2JI7/WOvlx3AkffMve8ewiiuj7LZyEOa1fL+fryglAxuNHEimJOtkbSGkM6MMGlYrWdYoJGvf
rSOSHVSJWNT5HnKFa7//5W6EUgeYgC5qCGegTDyDSOoqqEdUBBLAKR3i2xk6xzmpKGYOuGqOLz3K
kRSDjGU7w6EHjqdsNeRpT8wLbbWsZU2Jb+O0rNluZN6erYbzMnsNWCZ2hyDoBn07HvJrualuRulN
dZcXz9FAa0fzXVhvg8e1TcikT8lnEx0ZnNCqW0vtbYJDS5l8pHM2UN7KtXuitGafYy8k5+o/89sC
fcSEJDMFEgpGZMH/d9QX9ze5Cy50BUP1eXbQhbbDp23b6pX7fVDugXT0HDS3MPjYbUdq7UhA+vOy
Natvt4Mb9o3MoeUcmzla+BGn19KUQ/vA6KLxhPH7oLs5kd8eu7/9qe5UadpJsB2Iy0ZJC4Kx8pAv
h7B0Dz7fEDj3ijDZRlzVh14hDA6JGhDQ19/9Otz3vUfFFjsFMFxpd6Cje7ZK+iXY/jE4KxrN02zR
pke7NipsMSGYBDUMJHBFeLr9foMJUynxVk7a0PS5czXISv+V9Zg4jPcnP2oFKazR+wNG/BZUX+IJ
vd10zBv16mWHGUUmUgw1iBBi4jpHydIPdmKeJks3vEi/mzdCMNp1ZO+eRbhkF6A+pqvIBAQe93My
q3gUJy0fvVqXSGWmhW22SkK40x9ydIckXCU5LFkSCXFVAUF479Dl6QGXOjrohkujBQdhs3E7WC3N
g0nj979xcvOKFvFfhOD7J15kfKZRDB+fqFnpoCsYV+hUzAU0G3TGiutAxCSc27w8XFRPqG+OWZy6
rwR4JPOh4nyjF2FoK+lCFauWKyeqaZOMAo6pSi8eYBqv7gWJKh+ypirka+PKaGI9nrUDJQZ8C8Dc
/987tg82Ge+60BPotmthtu/XsPahMdr3wZ5EmXyglogkLMnR1yAm9xMuGFU2HIG83V+575s0V99i
qYhJ/1LpvxUfs7TXBybevy/tJKK2S2RFWRmVun5VAB4DVK8eKi9ccVHqfX7NkIF/UTn2IDhVU4E7
1H3aIttrUTfGQw1eak3x0cWpYi4ZMlhbsVf6X6FCqjXHI9sWfZr0vTo8cHu2a9yAr0PdxJAu3dUa
BYIsmHrcOLlvwaQPe17tjB9eQ2aovmVFwq2q759QwiVmbyT/hAUulWmU3uw80bwfoV4uG7OeHscu
ffygQBQXDfIwtOlvysE7OZVLdOBN/lkYYLi+FAZMvYyC4MGdIYogZpZz5UKTzIJVZuan8hq6zO04
tdNAkm3u9SJQ0cZRT+hxxS5U53+KkSPciYxX3t8u8Oy3vGvKo6JepEkk8GzDz4TiJ+gwtIpW2qPf
r2xbgJBAFf3puAsgQhB/LI/k2nqjnHp4WRjBUdB7vKXS6kP+qnB2p5Qq8y6jQd5w69oxWv0RRKJk
HPYvmJrcAsbObLBiQ8hLGNNzC8DXZaYl0yvLYSH1PYgpmbOF4onM29OWui3t5yP4D7SGgEzN0ag1
pXMnKK6sQfVVgw1AzF0yoLpJwdjD6xVgBdpV1M6oq0qw/+tT4hGiYFh78bdbVP9Qz0PNMt+QSmrd
UVyRNSGJDidDIeShg1euPZUhrxQ/iHnwCoae8VMrT169pu4UZOgUle6CH+kQPsCVV2zjHred2v83
GwL6wdK//jj4qXEXwdCo4AG7xRGmjkf6iT4gvVQA3zdbb5DQXasUztawK1d0qkAONK4qUq1LdSGr
TNgQ6DMiUzNOdl8DdET2AWtvrIPfzUkpBszeovcgpKg4aZvGoP+Lj2jxloMbwww46X1E0cUjyuA8
qG7N0yD2dJulaOoNZSNmno04HqbEolQSiZ8dPhsk6IAE/PXztl9Ztb+bPtrcLutYrBsW9O7tbb2G
l35RTiuHFFYTPlP68ZQKoVhNChywuYQOPAkOKbizVfuyg5+mkprNvrAB4k28AcuH/AuMDcUFz8jr
Hx4g+QjH/tDRwUfLM+pCUlwatTWFFqDL1x+jaZHpBUG1oP7KToG2ftzE5CA9BLtIfZDhy0Ha58co
ydOLWMwxKozxTy3KsnDB5HWe8uRxLgLVYImOx2jCyDXETQFqURCMl2dBTCX2/skWzsDC1ULZ/euz
SoBgmn3w1jsbC4Jp7sizsYPj6fvn9HMCv90h1s2bsnmqFHQn0W6yVT+MmeX3XlRZ+6hQB5SW5GTf
Tu5r341VmnnVQjF53vIf6IlncUzJv6z9tgirUHh/DYOF868WP6jAqsKLu3GefxGAFEMrlCYj6sF1
y/rf+9klL+CW0PBLP1slaPjcYJjRCj4sQJs633Jg5BPhfSe6IbeqxXP5qs2sPiHSlJyW9959MF1e
4kZznE9g6cnWiMmF4SwhPSY0UGigzLsIt9ccP322bsXO8NL9g0F8AjKKZZ80429r7J3LIF80J6/0
+cFnT2Ncb3sKV7wVTjK4mHw8QzxfngUUkB/uGNBCb0r1a+RlwA+pAeTuroFn0p1NizEvt/Wkr/wv
RxGh8p4F1zP64hzoNFfSGQ5La8j5oALSC0bJsM5p08iNzkbPWRpLNWJ4xaoNML3MRaI/sBiIdz+P
wtfDgtIU1mp4eEZD5HHu/uRMN8PCza63r/ISLUbIQtOXIZlrT5OlM39VkJXYVLoIyGg3VnmqG24F
b8/Vo7siJCcoivvC+13jaH+wYS93dDcM+4ju710IUpN/wxK6mkkUScrSE6iWggOhk5WycuvIFNFd
LfPWnR8c+xLYtivaeITjnRuMEXSXpwT2+b62JAPjWhsugyYwqPkxHTRBZnNI4SPtrOFp464BzHsa
xl4BUWhBDz4SagvyhmlR3r+7oZC8/uRv7sICWv2aLvwukZGps9oB8YWl+FspulbVmNlPKzpboCqq
F8ejUdic2CFuXmNPs+Pkuz+dIeRGKQHU3gFY+ezPbLu46Ym5Qbi42sWXDhkRaxrDezbKwKupEpOc
LEzdHblS2lhYaZ+Xj7HkX1kHdBGE1QvAMGlEeQApWZKWem2yXPZHXw8IP8sSIM0mKsOJcasVQtPU
LhSgwcanTMlgAKRL9RtpodocwD0Pa3gY4gfVyQO0bVYObiJxVgh7r3RUljZHaMskodF8yg4JBLRR
i+J9/rUD5puAJYfGa6sofmSU8wOteuhpsF9VsXkDP3wnYCBV4bO2kv3XzvCBlV7yyBUqWB0ps/yp
/QD0JW6F+brOIpILfOqxfM7e5AJlv4MPd9z8/c3oHH/lvmFp3Ovn21eEQr6LzmwuW3gfHSdfuEe8
P/nD8p3CUnM2cotiR8VzJLaQ4uvEPbdTZkoaNYd6OhJd+21XQY+qDN+XGYFuDEzUvnvvCu3O7uOC
tMFhpsn/QKoRARm/LYJOVyghTpKwfquKmomvqR0XWfOUmOEJwD2PC89s8DfN1zLCGW5zaCc4w2si
khcGDZNCnTXttrpnzP+ufDs+IkU/RDnoG5lpasIFhZboORnOLI6dR5CAUbiIJiFILzo6PJxbRtFb
xFUVRKZFQIfYGhHL0HSuErj+vgVseUw2T8ZoPRxu/YmL4jFerrF325ryG5gqzlfVYeAfvqfTYBAp
CKrHvCQW6d6gSTtrKImESB55VC3TcmJxkGziNt+0SUPagACHqeeXur5YxQ6lRLINxE7N/VpuRndT
vR2dPWqis2sYeSj4sOVopAYOYfNuufgi4Lod352IcOkxWCK3HXS+RTXrGPPeRWrNqUCx4ppUKkwF
PWqH25ZKN1zKTgdcvpvf0nNX7VF2Zi6YmfHREiIiPTbiCF98MoVR/X08+y7Si0R5H7qTRNO9f7DL
3YWJlhfKVPewcfaB5fUYQI3y2QycWFLpzv+00c6PFoSv2hXbPg7fn1IaVLoRjLicL60vwDKJpqyY
ek2Y7zlplGlSBGT4HYswAIqDeZNZNztl6Lb7n3iHSKsFjnGbCHD/vkwcwk8oXyuHYxVa5EIAeKWQ
aBU0IWEtrKua+d09jFN+KOLNCDpl4svqQ3SVOmCEMz5ectf02/2S2Fqg5IEaLlFqskHOrDYUm0Bj
4Jul+w3sJhIST1iong0lU2z0iuyIyfaCtxzQVFqgbXeHE0stvqqVmULP9BW34Umr5fb2rC3zsAgA
m3wD7echzSDfQiTB2a9QNVgflidfzLU5+oumgdPwcYhAPq6tyj/gD+jQHyErop7+BBl/24dicLOr
gzieo2awh620WZmGEZBLFllN9QiTWBooFm+LHNiyPwlPU31T+v7JNMhdHRjMLMd6BiDjD2gW9uT3
Sex82fz90N6sqVsq0/EmhznSbt+gNvjtkYbeAeX9sHo0Ki1Yjd6jL1xJ36xrs+CUEnhpzcvgiRay
W5pYWoEeDR9xRXq6ZDezW/c6vUS7YWN5T2B9yuHn/fdwXHJu4rQHGVyH8XF/BDyt49iM8Y+AXEq7
PGXyJEBf4tDbYnPWBUo1q536jA38ey7HTilGdLW1Uqd7LT6ENUUf7TI0bTtKqbTvO1Fk8PvKQsNL
/9p9nLMza0GuTt1n5wQlIec0xgpXmpPyPgHga4e1rNboYnQrZWES0QQndTfawEx8qMpXZnkXMDBm
TDQrH3xYUUOzd0K/fVtBwTj/nFZWHMqO7j05RA2wqsXlhv/W+KdIKvhLPh15iZY8QQTmBG8FhJfi
DLK6ssQ9l1sfRM529njpwfGa1HVHLmEsxCcbZcVzO2zTWmqd7ygxXS9xXvvqRZpPYCHripKF8YW4
772LmWdKwrz2ZLNBQwHxbX0LlWGLRrFuWCzVVcR2GupRPuMsNYRBRsv49BK7ie/h3uyZcAyM2i8I
OLKdgRXIjuluM3aNqNBTJohd8f0wAqrUXoS/E4FnF8eLsdOMYo5hXSaxDkKOS8XHrfM4afRaYJ4f
W1+yGs7yEhO3P2zUrgmveP4M6OKoBwgC8q5qB7ML9+qqp6o0Hm7jTAfUoU7DWlMeh9ty4ZcCVP4m
NYPqNlssVIWgqgkjIjJcmHCqxsiimIzbTK13/RoAZDfVPgU6cEkdq2l2bA5k8ehahFXS9SbxWsIX
SCS/Lr7bybK7fV86XPJB6JrgYA1EMaVTQAS32aR9ZJP0q0Ofy42TyvgXiS8f/zNv6A8BqQ/ekfyV
RzJBZf3ia3Yw9zMACNSrA56pOpSiQmrxZ2kFSApeEqSG8CTlhhkQeeJW0wGkZ+sfGNDVwBgwmY29
45XWudR0rQ45lGh7tuMc5dVm57J4dXY2UtDpfsbaxAbnW9LQJxEElgxNa/HdB/PH8F8WA8ZwRzex
fLYESDF62wruZOmuiW35z7YsNpOAxdWqxJ1yN0y8NjuvrHwc9Chk6YMLNgumJn3S2iGU83jXxVHs
PfMQK5UKgNXCMh+3esVxF599D5bpW/+E19NU6Q43KZFmb1smTU0v/YjnkhWWi8NtSNmqbNNSJJUx
fbve1lXDZkZ2MFn59QzfPnP5DEr9dEJAEeVXoR1SsLU7QvFXv6gjNrLYfroMd+aROvVRcDAOZ2C2
ZMKA5jdgugjT4cnyfC8ab9oTXDz2wSloxDbmZWzyoNLyWo4mYgVYFKYKeyGm+R5MBShHdwhMSSaA
2v3N/tWLPytOrdfUJFdIQ8ag5NZG9lRqNO24wRnF/YMwNf9g+1QtEq/EpElGg8+kSb3DlzcBoV4g
AoaFQ9c1PSF/Ozz8eNA3qk5vE0sSkfuRSHXJ+JWcZBKr7NJAIbcbzPf1hVfRtc32K4lH7wzdbfYS
FbkahMAqWbLnB+rZa4b7OhPBfwBEDzv9yl/w2aL0iQ8NvP7N8obGYGwlFDc7nTWO5+5eZuDCMnJC
qveSGMecVP55O34pDcmMWbvXWmYvhCTYSJV+mpIWbLg7gEJrMYUpEb0WT90ndyI/kh0P88UTv/xx
rpCnv1niM4Ivyeq7YQxK6AM1a7Q2RxX5oP08BuAHVVlxSd51SktF0Skm9bS7gBr7cFDjb9hBq9zi
HLOxEleS61wDuJoVCz0H2kG3eXCgN39CtAppE5iqU1NC0ilsd9/EyQzp6ErVmpWZ6HE+FWJV5cOx
itUStoNn0LTG30aVGs5ERfmtbR4Od5STlpvBel0XWRnoB1t7et/ks+ASBvqz7XFRjhr/yiMEkTP6
t+ir4yYmhe5xDvR0ot9pHUJK4M61tQQUdx6SDYFUcAdx/z8e8iAFgUVKCYeKe+BZxJviZzwWL+VH
1FWnWDJeygUrof9/QkC7lWnO9yj/bhlBfEOaj9nmmAwyRJAXhHgoXzDcNUv/KSg7y+ZraeJv0B2l
Kx5C78d/ySPbeoU5iTfQZAl9/ktpVM9+pdmk1lFdoHZUqvvTpRDl8Egu74MvGLrEYmSUrMpTpDeb
fFfOtrtVTWPw2PqMuHTL90w5uC/A85cyinxPXalFYpVRZXzjjw0zv3QaZI/li9msGsAtDkENqkm/
sIanpGSta8HG9c0qxzrpEVWjGk8o1NQmnEORT1S0j25k9Y8nfQHIqDuGuGaEaIlprq1nbaNiNSOA
hHT1uBMXickVq3NXZp5dx49ZGDnnHKWil1a6slofbNZv+i2QCpBL5MNa6zoNmbTKeSH+hbGB8ue+
0GbUoOq9y+6eQPf9i+3aWpeS931ejrwXVRd+CWxnew4hWECg5hVrYbc/t57NX5UhAKkBuCNQVcws
hsJ4dhjD0g4lZnhN6xtcWvbhWIn7f4UqGSupMn+hHljE+DxerPms7MN55F0hQFqd0NceVG3B5CUR
gmRbpea96B6GzV9sZ4ZQ3uSyAVYsv/OnYMRf4x7TLZFdC4kOspLXdFx5eykA2Jq6VXFdkgYqPTix
FhjAs1mLbNcUL970EHq08dSwrLvYMimkgft4ANOZVnYyfpgOah9alCP7ymckef0GpmR6SDbfDXc5
tlsPbc46uQZn3uk3rdY6wv//vYpNuBRYs3Y8zaT9s8xJao5tt2dSUeSC/3nmg5QR/oNBM5MHV9xM
55lHB7fq9cexpwRf7gK9Zfgxvl/Z8lcz8DrByBlYMf5Exu8OIiYp/uEnur17diMYvHZLuvHUlBBE
qFYprZD5jSWZiYmR0kajKM3TtQCiaguNTB/P3YvSSF7lhNVkSY1NnM+fiZJT/2FqgLrAdCwjbjgs
VAC/N370uKwGa+57NMX9mGdQBhR54OJyxZLjE8SUR8v+Q7alPRKnT1OuXPPXf5dKDQHhwS12tXd9
joHgMZFZqklkKX/UhqNt8NebAVtQnpuCtMA1I8Y59WY9kvwW6geTFHk4Khvky7pRGJudWzbykwbY
1/0ze5j5Vtpj4eR0daUZqcUysJLXvoRGYGIG198kQC+gTHIYPXtoDvbI826tS+x540rg9L7m2LuN
KY0bBqYHbEpBLB5EqRBxxvJtjFuDzoM/snpGNePSYKok8mkUlkEEOTKgxgtUTuxJFyaJhGFgnAzl
LGtZL1fIj9bqkUmJWHbyPv6Vau7InZx+M0fWtMTZs54ng+DALcJjyrznQ61dnLOSKqOdrPuKR66C
nUqL5+Tm2UjAtFpqm5Aiob+c6cbNFafhK4Ki/nhFSr4oTtTFVlHyilefDJnNfI9rB9/mp3Pj0Y1t
yO7/c4T+Hxr0tARkVOnCZ1u8ffKe+aLrTmZSQftHseojCFd3cVnM+dKXDoflPyFb8LaVqeGbAvrc
jSHhc/SYMI8Hd9MgnB656ufsK8o9/Slag1DC6csMcVZ3113C+rAaVAzAU7n9BKpUwLVZEuzeUhQ4
QO6lxDCnxEoy0hE7WuamQ5pwmvMTyL7YFNTiIC4cgAQI46BqRhqg/AUw0OlWdjHmI1hyq3r26lx8
zgzlHOknALgKLLTBYfhm5eG67KOAbqTi9IDBijnJaKHG9BcmKYuzWoDHkiHvenZnbIBxobUZsdz3
KlVWgvnAvIbHfOAH1CbVy/TeuUqTt7yQnRCrPFSW+42dYVjBmI7Bd5POB//vsJpRBdTnnb6XjOBB
GQxixvvkRWpvp5LNmilhEs/09ZBYIv8T0Fa2RH2UJxEYcveTEnehkOoYw2eW3spAF6bjXfsPxutL
Uiaf6NsG2a7ojjjt5KMgGN9eZzt4H9yRGJHYYvh3ZMKRLU1MpKbRRBFIq0K8oj2a8OQppM5jsOTB
wx2taFL31mBienJUUoWLpKiPcqMF/Z5h3J35+YH76h5OruJeqRGAAJPKeCXFHGzSiMSThNJglm3l
pwNUMuKWAWphfcfoH8d4lXPK77w8nWSwyuCaLapm3c0HUpCKh8+KtEGSX/mMIxozc0xrXjuWKBmz
O2rBqoDCsudOpgwRLJh5mm4qQemStkpgzomWlOzi9q0Z5auGt5gzEjGIg4gfONoocOAHBAz/KM9I
w5UOPB6kyZL+8wptdcBGSobyRqCFAR3f/EtBTaLarNePL6jJP+FsfHHFrUacxRVM15xl4e3+fSK6
DyfKl7ayy9PwmkxhFOY8I6n9aHtYJqseZIHm6OKY4OG8su30gZss+tCai/WntRJ8/BMjeR2iCUSY
qqHdzFgdjxPxSAmRGse45ZBzNSmJ6a/VCLyVPjtDvHX566qq8pEXJcXC2TLnPCP12NEw0dXObOjG
dnIWnbG+ICSJPIRl6vOdF2CICyJOI13buH+PbWpCDQnzYIKT7eCpGfh1Y9RslxlwwyoZPXCnXqrI
eohWT2huIecy/Y+9twKm5mSnbxhXoSz8RVWDecEdZraMz0mqDhBuc9zvjRdPj/3UBHNfzalGaQUC
u7cBsyUsg7u6VN67O6uJBXpU7j1ko5CAjD0cGmcx01xwCveYho7ohmS+YLbCpj6Arw1Ugvz1wZhu
YMW2F7RH7rUGW1ZUdM61HjG146oe6fOa8vcsoSsEvBgIRGK/I127MNIYLDlU6rmxdD4PC0eiApQz
lgxSavzVA/M5QVRxiERW6c/kPeJY9HSvavdfQ339IRQ13s1ivEUuk371YH0uf6OMITHfOto9h7VJ
TvCJYIjGfSYthLQjNzA/bY3+dqYnvxKfPpSjUy9HreCmwKiS/xkXYpIn0uq1HvUOedS9bk9hLV1X
0rD46uE9cMUajWAkzwcrooLY56ROWjewzIObUaFzyqzHhY4529almj245NwphIJW2X741ioxV3iA
YrUjHxoMFjfgwHt968PX23YVGP+1Q5BhTIh1IKPWX4qlo8ytI7/9A1zXQfpCXvMP2JAw4J/0nrpL
/mXPnPR+0Xv9IpSbWgkRSRjS+H6a7YzNjo1IT+6DMRPrPkvts24rv2NfB/ftWWVowoKMY/xHbiwu
tqSae4aLRi6YU1rGLqY/iZTxFl1Bx9xguS3yJ/3XVZKZeY6yQBruTkuHUH9Dot97tFbNSmmR+JZz
3XMWR37rcqaT8Z00YiSN9EmbLzF0aZOy/aXaoB/sf0kpdil3ZWQ06AeiAoXoVCIYVIn+TG7kaPWd
edwGoii1gVoBunCHpDWaeQXS5J0CmptNJ89b4fBRQ6CmC86u8ohJUp6omMxoVSSH/2S4sgS3J3zS
N45CmfT+TqTw3nm8P898FQW4iYQtOrFZV5IY3AtxVOF0y2sFmdSnymEuQyaXy8i3VlY3AhcEk4O9
xDU0AVUxyGepbv4U5gC09Lwq3ECwrED8J5jjhix1hopOKbMcG9GfpMYUPCGCdzyzwtoAyMMOgRZF
8DkSrNzslQKaLQafMNm3MV73lVy0+jv/4NwTKYLOofqgEOZ6aBGltmInUb6yEp5xWyCFZrZxHeRG
weN8gMM/bBG8tBXeL76BZr/rmWotbzTdBRyRrj73rrzR0NXIGEI+VGuZNPvZB6pmjaCYkcKoDwDW
zdNx0/hLXmUQh/+fChOuXwEBr+IkUfFgrO1urIHD1nv5mip8W9OVXP4S6jzjecRFztOAw0p2t4vk
Y9rReKY3wXe7/FZO5FxSHHp7THgZe1KX8CvgXAqnnJXO09tKPpJ8Fw0KgTo/ka8MLUC8Hrez/dpM
dWgP6r0+7sGlFXGaHXfYEhFFbDnmvOqnb/5B8XB91vD7Gb6G667Hh6aQkqzXR5FwmO3IF6dxe20G
0Zj+Cqr7SXR00n9lcdahgCN6INETxv2pe6LIi7JNxK7Bjuv763YjQ7cR2Yip+zE1RsJ1RyW1ltSw
Txdl4GRCp9f9HEKr2sp8nwrrJfMFDd4Bhwokt41XdjiK2IB+4w795HY5DK+I/S0jnQ77UCxXOz8T
4KcaelzZef7ptLpy1m7BaEaETG2WqZ3QmPNvzkqKa1tZagS+pX8n65FyqqenmmRtz8svM8axo+P1
MpeTnKL5ajaLvntJdRN9rc+VswhQSUHjfWmaLakEkHtLuk0DUYaQnmJ2Bc57QYyu8aQafVVI/NWN
ODLc9tFeywWc9XTh1kfhaqV6vLDrygbUP502HJvpB9tQULzC5m8kknP8X5XBRypN4o0iK4JQ7h+f
7qKRM+w/GR5gdA/Ckh0phAap5D+SlXheHl+xBorG17y1NZHGSnUYsRH2ZvBcRP01JEVjChH4jdcX
yeKRC8uZlJoFzC75nLLWLcdxFeNAAp2R3JTAg6wJiw91kmo+Pb09aXihGDtdA1OgP9maFh1/Z4pe
orDVrYylqYYHsMYgSPfNk6/1SlEitFeizLHPwSIUdIbUxY5h7EXFyH7x3JkbXwjcmgofsQNjwbA5
KgunLHwcXYQpyedUdi53b45+nW5vsdzNVd6rnvx7TuvNJ0iIP9XOFWztRD+ExV+Tl45jQYZBzE26
BEJu7bQEtQZO3K/DOyrVIeg2grswoIDG9HqZkryOigfvWdXUvoRSciXs7haBCtJYItf58w3GacFj
b4P5NVCZBomtazdG8533+w9nX3ktWi8wpS3k22+RbsDiLE2ZFyQpGXHacUf+DVdhLuxlNcFXmIaj
edNExvFKXVyLPTOGyl2ETLV0p7C/BYcrgyE8YgalNPIUc8NXbL7daKjrHBs8Z3g5qK7uKC+EKR6g
3R6NKExKo976xOAF9jI2HpfSls6s/8OBNfpdS2hLCfhx35OPLz/ME2TVIPzQC6BHKuYZbTqRiyG3
Ml66yaJsZ9yDU8uFMpV6cK62rDB7QfsCRxeXMZTGzin3z0sIPzC/e8LRk6iARDlRxtfMJbcKPYGz
MPGCHveVZLF1ct9hiozJfxJShnPGKC1vM4YF2JjudIW/RkzuC46lzG/SfyaUPDbXww8tLkkxCkOb
Jf6rFjKIhfAi37zoRMnPPYwSe+YTGDMVlJ7yEfgZXgKL04cTpwd2KlMH5bHixW62GSs1fp/ITUhb
ITQIMOOMHcZksWlpNw77pIF+2yomXWUnMh+MMW+jN+fssbo6zz4hNzK1JOPfB+mqtAPEg79jBVsB
oxlxG10D9flc/mCTRpCnLqQ2p+VwjOc7VNqamseMgUSPsySVXXE6BobA0JKgYbLKC1NFCLRHNpIS
bHjIn+hd5gUujeVov7wP9PaFbFBqqphRqN1aUkOtG81lWK3hcqqra1Q2tO/OewRvA4gilQOoyhLs
cHNoSipVESM9nRtRzmMZila78UI9k4OjSEjY6+R3xeJqxMFqPfeB65rOyZDHmSEtDV9eBaEBL7lT
NCY4p0cPT/Ji/De8cZBGai70IN1ibdzelUkfhxUjjslYQVLN5vcJQUi1ARy9RYOpZBOeXkbvrii1
JlgQDMlh9T/t3ErOtc8onZzvWPVkqmFYdhLa4Amt6Wf1Heh0TSBkgVAIkun+MYf5otBAenQM/+ZD
gHZnmuoP+VFIlJKsgdfHdFLydjj+jlBjKz2H5emnfpbxsOVQs97r9Mlpc3F7O3G77baiY39ZnCyg
5NNaMNwHph72fetWR+nHpcJBZK0J94Vl8LQAtJwx7LzRDXzUwdTEonGXuyUSh5aHE0sVdzcT3n6a
wIZhf7cOfSfvCcWKHWT3mYhFNqBwa+Av0PsddP3mlmeLvyNggQFJ5sefdldpMXIrexVDChLquAc4
oDP1fSv/XzuGxASM//glKGcqKwiq5bfxhxkvHwA9RLKMPJfHFJ98CjyZpFc74UiILNx+/O6UJRhU
dLJrhgF7Q4lW9KUBJJOZen1q+oPb7IApkMVb8XbWIVlhoh89OzNSEEqIZBu81XlK2jsLHiRX9VP6
o/Qy7514Tnei7OicyvmfVXIi17OdrghtecHq1Do4sm2RmxH6nahc8+24oCz9p34bR2OUCM+zBB1q
R+Tg9okB52V0wtukwKHDIXEaidaFl6QGBsE2Ti6SrlenCbpg0w0GGoakd9UIx7lgZG/vKeWD3MOQ
QZSlGk6zCyvcQasdgECGmOEcI+GcgArVwrKbRWhBQsI4fulkf1uoN9V/6+aBzr1YVStiqk3SBNz5
gBi7fjNVhGY+HK87kLp1Terqg6re4xPYX2DWdrtc50BJOeXpNcjDVEmFIquoEYnyPRaKMLf2hpi5
trjT6CI5UhzfMU7hjK7y2mv2GD23tQ02H4JYENZuGSjXJxmPVm58OsQvMfHygrbRTo4VisF2FhZY
Y0T8oq3UL+oevzekD80P4khpNkGFUpItM/5lIcBT+Wv2xJYk+Z8DAjHwQRCQN4igL5u5ZlJoOCtV
6ozhzQpVvZgoG0xcNdaoiOcdgJExGQofK9I0xvSbdqhFr6cwBqW83FyNIJRhMiHTugUx0ZmICRXN
cY+dh0uc98sFl+0UH8nDj7wJepWq7qbC0L9CwREvUcTRw4yaBXmTBU1gmOih3rLKauEWcaLIA6d3
6pXFGqhTZ0IFw7vUz3HBqOHdQq3wrNy2uv28GJymr0b+WFaJCmeUxKyZuQSqIofOZsU0AAlgJVoK
Cu9SqNezRm2d/L7ydRKLnceiVC1/cvHoMFby0J33grp74T1njvmU1l7m1+AlWmbJXzUrYO/D5qfY
Ns5bmxjpk+wnEx6HRMfWzO3XSZIxZGLvrJZtdwJBVXM47l8vM9TBDBa/XD8DD3m3EaW+xusWMA4O
YQTo9igfkVJ3hYyk4kbEwJ3/2QwISPmIZ0jUyVmvLH0+Fo0NGtGkToyGNdzM6GlhoO/T7PwDs0fy
XOWEaMTWei7Oiz0R56ZEqtCMGc1KiIs+mYuhWWz+wNKk2Fwg2d9r/DNVWtpVsyKUFOIEqYE2bUu+
h4uBiR9ypeysJmtAAOdZfrv/CVXn7OiBOsVyEnz9mrPrHu1XoLiI57iU1sasFNPKY1NXcAhmT1bq
447yjt6c8RVXkpgLUducCCgksq3rU8axrurAZYpU5q8PbbAqneajcZ/Z8x5HHptYTl7vz2vD7HAu
tmHKmQ4hZQJJMeBsp0iOHRcTXebXc+UBooJTqqvON+lUsihwZdauhvBAb2BsF5eqBO+Fhy8S786r
30uWK7Iy4+uqVT1RP8jtRCsGlWvyc1aoTR/thj/RFlBAqmt5IL9Nm6yGRZq+HNLjthmaJ/BFwLSh
E1LNis91vdhEETnQpMcZBZuwekp/8uKn+Mn75ZA/XQBSjti4VIbrYJd/xWhaGsg63JpXFcBYPo9Z
aXpgk61y21Y4ao7LeGhqLE3QGWzuZhmSTV084QoWNfyXBiRHq1dNDk18Y8eVYEfHJ6+gG43WDmOG
4sFftoNAZ7qwD217peySQNeEVPsPV52vhJd+tROn+cNV2+wGCC2J8pREjDHHLaFQqjRt9d0XNlVw
r1PUS34/EpZe96FVwZ2klLEOwE9i2p3lW7DmpGBYtEUyJ1mOx96TdA4ou3kJYSwZd7siz4yMqjTS
OvMFxoKc76Mmdmqcvm2incTr4wLCOtkgfR3e7zaAEdjDOPY6bXAXvpqUH9NNMiYPqmTAggKoi2vQ
13wyGwFqnAuu0trgzldN4+xT80g0eYTduNxB+/TXinFxhu2izWdwwIB5gUvcyc0LxBaUgZf3Jy63
q/PkpwMryE8bnx2zUaS0IPHZzaAEJ7zfv65J8gSS+Zz987FQQKKZyDqosfQELx3AmYTAQW2x0mAw
H6RQ8ugOjIYbrECPn/RkqfTdmMxWls/FH9OiU/eDRsoizhsCGNHqP8CC5+l0KE2S/3yTRowfX7Dg
lnWfCpV52hUFCHE1g2X7egZObwjEGlMGKiKbXOsorsl4NjD6oHqjB/hNem6dzZcC6hD/vYAjqsh9
aW49G0EKQG5VylHmAiiYeunKAO0VG7p+7EdQ4MtzJ7BkiDZzcOfTVDwAJYTgyh1g9TU3wK10zq2o
QLXq3j6QSoaZaJzOKj+7ESbIgNi5VEsoXGYFIuHDEz9lSPschljzioN/xEln/EJfY+dOZpNgIzf5
2qH3CNacT407HQeN5RjXuyiE9i2zAWKvtoQ4nJcBSJINZep7JTzDGDqWTVdnj+gVIiQ17o/CryvS
L/SAiud+wnsDCHgQD5/5LFOlI3PuHhflYEg0NFklGk7Vzqbzfb9FDbSt3fAJSEn/K0sh1UjTiOZW
gN1eahqqGtAbAblTUP1OyEAsNbklCemzhe9t1b6e0bWBlhp01SgDXMj8PGkXvP3mH7gl+8cjipIl
z7+YgZFFQq1jHKSYqOufGMXA7kZzG3t6tv9IOU++wrbaSwuJ7cv3xmeeq+Vq6SI+FE1SIeXrYWV8
qmKOtoE6cXbRrQ64LbEXhq7EJbMSl3WNNbryGEJj5bdp5v8iwalWvUwlMaEYWNrz0LdJg+S0y4ZK
SfxwZE+LX4SIgBQkP+8LtNVL0jh1J4iUShkxxPdrWFiBWKHI3lhypz3n4kMvviSwG74prrMSp4FU
wdGTNY99UPa6O3weJ1TRIegf+8T8qrYo3MQbPJ/EM/3gH2n4ils61IiGUSbvW49XQG+9Bscj1Qht
eGgWLKDs57crR0vZUCcShqZpGnN3sKsLPcsalx1vIn/0imOaSUgHBq5JxpD1BHiosDfQPQg28h8H
//cwVu5tc43gmiXDQugmvx2ROHsojIIAL04eQLioCTAlN2dvyq6yJ5OGRoDcO55P9mHyQL1QenYf
PgfN/8HZ3r/Hjryin3mJp5yedRUNq6TMFm+8psMKvqxZM/FxONwgvi/qEY56gwJ6jySfI+16g5oP
qabovBTdBTVpuj7Fz+OC4CZbGJ2a7vcWma+VwJLzAnqzUqYU/jTdazsegtwUQ8rxiaa+JKksDt5p
49lVMWDq+5bYrEZEjve8KmduLdEUhl0JnNh/1FXNedwS1fI+1P+WucgHyulrLtqEm7l1uneDHoOD
uSFalDdwW2T6fRi6ZB5IAmY9eiXgN+ogJdWmp3AHo09/N3Oo3/RfSzqrJj9TTdKTnaPkjtRjZ0qa
j2t5CKFXIAO7VGmXxbMT6WH8e/Hr8/M0Gprq2sK+o1P7oAuglhA6TtH+NPs70HAiVY+xRorqPt59
Wny1EnoPwyoxrhKqwYH/fKr5Lomg/5E9k2JMQZSb2NHAu2nTIWpVnamAzXKxugYf22O8oaDK0g5J
rS/j8XSdBTXo0LnqoafNRIKNuFw90X3MgxWyopo74WcTLKp59w8fA4K/Qxbv6BQfI8CNkp+KkPIA
OE5mfJL14VnC+hS51CxaQiXfv5SSP2MfeCa4Gx49KIDmPipwo9wOShbBdPk5APEBIcnGjhJ+DZ0h
ls7h6AvNntf71Dn1fD1V4smYJ5qXhotCKpRilI7xFBtSM0LUlgZhzErqG8sJDpZIR6ag1uMurEka
8pdtYm+lxxzGwhLB4NPIel3546YXrBxo5B0Iq8C/MLXeweJB+szIKWnwS/TWZVmZkIeKugva1UNV
rHEzUirK1XF7JKHENk9iOb6rj1dAsVfhkXE/o8xh2NJuC7J2uJNpo7Xw5pXWdR/uiJcy1B2NPjl6
KUkMpLYF91x447jecJ3yPj70WyAELUz1F3aDZVpu9SydwMdG63VBC3Dz5hfnb5q+IDpch/kfNyFP
QJTHMynOGsrqw/eM1Q1857i8ATnYZ5GWr2V68xjPwSy1WRHK7dITpvO/hcXSlVDiCGUqcip8Zt7v
mZjLX1m0APEVHxc0A9Vacg1TOKCCDaXeOxYa9owfANCWa6MGrwYOjE6ayMj9S594aaif/jO4R8yw
fSF5QAUniGw4jk0AVzOHkOF++5GqYHQX1hkMpRWU2q5sm6DmMSNd9WRVToAlwv4uSSwGgOx6uwjn
+Y+6uxvpO2T7CUvTHR07MIrPlh1PxJp/HDFGbuln3GipfD8DcCIYXP1wjGqqm1PlwHr8rbEAxjBs
/yciKTjvHbX48KIyLl3XziodQeq1kplzmWfSgMjXufRlxwmk3Lg7CHOeGNmJ42A6U/USaxj1g5z2
P7F3OUDEQ3x96S5ldH6bQOs4tuapirEgaoMNuuxUKM0gxozRnQbXIulPl9P9QOdDokRBGiI9YdTw
FAjJ10x9lFAWVgmS056SCrcZJf6UWyA1VsqMlfvJslZzjSS1C7tnW5/Y46oXWhKOIeH9FqqB21zM
G7t8UWk+P8tsO0lOLNKyU+DXOhGYd+r64snLqbqvV4KCKHYgkA/OrijPFCxNG/G8FgE59oBbg2d7
sNMqUuuEMZWjAMcC5U37xkD11o4IBtIpAgnkZFdL5UhjlRauulYs+VH/LzocM/p04AkACD2kPz2z
/wP9jxNH2rwqrcFHz0fSOprnFfT0QoEB5ubh/8xR8TrsaTyqoKAu3CjpDkf+em2/ozKeXvYudrnD
lUJxhvvkkLLDpmpqkJHC18MvsQDQctMKhcIGYBNV4xGtYH4Lu7E89shxVZJsOm8Lqo6CQXV28ISN
4h8uc260TQOFK32p/Ng8gwEBD7+ynBTtasbC5upaJijYfOfpTMooQRw+p7lvPFUvd9Q5FWMgdBNM
Zstet1TXdh0cfU4n/LOKJoO3oQ+Jkt3JUQqLnh2TdyXo66R3I27sA/JtLe3CZlNeiXbsLcPcMjV5
AQ1BT3+vV3BsPjE/7jt8aTm6cgr/pjX/F84RZHysXJwdRuL89KWUg3GyiN898p4toO7ac76M2u6W
S5i7OahnZMiRzYWx3goezgCiUb6CS6wD2jwu18eYaxLycOf7jEkmZBjixig16823KXZf75z/SVgf
NbU7Q6+NciPi/eh1lS1iGgTMFSNIvZ/z75oKvG27WiEJ4tOA/787H5eHNIdIrkFCW2dkmTZk0i40
AkkWoDKHg3sYtzPGVNoqDlPNh7uIAyuwOVw/6v1PUOtRcs6ZeC+C/a5n465bulzf078y0DQD91eY
5bR8Qa2TrdUyua4XmlNVpXmQLtl0gt+uFKPhO6Nr3SP57PYdMN1sxPt6wgWepoCZ++c0qyPCgwqc
3k229NWsZFicu9ZRBz9l0AVZgQF/Dnbl6xvtoqGC+yqfGJDS1NNKorhBG2htphU87VXiztD7xsrS
4tdvGbceG3S5A1dykZmq5dGIXjAXDc6oagbq59+KkoPmUHqE5hEmHI1ve2Yle9dlvsz95eauF81c
rfBqt3gXgM3r4f9rLvcT8mduzR47mvVEIKZAqYuOWRJYJJ851s2aZmyQxCamjLrkYify6WJapub8
E0/fw/HsUoSHZH+uoflMucxqR2Ewroek+Y0lJ6VPcdpcfu8s6FdrJAGq7dgeC8COX9SlpahUmMOj
4RigY8KzD8QNEfK2yvtLIsY04keaLd/TsNFDij3rW8E8HKGeBMZD0Yx2fn90274lAFkLnx2f+d9d
M2HQDraKqOlrsoLI5hV6aArW3kw10NZgDnJZsBvBOyYILpU7fXiqFbdIq4tCQRStQ2izJAJ64tj2
0kePkNanSNPw4gYdAk6U3lgZ4W7cf2wLzMDO0SJOSWRseqkvZOriOrEAp8bXezi2ptKxHvPuxO8l
GCm4roJTOKne7iTJjnszlc2iYNyxJPtC3fk862/STtT9wUK87TCZWqjlau7FRtAqvgJLM7OhCmGx
FPRjv9eYpFHLvTn2ELXLu29M5bPWrQEmIER2RR55b6xcS7BgpZnaidRfh0r9XoKQf3kNhgOshERm
ZgWCw69Ub+1NwCwZJDQlVC7K/rxEZJW+pP7txKgruN3AfoVUWl3r1bfW4cTg7bibmmeNBatstaMd
ld72Xj1fsoAk+l7kgzgEH6o3+tzv93tTW9ZGlqxPS1eA/HhPLjjhkXIlf38UwLrGZNtZDV/uBHqW
n+si2Hpt/n0MCBhgab4OEKDl4I0wAv3Qug5YS+wKiukD9w3YpIyK9RQCf5BHJtdtCoNS2OhtDdCp
RHSep7OYSWfK820UnniW4483ezkluhivSMzYKeIvB8t0PzJ1giW5kHvxnkQz2j6vxdbXGi8ne3gp
msYN99wCAlknm01cCZ1UEDDj1kSUCecud7y14e3IR5FGR+8DnhGT8BxQ6WQqyQG50HjvDt2STjqD
G+itWdnyzMp9QLxHr7NUZ1dWdouOPFCddVmXrdPsuv6dY2h8vorpSiggl//UHp+XvJmWmkZz1R0a
HViKmdepvvywWwKQx+6nQul1zho6un4ngZqPtL2GkcZPc7ysBm9bV3dL/OZ9swWXs9RFZB67PlRt
fcGxSMUhoPHSTVVrIpvpAwp7BHz20bwQPh6lfH6j1D599tvleS0Z6N20ZeROa2BMxOAWCuz2Xa6L
MR1teHYF0KKd7SFX/tqjwU9dgr7fUKXkdSVH4jhqJ6KIv2m6DIQRVjw0Wh95LJKYiMppqzWAuwSJ
yPimx8mFgxixlLXa2LNxPCtAJB96/nBObKAoxHqh3eVvFibcRFCLUl/RCVyrGyjmsfJP0YY6dt/I
4ZlRbCLMjDJvaIjaKgftQj0aA23GFRWPwEZEnNz6KkuxTwJhi7R/IA0FpOhD+euqOIObD52Ll50r
ysvTHA0t+CRbuhoQJTfQHELlHz/gc2g+zeAF08wa+EhpXHRu2h8CFc+NxYlU8srm1uN+pEivv81W
Lnh0Q2A8cTtBbzX4Abrw7ZXFM6eCduIPraoIFQWjBQCAKqvrVhlBcXRkEtxzxx9mMtIoz18cWFc2
24suHbqk3Q3kxl8FnKAImOrNHLDLnDWU/S2oxCcuMfqQrX8iy+V5cFnmAPTLXDRUQU5CgKNx6rWj
3cc7oodI6atEIFCTgcJf+kGmjDzEpbmeGHOuAuw8PT4uGjKqx+GlCj7gx/GihP/u5xsFixf7cKAd
sQ+PTqbvTTtrBsRBkA3iaT5jqRn+N+RlIf7U0ERIl0mFDRwM8kzQVrmDsX5PoJAGFsLYv6tERAQC
Bt3Ry/DW2cXnaP/eHBcW0s2loBEFqXpiHzuu0urPoPNNudqQ5v47Gjb4m0b8hi5uPmsZ7OjjVbTu
qSACtNTu50Lt5+DYnxCAjt3H7k3jj4UUkFaGWPz4/7PPfAo4BuH5qWAc5p54J813LiueZuhenzkr
jOGfIajKsaJqIQGQtvhaESqDdOs8XM8v8eO75e+W6i9si6oXLlyvpH0Zji7QJVm1PO/oqGTCBo5d
ECPhAhljMIJeP0yruFDE/VIznEVDUhg8EGHNu1OBr/wf7VeqxnKcQ5hf7lhQp+CMiuEleTGvuM9B
13pFR7uJ5v+VbpPderCFTBwkTKpGllUnLIO5PtOI80TlHNsqxt8IxESYTCHM6WEKPbHPj1s12WUG
82b66QYDHztgWmrBpPn0x8iCjFSA/uaR97qa+CB+t3omVzvoCu5nqZcB6Im/pF6vEOFkOJoq/ytQ
QzIbkO0nbqaMSiHhYkoAHfxXKF58PQmAJKx9jr5P4sLfdAOmmmFqZZ+C4PMJcdIROLGXKZmk/bUZ
rfQM8Zh1v0rspegK44Fkdmf4NvpQvFceJkyTbtZ2NRuNzvzYZxwMl10cMKFSW5GkF37Xv7jB7p4H
6MWL743LYIG2CdmF+wBKTIAIobd/8bvl0BldotKOWSQ1lBWI0C1Z7BBavrPU4SEaRK7MrsnzaGkB
4ScW9cOLEqik658v7b0pb98TAenG2z5gkAWHGmQtBXquYPRipiNrJfhGpPccZ4swfX2yME8Atsgv
NW6IKKq8ehLse2Z8+DGvHVh0b1bsq4oTWwWujNlv1hA2OR8T+SzeV2ii5m9nFLk5qFl9+KDohTW+
fSMAekLxw1PB8wHfXcm17P+utejPmTeNYUiRdl2GH25UgFqIGg3iFTfx55e7M7nQKj3JnmKRgbbf
8xCnkWSSx38/H5tEl9RmCxWTIps/3ZKYIt8Q2LyGCaZSSp1G8PEaYMkZ450nh9gdx06+ORBJewgg
PvaquPqr9BuUNbHOSyH1SGrqhysEcrSdvI8/oq5NiGw9qY/6ibSubbF2vthwKGXSJ3RM7kBxjz8K
1TuUWFBUsFQ+jb7uU1FSwliqWjYAeyKH9bRPEOgUmpR7Ghktm6X22mpZ3fUujKKidyXdlYjDrWkR
ydbgPWX/ti/+AbVko6pi/QZP2OuW4UuEbWreMP9QPhyjdf+ksmiO6egosu/SmW/hxcl3SLc30H/Y
bR/eNrp9TyuuCyECbYbApDtFUKkMaAFZ5bPMNE2YAnvaPTk/JWMaBdl3b9GfL1d3s04ljBO8yg1b
zPqKbxc861XWq1KArUXYJprF54kODgfy3di5M+0gguzjv51iFsOT6+WUbKYxYLMi8Dn/JuuLuWD3
sXEYob4KN5AS12NyqtLQTOUGODQC4/TnJozAJnAb7Zz4F9wuSH8/s/kmW5A29Ja4FSsmDPb8jFY6
/yTv+WXSm4bsC7w3idEUJ6A7k3If0KFhbE6Kk6gXSEAph9g4+ZepA82BT5tGdZYmSLkBFrNxY8yF
3KOduwa9Wi//8vEhGxHPmp+kMJ6O/7RZCOPvadnFE5bqSBhKqw9uX8J5pCr0PAQ3irCQQPneqeWr
gjF7yLuo3HDlk24MSSwkIjq8vbP+DyBJixlH8h5lEbOnKVDF7HakZw2fLamnDhG/tsUQ8OQsjrLp
KoVEjntnXdLR+kRGBO7InHkJfAx1aUFPZ09dZnjsJDDNs7oR5PipGenGS773BK4DykRw2UIpqTRI
sVG/4eFnZ9VBlVYhoC0AsmZKBeZSIO12JAErVJFJ/rPtdDINyxpnSOcVqSMxkpeK9csqu2escN9K
7fxjRSVUXYOjgdwVuC/tU5SyoAA0MrRG+jjLxiauNXICEFI+wxgm1AAq3hGz8TgJBdF5EZWVN1Jg
ynminHg/RDGfz/u9hqbBO6ma9ruZoyqZLVxaKCb61hTbk9BSzjwBLcAdHohjtwXfwzDi8whV0403
DRpp6/IYGk14QC0SCDbseVScG+5FnV/uD7WgAtsSr8bgq0YKGHI0/jKAklgXCvjsGIEzxibdni4V
zK5HfhoyjRb4+PtyqJeoBPcjDDNPRiDVrwfF1C7QtOl26WoHasS6fYjvt0o0HbjYGrMCFEzJqF8V
qwcdTDwwSd5puCkFWSEU9WNYP7CzgrV32EV0oH8w5/FbRx2aJiIm+8r8pGK8KDLctGykLn56gFV8
OYuZQ1yAFIobqIH5uB7M3sRxXACDwvZbhLMDZUbo2z2wSAr4SgL+l4P1QexGokyYE10Gqr8b3Pez
LeMmeHo9LZzRx6eL/iNqG9SiupiBVdZ8kNjzb9/6xciNvx+VGYEcNfttjcSBgT/DYMUpN+k593ua
MoQnvBwylbYL7kvDmyu4hF22ffp5ps4CKWz1UbBpb51QzwuODij1uD1RgxpYLd/TOaxiruUpPzyY
OhjK6fsv2/I+PWa8P5bvq4BBTt8jhY1xmEnezT1PRFscsbeUm16lx5N7rzx3W0Bu0WLuImmeINNp
AWy6Vi9Ky10+4Eck+AClHm56lUJH/vyeCecWZSKJ7EAgDGRJR6oAkeMD5m8ksjE8m2jdos1FfZQU
VC+JoaILNSMIOLUXyzKv20C6A/5SFEZG2h+thK5QJccL3wEBBjCAgPdzgMtKuNzGOZAnejPB3r3r
3SVEc+it5KT5dhT91KAG1ifk+HBmjPiftrJ5LGyQHpSylwwQ4a0Cg75ZgVOkhhAdt7/Ekpp/1ajp
shuBC+h38gVMDYeS+HjISsEWoe+WzPX+GlS7aG5o8wJN9N63+8uXMwLWxC8LrV5bh5EETWnFofeJ
UKBNGs7GadnU7wMwGGyNU+szBhaAsL60ELQ/HgZKg405V/fIErfUvW6WDv1mxgk18sbuVWclqh1O
W8aDy5wAskLgAZPr3lzR64qNxlhhUMVspOXr1t6AWWlNN8nIVjNpJUrveqj8Pf9JtHGpJLzSt1A0
5N4MCwhk36PKjLA5sel9iD+NHVRT9f1fY/kkPs9S2ejM6Q8gJd+cXq6qgCydypfpBwdb/EonCaiD
uXxWWOGsBYzj0sCQNxnttoWlEnVJrl4xMuX5iTvyib0ur/w0CZ0Ij85fmGH0SUrKRidL7EtQYdJR
HqkCT17bN+87+Fb9gWL1iOV3zV8gYfHN8YNM6hX2wZ6n07UeFybZHi2cMR+4HTV3TlDREFYl/hO/
f2jxX33GOxkwjFApdLDkZDm+ZLE3uix+N8Urb2PAV0byZ9W5C9dq3rYgELNq3ySzMmnt0ZOaI/Ng
qADXv1T0EWmcvzZz591q8KumYxAf2nkjZB3QTbnlvKdsZ9gm6kfP3+1IQmf1ht4mAwF5Zpxi31gD
wc6OLwY5iKjGm8ZTAcR7fPEeyd2mDALlyfSrh8gDR/Ru4Vy7Cq/K81gNylzUcuENk1ZVihUxjL2Z
WFe1mfzDkRgW1e7U7JCbq+TzXRjGRO1u3DkIXwMEM1kXAxTMPYtutkzpZJxGGe3GhARU+FEGHyhO
SD65SV+CYNejDLow+kJd8KsuHI7gaN8qknwh93pnqcxU3BOo08F8AFbHkJvQPtdK/hamHqQfMFrg
vKvq9GydYxJaUkAzCLwiTLYUWG4p3pBFNNrVIvDySo1raTp4MBFQjLQ1ONqHG113GhYp57Qe6b5q
m/vT52Q1Y/d5nQoiknTBh5QZAa6EW6Yn4DU6UAMlUiP88SqOf08pgNCoUIebiQmTV2kTOl7GVioO
fg58owquGXlLRNZsiQ4uQhnVjFmYXBFyZ03rpJfUhl65ViJSFi/yjui/74OR6s9a9umQaUNSz4r4
+jZsxUdCk0+HKu5oWBfALtW/zfVkPo27ARR37aqw9lKw+t66pC/9Vo1WyOcWtK+vLjTtURrx/D+n
JZjFW+2XgFBEjpk1dC1eU7XKjrwLqb73Xo+zcXntdD15EYiCd4VuqhZzz0FzI+vqreG6BEKH3net
FRD2Z+PYaTMx2G3BgogK1fO25lzaG0p1U2Z8kf3lk2ntHxlTEvg16PhyQokMvgwaFNC1f1EFclnW
iFn6f3DvG3KFe8vC1ihkhGk3OO0MgEgSMSXBNmyoUPSpHyKAILukB/1D5cszDWb1qqGQWSJ9Hh1U
btk6v/FxEVtkbJGzJUlDnsNg04N2MG1eeCDXv2yQ69kYKx3+Eam4tWINwRENdAs/834I0MkQJpol
gKY1NhJ21ofRjV/u1yDqUtkpsX/X8SshQJg1j4pXzobiNmgju8fbnqd38Tf+o72sstVkT5UrUqII
CgLy9FFPYvzagenvrekOOp/CeOqgFeHgWA3a3+MsKYH7TJxiz3YaElHfMRxdLQxtk7sF8DjtAU/x
bnLMtNL6wplJTLyvjM4nIAMfTGCaoR0uGbYYyA0UCKEQ3fb6WgYs270j+oxUGKdsnMsirLvQujYQ
Dcm3kwpCoCExVvGGyfuNsWwh3sWNMgRpsFh+OPgZXBfTBkJYd+wO+VEGUGYNhp26BvlkDwY9EaV+
L9EihN+HkEAuteHm5EVbGQRCfVUltvsOx+2RpvpYmcuJsbKxYpxh5rgnDOIqvSvqxZLucLHbnJaU
S7qQY7KvikGB7aZzoEZDcZbSgGblCNeghAmNVz04aSXW6MlC0sttpgpyJkexRyxtLVGy1nUH+qhD
CN6+Bwtin8czUf5GmKcLUlBjeXNOVW3j/rZ1nlHY23TQz9KmCylPPXz6+ex6NgZIeuM5eJlKjFgV
gV10bZHEX2VN032Lh7EfK1RLR8f1aFkXnHXuodOSFtgp6lL22gyurWM+o0ZUDc3ixgzmQ4HfuHdg
Q/FLTwKhrGic5BaoNfWXk2ZEMJox/5rV1WZr+KHTZFO/i4rbD1QC3Jy06qaN5052VbkUUCh8e51E
IJYUGYtSbng75zXNBo6w7BmCpz2FuVqpjOxGFQo+a5VDRVS73ZLde6iXlBc/Kze7blF2lioJHSYi
RvG47u+LQ9epyNB87+hc+fhA6eC4Ojz0W60K5rNfH1QMt20Y7EoG+uwTn9Tm5c/gtnxIsQfRvL0+
On2ArSF/AxiXMVCfiXXyzJXYAVLWi5eRWdolYqa/3gKc8PN8fzUiqQtmhM/OMb74z4Si8I4EPb2L
BQ04x1I5FFMG509RrWKviCz250kh9M0KDUdTk1yQM43a6XiWAI+m2BPKyYSpnJF53VWGmyZy6bcG
CcSrRKiIlZ+FCqMEweQG805eJ7ER2r++d1htJhzXCtLD/2M00aGXQup5iqn7D9tWgLO3Ai8P1pm+
BDmyywXFYRkwVnSBgtsUlLQWLUKrm9Q0KmW87qjg7VRriQSw5BY5TTZu751w+BjAOhumMo/JebMe
+HAO1p4vigU4cZPmq9HClmngaKiAlOPfyJsgK68PdfI/eVWzdmolvZMkDE5yEpNYnwkIOUbw2hFn
3b5dUVzvEk5Z+VneGV1BLPD9BCcCrzXeYtuu6hzqnz9IyrZkwplhGYWYwq1+ByvMlruz/OzMZ1lA
GUl0WP3OMToV0+zIONLJOgwR9PaPgO902SGGfAqi1wTwoGmvVCoxd2OWQX78SMCibXrqRsj22Dfy
QBBEVmKR1NBGtsxVLhZr2wjiEEzWwSdd+3ySXd9Qriet0bQQzclZaWzlaf8DoUrQ0Qpdo08UKsv8
qQh1EcZt59zGz44F5lPtvW5ocFdH0JQVmECPE3OAa4YlUnspJCqfhXZYPKvKUxW6aOKC9hA2YulK
zgYO01MhHc4eAeluHNrQfvwTnhYr1xo/g3uGyh/pIZtK8sSoGZTJ3NM15tqQAeSDtGnekokaet+q
SPX6Z4w9iFfpR+2xwSdWAfpByuSO7dgD8J0zT9OORZ1T6ZH9P9a9KA8dEP3HMQRLmfzFux83d/iH
0qfZxnLuy+WY0/QDywewWUtxjRVJgThwEeVyNmcnAfD4JpWy598e9DdUvgSoMJv0gA2g80wFbGEq
x/xjbWKgrBLP+Q3VBe+nJaRd6fF9ubPwxGGFKlQ5TJPr+i/cMhX+DMbfI81OsLXQDA/O3/Wsvbuy
DfJeIdyLwY5gO9BhrmhFFAb3fny4waaF1KuRMuCPQ0yWkNHVHaVnywbXgAdIXKUplRrU6vcd9k5d
U0ClJ/CYD680gPDRdslbF/dyqz8UOGJ/EfgTHcoQ6An+BJ/dmz784NHzo9okoKOx6Y/FIROarD/k
KO65Lzqc+Qq3vmQr8P6Odl9KLqFpAxSRjwM7/7PSkKY1mxV1Qn8VWJ8COt2GrDLNYoAz0h7DYzOF
9+3Z2MfO4lKZ/RmWkl7pS01arWSnf9UgOy2c0Vg6us38MyqhRKlFJTlXwMRgfvrDaXQOpG/g94eX
WO5ZzQV994hCY3ReLP5G8Laizv+K/D/cpJfyTW8+ADK/c/IxWFTJFXCD8GMkgXCiJCnTt/d8lSvY
lI99e5dELL993X7JaimNGWor7fEBT1VhsCh2UKnvvwAC2NcV91rVGY+uzMapOTyzxV2aUj+83FiO
aENGqu5sbxqze9DD2UMQa8FwVgRGjXrBO2zzEXJOfK8KBfHX5niMLbXwEbkoCO/XOvL2FpGzvwEC
kinUqnrZM3psK+RYEWFVJf/jwEoa0PI9oioJxYiH00s063onZF6aJfKYSc0p2/BXslpfz1Yuh9oY
tkbOwzmY0GdtSJFdJy1EOZoEmfC0w/1JFdhR70QkcIQbN0KLU3jzq2t/A36CGJFt5LOW0va/hJe/
w/TgOVtf4XIKo83zK+oOLR9emWYAH2BIBJgFP/XhJpO4gciXYmMqhZRaYhgE0PinHGulpDxrBa/X
Pq1UqoZsggbjSrIGhA4SuLgPVLp7OPArGlGaICoWw3n4bGxqJMjggkYVXpAwHdnqH1ZJ9eH3ciqT
u1gZUBTgetrwFMsq9PHRRRCFi+/80/jxmyQNFw7rPNToeO6dRxEToWOj/33BTgp3BHNGCbqIkTbB
+E2V8dgtOg+wdFtAmE5xB2f0ATF7LJoiuist0pNDQpPZ9aSTQTq2i1OQhW1ZFeL3WU/ZxsaAc3S0
zqzwLYC7qDtfsmb95a01YhF6qRZRsnuJHAc1h4XlgHf6FT9w3R8oZueFHL8pS2kWMZktJuYhOGvF
t+mqDQnad1h+8DsM776Fec7auuipsVMrjQ87QtJyfyEJdyuifP6AICVeEz5IZsPR0WTh9f4FzTvF
BeKoyuTVQuS8YejlYBBkQyUtEOQrBzz94B7i9/++6wORGJYLag1LpeELNPXymBH6hg2NlnCb+FCv
gNDnuHGTGXritlRSDxBzJEv/Cpjs8zK7UzfMA1wzrM3oHzRMxOmiorF6zWsASGfN/oCG88HJEqxH
+C0QMi1P0q0L/TOxa/c0+ESrjbwFu/YHQUpPRuJMVkmCnqxcaJIdZSgWK7boaFz00VJ82yiZWhB/
7Abd6KL+DYa6wyFKeUYXrlzNnG6VcmEi39E1alv4SYaSgbkV2TS04oEf9NIhinl7hcxm1fHJ/iPn
9+qWlywSDR79PpJ7txcJ5+U/PbYdj9NemoFt7rkKqP3AnFuZKBU33WgsfgjKSA1O9aUWHxl1yjk+
P66pvinbrOMQiv9K7NGGPMrN8ExSsJX5/qv5JPRfOFS4zCt1OD2wv6R6PavuBguH15+9nRNeHVJ2
v3qjx8k0bMXmGx2/NqMpzTUawxR+SSaZQ72zZrPqGk2hJCsex+Y7VJ/cSBk0NVkoDGyhsrWMdUw6
40w1Z4GDDCK5PQWRI7H4GODAHfcY05+FOqbhIq7u2ZXZc2QNQQzvlzH5jjRrPMZhVz976/mmHCFE
ao5kpYs1n05HR2N12YRbDllg3KFiYNwUKHscevVgHWYxBg6N0kkOEJmM7ca2G49ENJkWFeeFRFc8
C7dVf5FfV5pzM7f4Y/qhmHnT79LMaGVLHBN833yVYPtB5Bxv69veoE2eIHj8zyTW83RdnFriE347
jO8c247ZAMxwwXy3HI8+B9IlaLRUjK8n90lc2lY1zOhfumQElycFo/O+Uu+5qsLnYWEi9+Lo8NAg
/q8H5cTiStcxylbapktyldv9tBQ0t5i9ZwX6oRf2y9xyWO3qnggFxFassN2tWopI6/ELmOOieFs9
yj+h8S8SjX0YSicTqoMMgmxNWtnKsYryHxWEKJees4q1UfoZvBRpyhTg6zBTOVqCfDtb4cD11A1P
XMqxnDLk0F2oho92BD0z1T7Qgdkt1ualW5pP6T3zP4WudUHC9DUt4l3d/Oasuc5Raz02QU/izead
u/8faH5mBLKhhJp7spsv8XbWyRCs9l6Xse6WntcIZ+KolVxDUaNDv17/CJmv6fvMVLPDSpdA8DT9
v+HObWQHO1Y1kFrlqbnhrB7jINHd0cUknxwvqJFJWuUagGWHXUTawXveAWE9HwpWHZv5Muz1WYMs
lIMAQrT57xg09hW/ZNdCznlRIVRUnpx3RDMLoY5kH/pdAfGm42UpCDO8lOS6o/B6q7jYNOkQPdFH
s9vmbRyxotdG7T4BTLTigrOVeh8iN4LOY1uQbT1s1W5r6IVxkad4Pr382F57RyWw6YbNBSh0nN4j
PCUQ+gnvisE317TCuJS462ABt1gnatVvpwltxukmJ9BuGV22FLTYFSXeVbNSWcWXN04aBMM3KNcR
EGp+cKjawDxvbz1lbwlYs73k0HiCdYw9dj/jx/DrL4r6wl0FdwR63Ja93udNvdDU7Kj4rs2FBmpB
1/ALVUp2QJ5/XaHL2IYQOU86hvtKPTdH6qA6FJLgc6Dxyy8y7x8cCsARXs1ObTiji6TXN2YN5EY3
omP6kJRwG6HlQtzOechWh7eoUDiIfqxJGpJnSFMmz005BQWOz/ktR+4vawEf5ojlmRjWK7hCuyYH
oRgLInOE8dR+j0ra1c9skHA4zMCe2mf8RhxtDg+8emkyvUSmTNufirqFLgJKZv6abOC533UNqCZl
C1KzoqipWl1e0lzR70ThWer2JgFV+mqaqhrEFWqCPiGpv3dFkiEcIAGG8Y1BIKLZftM6lGTUz7ks
2HX+TVQ/7NF6Y8T5RpS5617Bf5QiRoS22uS4JaxXL9o8taFpLQEVuiTHL9dWHeJiRCxL2CMNr7cl
Nj+MMfYKdnBxYrfOCQtx82t+/hBcrF6pJiZLeE1kND8lqqs9gakc3Tghv++TQolWVou01jO6isuX
ro33cJQwCAir2Ae7Dsco5qSMJZbC6z0u/VMMmjGHRyLFxDtsqzSw40PepSN9RwAXWU48fvyWW6he
FBolfuDem8EbJOG7blj305EA+iYZ9cQIqvBMeFMmEbixwSqzn/woszwRYuFeJrveWkdk56qGFEAU
y22cUWItbv/RZUzo/Lzo9oqtCks2ruqWH4YBWTWoj4I2SJnV4HfTc7SULsszuSFF8MAaqq2Z+YUP
rmz5tl44Cht2So9IRMVYCk4AVoomBwvPeDITNYtZCKW3wiPQDr6mrFqJEc0ku3F0g0a79Tp7Tg2B
cABCszgPrUElOKZnbrTzhXD2USULJWBb7zQf+g83OuqFVlnbScis2wZX6Nkv4rer56yCT6xH3+zG
0y9ci+AlhKkhXx54PqB4njsj7rHNjGI0RlJ2wQLsrY5OhUTsSU4QiqMPVizxBeUrISmYTyCH9snn
+E8//OZ5sfnvUjLFRz1UA7Jv29A4hhKSCt/b9cDJozDC5/N6I3cm5ZvYtrGVWYmGH06xkixitEf1
77kYlFOGtZAGFnHKn3Kr2gJn4aU3APnb/sb2+AO3kmOYhpDs8eXX8hdaK9lMG9V+EtwPq70JuC45
1c3sTR8VrMyWZumh3yYN7xFdt2AVTboZ0AdMvM4ub+slMY2IKHPWtTSthXH31VAJ0FOEDaeCvFlt
TQTe0bNL2pSMuViN9oqL9vAf79IT90KkKPCEc7fUJ6TG8CW3Wy/TxqZ1sWRiq3g1fKy+xPejIi/Z
MIbpDmLmxnS5UQFckZkaSGxn8D4V5PB9OIl45neer2VAxJUSuyivARAdCdcJdouoQvbWrocjcipm
p0zjK+frxmhHtkd98FENst+Tgm9Kie41irEVeQN+kzQV7IwXAJkTQUsGgn4W93vSr9GvMTjEiiyQ
LFl1M3po4kJ0OanGsrBUgQFL4RHDvMNN9AvAk2iUgqK2AKJ9rbnFM48wvgONzje8lgxAUaR+837v
vyrkaBD0EFlp971xgZOcN1T/whtd7knMTKOINE4+qzqOKXaO4mZ8pEG8pcUWgvriIJY4rIcVQDSv
JWdvyUWrxVv9pyECqP6J09Gu7I1TcpWr/1OB3mjGDMV2fgkXuV+QJKQpxYHJl3hKvPT3MIkxS7Jh
Y6ASZLWOMqv2NK4lqkDY4/G6BFZ5G8HEyXUx3ojHY2npkqXwdJoyCZkArJWo01cwRUOrauZJ6Khp
V3OoEuYxhYT686qqNjtFsVkJ3rKvSLzxBENBsoNcEYcqIjBXl3NCMSISog9UsDwgbuXxrzXw7vm+
ne5hjOTDvV0SUa+0w/J4hQTqUUBY6UWZyl9b6jBySHMwIqL/jHDZtVolz2P+ouZBY81P1AR2DGak
bN2S+3tzDx5ceYxIbZruh9xGU/JKJO2YQksK6Oq2oGPDBlViHOYnJHNVcjvIZIBm0o65mC5lp1WA
0le8eE6q6GywF9lhKpKflinFSoOteXARBqv2gVaIXXGrLSu0korEshSoBWBvSMY4jNEqQ1wYdbR3
qtTeWgQBSwxbnTQ0wkTRIf3ApoyejKUzWqA/GsAaF+bgtwJIyT3pojZkl2pplExFmJjRnnJN+nqA
jnd1hjiD1a8yGzFsv9CTVszvLuLmDRDgLRFADRewHfYAmoo1zLMqMsJrsr/THalxxBnuBTDrkJfj
Bm+nWmnjXIKpPGCBQBAX2hpf7bNCJe1rJSWCxD2WJfAVraqxu9OPPZzuQU+M8GGL5kW5RVVP2pI5
FRooS2VKYxOmut0eVirIULZXETRxUMi2vwQ+0k8TxgYORqzaOapPxqF2g08WA7P+2FVmIaVXTAmH
lpD2y0LonJoahpJ4u6Nn4JFUb1VO3QH6In2qiH75QnY+TEC4ZeMnLvEy6LuQmLjn4DeBw3O8nN0x
FK4rzZ+CnTKvNLnzG3OgtUTPQVwrk+KSIMBO/lv0k7jYPdpprbTI9vAeY4G8vIIhVuIjyHB7vz3D
M02vIYwHzVroh643hmP25HW4PZCNNEuCki948suZheaNV2PdG291q1XiSiCJWydId6Cm/qup1++v
HEYBeytTjjB4CxX4r+d3b5aPECxJB3e6JUPDbFRwaNrMMMEUzrcGWHZrXgP94IXqa1+lxCbsjxRg
Ncwa81tQhta3X+BRacDdNqvlpHKY6FVjyX+MCARK8Bt6PaQkvpD5qABsbLFRuywrIjg1V83ncLCq
D9/qkmKdq53q6F1yFLeMvpyFdmqfkml0rrm5acQHRnsQOnICiWfweKHmOEgi6YLbO4PmfoHZy8yb
29aLJR5UfoiQh6ahiVxNDt000Mq/kF3esoAFiC/13+g6RVIGihbqTtDpDA0BAFZUi/9MmiVYByyB
H5U1q66jxDefxUEm9HQPlXypXeMRqbaENlHh3Ts0cfWvulmdBneknZo+NB6wW60WiTnKO2Y6WGtQ
uoN+glpIl2wpffV0iZFxj5DSe8kMJPNQ8AoW+Gma6514jDFTsaNiPHAUCPkzG/Fy2QPdhjUHew5d
lnGMPUYfskd+nwthDzei206oFSI0DWYXLjI66UmPiP/JymOgRcLMnLz6LuWjUMj2X6uFYGlv7y5k
1qOh6AyK8DsSbqIYacJmjXgCHFU4BVpW6BAcGslBfPEOvG49x9npsOHar8R9/Y7F1dvq8M+yEqYx
yhF3O/9r3n9FpaNGg9E6jYMqYMoyobnAUhmsJ6ts4o4kOaG5GbaICcCeIfUQcuih36NDF/GmAa8A
bmthAD/ZfmQFIjRDP1ueV/8eE3FrtbrtpAHsgux8XrLkFRASCjlPe3l92EKr8hxRMHFqHLnwgTQU
Jy+CQFRT7wa4N/W1SKNY07Od7/vFIRTIfn2fQQ//flPZeDx1Xafh0AmxCbeA6MkwRud4qqno9EVz
3wN/ZbV+woymURvKCrwvKcNtHUkqVjo6UtGSCzLujLNnY7CWBv0cK7VrKWRh0MFkkAwHxG/egORL
MwSYxQ+2ADvomMTaWgT1QJttRR+ecTSZVNpsAS0I1ax+QXnL9DL/y5sgNwtHo16JEybYnX6HM6eo
9NAytiay9qrAlavB5aIG7WwXDM85CqftNcSD8AiBTE3wHfLkloiPJbxJfy+o/6OYAIka8niM9apf
1UuRBvRrTV7RMQVIV2tHhciFpJH+oMF4IAwdyI1O/nFWjMZYOBDODHD1XXFTk9Wf5VYnbS9Lf6Qb
0LF+GyUINzYTC8aqlgv/rAGfH2TK59+j7yXGr8+edZUiUMkVCHHCgaSoSlfg2iAfIjXPTT0Yuhxg
enPzlBoShDPXRQ9DBwxuOfGSLy+9SbOk0QWyoriPHaMrmojiqyWpWpv3SCQqWS5gfCgAl5Gr0QC/
ORnnAXlUKAikcaO5NLXT5J6tNE9/ZnsPBQcuy7rYJrkI8g7LDOS2nDXa+lvnbGd0K971/FephWzP
sbByQFxedfRkraPZgdY+2bLeNp7xITmHG5vzn6YvbToo8Fks9Cj2mNqbijNOUrcspA0FO6KQIgTD
0wuiDET1HbhUrVjoLfBZnhdW/L0a7CpKAhqDIOnok2ct23p0aMfutuNXrUDVhPS9pSBmmQKgG5fq
lEnXNoK9Crl4V4Rj6fTtBtbqluGIyJ+V17l4l2efLJ4/LKWIHYsvpl/ctIHTO8NP9Gr+7HJzbwlO
gKHnXZVJ1vKHEt/SsRyri90NDRobQv2INNfJMgIs6+Ns08u73K+oCEyuOW/c3aWIMk/jhZ7s6C25
5ffGd7bzXLn8JaapD2yAB77Il2dTABwdXdEzOSrxx9atSNBtOqSSK8RnuKjljQQbe6rmy+bjZGM/
K4Tub03P0EEUp8SrpLCwqa5Vh7TduYMm2OzbcgVSnyw593vZLYpCTCnGgRhIL2lcQUknJxaSZes3
yyTab/USYYl0GgZkkleHD+enCOBQpbEDeWpBOrUTyicOE3F7zvWJVJXHu+iCNd/30+v3/lI+Kaqd
Ofnp5LG3gGGVzwsJTo7ZT1jCkqy0lRHqlzHwckrfVaH5seUQt1SsoWrU0m5YFCNSilrKyzXWdLAP
FN/+JkdGgngq9K9YSGAKj0eXQbuGcgPkTke1mKGmXmgjDg2A4g2x6Ezr81hm/aaqt9g4HxzbMP6c
wzpElB6o2u7Zpm85iRVodeKXzJ0fUQZUfjAL5Ps6LqNQNCjPOVNrF++Ky5aCQomUQJuLu+e6fK9N
6a4BaO/3zb8jK/2bPVrJDJN7i4KZ2xlOwiWrbA1lnE5br02RjHYBVxORwQDPIRXnQ5EJ7UaJOKVg
d8ShEq+o8sVWQocG3lkHpsKXBLFaKqVqACqrWaDUQD2Q1O0R3h12wW0QjRnPL46MtIncXQupJaRA
H7CzMs2e1n6D3V/S4qxP9g5R802t7TRcKvjCcqn68/rQeGQSVrseL4MEgEsxfpIHqDUFqJP3gFTZ
lgSceWFMfp83H3HNwVZFS1gQOn9leKY+TZgdSa4vc3l4SPcSYxpoXqmGgKhZiLKvLyMSeddmHJY2
LRfdPvTO53pVsyMFZeMXYnVmEHCmZwdaZWqnQTV8bUo1U3d6gWdyPiCW9ODA/hroXLWTNiIyQEqS
P3NCEydEqhTKrlcggME9QBqp++fgA2vK1J3RnJi2tv2+elxjryy20Q3fRd1o5htik/mhBqPKzX/j
ZDb2/O1TgwtksJkHN3yV11VerndZA6gDTFPtU3anKYkdamGJRgVMS6RXT7cIhO7nW936blKktHTZ
wRKx0lX7qc1r+fFtZIVd5euzuGuHmRobm6Zd6MgrGzqsiC3SezdjnFqcWrNG82gnMbMOZTWCp9+Q
iDDwqjPQfliqVWd2pZg0flnkCF+wXvBSmKt8qO0P3sNn+28R4QZ4hfamjoJZbarE0VBSdM3cqRGC
RVrQzJz93tYEY7bo0y4aeoS1EnYnZBEICaHpKMqcc066yFO4TiHoQ5Z0Bf2bvNthbsCQsbt42ndU
lq3RPGNrTty1EKfesK1KwuwhMpqUu5hmZPOMqmpFruqjIPwWgeI6I0k1mLMKqoIeTEzKAn/vT1dW
U5E+Ib2sc0K4nCeZzvFfl0EoU+9sDzSwmxFsFFBDWxCe5pXfPVgEssNR0qFGYDX37G92WBktkP6z
Xj0Bwa5/K11ygqXWcvhqUUV4dbZhd15/sNUAiiO86Vlk0bCQbj4j698xoeVha7sXo2aoA7UngpxF
wTj/Q1yM3ixOLr8rqMk6xZkYfp6KfKXgX8UtNmkaLV4p/t48ZT0JJmobpJnFFWOcDeqCP2N3kDv2
B9OrFZLpEPDdwK2JXcGmCAqjYKKUd+7sXsEnfPRg5en38aZrl1YSrODlfqncuII8K8k/SVs+d1aX
ADQk6pXIzS/C1t1nB1VrGEr8MP3jtjsNjz6mBKj+dR0sdGFII/qOt5nAjZry6FgetLDi9IvVY4Tt
eu84thkDtTTgu+VXdLTIjUGlcNPIFXoP+U7VVQfzKgtK9OP/UtkTrs+5rgTTORmXewwoMeAb1XIZ
RR9XICTDyXEvhH9BAo83iRG29Cjdjpg8+oWuFAODcHSneFWDKQ9cwE3zhBe6THIchxOdYz2HnbbX
UpLbiICBOchlf14bFTJy7ZV+qmPr3tfBhrt3J39FQK7Undx76wuHQJp/8VZVUXZaymJ8nGXGMk3R
WpvZD7ddvgNHKPp00HB6UqmMZmJp13RB7Ai6P8gdVXMnlGwCjs6yywt+jYMJ3Z+EhZQD0a8SWOg2
Sd+otHPmU8PKPQrJaPIWWfO0e1GW+J4nedtE1yoPAbUCbnUHpTJaA0Iis4f7uL5mn9JC6kosDc5j
AQadcOYT+Pifw2Hwp88mWo0498dBk7h2C2q3sGlJV7fKA+tKdY0lXmpJBjlRm9oxsVSlt8TeQZqF
eGL8G3OrXKu6Xr3Z3zs05aO4uONAgTUbcLfhKv+vbJx/94PeKMvxaHxeFhNv7XYEJzIOIKuPJdsW
JTM0WLYjC/WzBS8Mw5QM1qD8QiNRVYVbey8FrPIvMCvV1yvD+r+YIj/MN1GYr6+5EO4201DZBbjK
Q4FTh4KanXnSgPPVn2WRJdQXTLGugWhy5R74JXknx3LTiVdAO3krEjQcBB8HPKeaXYURYAgFauK0
OI8Mi/NSPMFb0Ys7qlWVi3J2ToS2P6s/cWlAvOI5YW1Iaj9STz6jteSm8UHmGHNbnFN1fQXfZggE
ZeIhex1wyPMtuPCd3klUWnFNERMBlgtKE2he3feB1AT4rvm/KitJA72LQLte27M06jkBhu+ZTKIU
H4KmAioB6Fo92oiKMPlr2yU4bnGtUlaeIPfXvN3M0fpJiRXtywzWSRqvDMZgM16kBoy03+3YhCZI
STMCUvPtniHBqGu8MB+n4Q4/Ef73wHtjP+xS4Qe3zL/b1ce6B80hri83Jtdp+e3BWVLGD31mC/RN
8YHqT4v6V98TzWTr2QuVjyBdfDUlHrvGhRbwA3NKTD45SZ5rDqkPlgiTNVo7zAm5CCHMPHmvCLKO
bMzY/85bfcnkjr0z2AR/5ZjKfc/Fk0QFSg1/DYqMdvwDHCvaLT/J8flY3kcyCSYWv5pTr1K2fzNx
K0YaQIYFKcWjbPxsOrYpAOTJV3mzADigQj+uHsoin75+L4YW7B55QqJpg1VkwpsdeeAwD/ZKP1MO
vL5L69fq4Oc66vhGds6KjRbOOT1GQQJ7YlAeJ2187gkkFLuno0iDNUhhSyQNHmgtBKs0wjyrblTl
d6e57XwAILSjAG8W2p/PyupREH3nti3tvALMnVivhTTsk8ZexOK6T87pEpjU2YvzlGqBHBeW820c
VZJKiRxj1LJgCrQ0+YSCpnM4rCnHbpPrE2VLUnmVF0tfgmOFd4PWX/7cgzdsu0u7Dvh8Nxq3awr5
CMcqNSObn6Ve0Ld9RNR/Zk7Mw/OPaK/5d0ovIUAvSxNCONs88tfEBDjD3F4ATl5yG+NI01guVaLd
LRjS3xXWYgQEiEVfAZx1qcEwfYeIzhmDaA/09Tl/CkJ2gOnnoJJuyH2W4i29fqdwhvpcbqIFO7hL
Si/7kjRmv3pdUCUWlSgr1sCHUF6TYEx5K9yLblXcCVHG2QKWiqlXhv3+HKF3Z4DmnxaZjXFRflWb
/qiucLP2TBbO2KvzSn0d4BryxyEERgKfUKiuxp/ylKLMm/AAHkMyQEtdVxPc0Elj+a+WhqaYiMTj
sqq34lMDAUgrfRsAYKi5sPqzbJAYkoI3v9sr3b90vj+FkGMlGA75V403ZTko+7c3/E/yquZbe12H
krwJRId/ZXCvuEqH7DJWCbBTpL9WQCwn2g3v7zz1dReWmVBOlaP10yw+w71uVeRmaLXHAUz89z39
VEBXNGK0MoS6oDKVPKvE3Q1rf8qwR6JYJUbsMFoCMR+/o3uyCwdII2iljgXGmc+52188hnOsuMYl
gYQahTJHAwAtnAnBmksKsPu/2OzIINFkU1IZQx7P8Mk7Jrz6QpZJwWtANQUZLCzziFtK3cW0qJ2R
18QKFUxKPmUvOa+PUT1YmyhiWHSqNR5ukkIqXUdj9TsdYZPa/sFYsy/xGVrN1WGJlH3C0GKMGG0R
YQjeUJ+S1VQEhOYeCoJKvjQDewzCKwEP/coL7tmjDwWdgjxN+NTEaOUv/NVSzq9ZRFbK3xDdkNGM
ddJlItd3JiiJUBAhGnvxtOOQePvh/ixoxFoSDcMsa2DfFYqCVmLunAts2W2v8ZWyD1QRiXAY603O
lCSXkXIce3lr2GUjlsIJOVaUvVG9ctZmW2xzIOQdYQwy71NZoDGi7fySo56723a5iN9M6IQtkr1+
3Fyt5JRa3VpVr86FqfixN4/ZK5rMa5+zqQ+kI8zLQ7uwTPiUZKb7M7C/fQ/PgOwU9dRVU19qi09B
jvEU2RolW02N4pcUEB4UxIOjmI30RJSJaZdOLGWgEjCsT19Y/wMiWXwB/UTYQvC0Y/lqBH+mwDWl
soWNO6bPr/fzGjUHQat/NvGH8rwKuDF/TEdQS7hBaKNx6m48EI32vZGEbcSfsqs8gaxUMyb62Ye4
ntJSVE6W/M1SLjBVeW0IWt+2FJGCmpkaFlBinFtgrP5sb++V9V6TXs5H8VLgK8AIcr25bdoiLHwE
PEy8XGxKQ4zHdM+1l6emmtv0mRUbQihKHJTqK3a1+HcBkkeU5nuLcKDwE7Oej+Z1xq2oZEe8nXL6
2BEOeYVYYgo1a2ry7JLiEPDfZ7soW+76ZtceAgtGNpd/aaT5Tx/rJZ7J7lYJfVKLoNAFA3XujlN9
+veN5h09QCylj7xwZVbpwjiECJ5gqFjDxD4ZBbAW/hHeLBvuiNL9JVoMRlsrIMTz8SFnjw5SPGJF
tac0mWVQYJc2epSMsia9Mewfj6Snp2CHmIwRyELBN7J3O+zIgCUNzsFrKzWc1n7TfnJfo/jYWzT1
uym6zHaJvHuW4YsF0a9BC0+lJlZo3fuSp4FQ3EiTF8ZIOv+nxtINMr56wpmbXR/JXNqwe/zosbkH
3wQIH/NcO1lfLls1rU2QiQylULGsf4cvSiNL07RVEmR/mAKLJibPtCNpKtm/9fnrFmd3YnskX5yR
d83HEzcdUn4p0Vu8M77Sby8gBULNnFdWLmIiGjlJOZjfQdOnJZBrCx8CmBrf914qKUqyfawe6dTh
kU4qfsKOxJH83zPBMZ6rba9pTRR6Eo7XF1O9YIcYn5jiGFIdTSEWfx7+GG5v6m1wLfHofMjIMRB5
AAxdcZbTBC08P2BR/7CYtorO1TUkW+CjWsTGcHhJQaZRG2Ey4eZf/Vh9/v6MyyH9ponY/rTkRHdj
6Min9Rq2jRe01pd6tcg8hK80ErDRfHVABSPR6c/ZpFl0YuQfE+jyJ+OC4PtvBRYu95E76tDXBoar
ydmr8kJyWWjPUnig5ql9xE5581Lg56xg8pdbbRdR91bk9YBVB0drUL7jn1JSsbxBh7xDyYtekxPE
V4geH/kiAIu6hipJc7KqxnlzSaQxOr3qYB8vjqFK5Vz9ph0jjunpkzglsB4EKhn8FNVW6OtsJiy7
IZI8FBxOuizAzAvBRkO7ZqyC+DuVBZ2t5zQdzlAuybs9eJIJyQSlK2/tjBh9ZCGras+VHKmVeSpL
ZoTlUpSdFpiE+PsDzb9kc5qOFWy8R6AS6wAffgP9WAUCCCNkVqrZi9SJWjLDIYpXVHP43WiHzDdB
JwIe38hScCS5icNNb1zLF63z3ltozs5kRgfGD0AxMNp/eiuCqEpe9+tgLeI1ZqZ4C1tw+fGGKmLi
uSVyF1y87zEPDAMTLNU+G1tNlvHZihSGb/3hP0J1y+nn1a6UVPcp+HsNIhjA96UfL3uPimQ8Bfyk
UeG9qmFItqF3/0HWrzlfPJLZj81S97xOKhDbPrYibdROrhc23JHz4+YyxWcpI/BRII85JDxnIMEa
WEPwbZqf4uL5idBTZraC9K15LkfCRUfYC87eb18qYpoMktopgXxdF1m+el21D/6XGRmqjEAjNiYh
LQbBz8O0btm04NW2glde47eovxO4KUqAefSKycPsDm3kubWIL3yBMRfULgSrHlqYGw3d/rNIGg6u
wsa+pgZS7mlENgp/9p12+ryuBwLrrLHk4V2zEdMpp1uEzzFDBwfAVCCQ/AwK83f9D007RNC7pRse
r4y968zukvLhGCqTyCQLUwBBj5gTlFRG24DGOUnytmdFKPBkRtW+WZHhEKRj992eGT7/e36GmyLc
r4erEdTBqhaa9XBAsz3Mz2S1QU4N4JIYvvBHarl0uz1aQ2mu5X1q9E2Cf8ZmrxmsznmL3cEdDyk9
gtR3AzP3ArLrRuQzTte2UN2LWqDv/7o6ZMXQXe3SsduWNunSNVtZfNPeCTztPVwZvuwKAoqUEfux
88KnYdoTJIWGP7M5PW9hfQN7qlWthgHzViZeo6FHPuboR35l8qwt+KN1TRaadNotAHO9LSM9Ntlq
tRbU3na9fG5YJX9ufWyBQiuvKl5BOM4/81BHb802QZMczbOiuBJS6nDSZqq0kX31+EidtAk+Rv0/
O3Oa+dbYMN8sm6nu6iE2dhTZiF24cKCBj38ityzshy756kUxPtg6zXwvxw4cBFX9Acc8v2lgvM4X
fteQwrXy/1wzOfNX294VXiy0YP/RnTOBmn0T0gmxxpyTGET0ZL+Cp3034FsevcGRRSPmz7UbCZvr
K4Ymgini5RKJJnfajaZmR4k0ZBK4v+DxqY7cxpIOKt6cN8+Wj/9Z16428WmFvhKDa4Le6Nl01bVd
/fEufd8e4jlbxvxOQ3qMrhAUHymzaUHCYpbn6J+A9gtthIrDMhA5LBKptky5l9qD/ACQ4fKzzfRo
UuIiEerN+nylHi5zvyy84K/X5QB5dYDpoIShtb7Yvpv8lRSqfTFezvpd4K9myA6DumwCzmN49BOe
y5/8neC+ps1549pm3xCkDD5csC5PK2vjtp87Nq1cw9ORJyfo+yvqeW6zR7DF32m3Ht9OrdlX/FNI
j4+XCilAP/W4nuUu2GXvp8BYSgn9F0AR5SG6+PtVKxrOqzmKu1AyJMwfJJNLcfvHvX63MnUexh6O
9RW55VHX82fyrBNxdB/UwsMrT6M/1UIQjgd8U36GzI6iZUYo3d7i4KQK9p8eQdthgjO6V1mJdm81
jt/LfKQtcthnM9FlPi37mnMnY5dUV3VH8GY6+VBeuzx3DF0Pg/8RdLXvA5Po8U91fCecOsRqZta6
PFkAS9U0aF6pQ4GM6QcQRjkCKTL1UuXqLPRItVbhxLHM8vqib0vog+RppaBNcQH+bG+37fqzeMIU
9c7aoD1kUFX3xYD5JBNn9oYXDshw+VMVtkT694l57VfOivs22o64lwHZpt8/w+IUIx8Gka4NarnK
XP/8oPCgK5ylbHIuMem05G4VoCp/N1foteFE+H1H3WmpT3BSqhGPGoSIlEVhW4lRoWDEIo9N5cth
FgO9ddBXM8/hsNHfQwVpCp/fINmSgSVTjGaBQtpVislEX5uWXjnAvCFU8maSmr7I11aHNKfXEOS1
UhXoTx3gObUER0e51R+WLQvL3Rqkt9IuFNJiqbGAWx9UkdHEmze1l4VXm8ytXVZIAMUh3hrAVSLr
fqFC4x7wVcyUuG2G8Q58Sh1dCl9envkbPcvRiTOsRMzui828eMO0DGWuVgsFHSK5wjBv3we6mBf3
zdwiyu8MJtzHr2NcQ0vpDb2kevTs/MRyURO+cLaEixxFDijz4yJMfHGsEGlLiZ58pXhgkUZk6kpw
qBr/0vksdcYf6BKrnqFEskSblRqpBaqaPlVzCcldT6Tdv/NllWoy2ZOQNddVWmMxl38ejxLnyJVJ
blAnijfy+PtJ5BPHLlsgHnUhvqUimI8rBDDSFpc2Bzh3oarMeBUCG/hiLkl0lIXf1cqbx6JekOPR
XoGi0/4mmOJnFmFjRGtwSkM2EeJ/LZXxGPR1rA4jSbl1NZaXHgRENh/BPSZ/qYOYaP3Uc3hJqMgN
Hi0Hmu7i161dOTjhIHbQbxTF/Jw4dNRLgAEL/9zm3c4L7AD/h36mgapMLiMwE0qpvK+GAIGbIcFC
bhdCL75tFdmYV99UEQs7qkSFiqJam1/sTcFJAuabmVvmiIbnr9wlgH09Qx0U0T3ieQoE+tgFsabC
+2SetcJAKqeTDB/tdb+aeBP3FvLT3MmWDoJynKxhRv/VgTvd2ki311G8MtfN2Ro8VBg9a3nb1zHI
aBoMbeGNB1GBDs18zQ00ZHaULxaLA95/SRHZ1oJrrPuOkyOv9TdUuLre3DcKVHgqrtTn9LP+iLll
SGTJjNY1nmn2ZThV/dG6GhKve9xqhcOCWIKVMwuLT4L9HishvXL0GsjqSyy4FxZPXqJkHSNdGTs5
HvKTyIZYEjuyxSUuKERB72JzdNd0RRQHz/L5x7Elt/zZmPyIBr3YGLZZk6AOkNNuQXQca8m9jS8J
YyNn8tbpC39v+dGLd97Noo7sYrtYaZ/WZ/15BLxwCdrvmATYNywBqQY+uZYGCT45qC4bTbH229O7
epAgcO8lsQ2iU4/fmisi6FZuMbpnfDqGR5Y26U+a9i4qF2BMRy2bPNx4plPzBRN0SSzqOLqDa4iK
exMMnyCaOVuE8ap951dKYTOQOJ2aynxv9jI6OHCfyGbOHIvPwZd1ZEk+MloicTDeKC01iAwtSdJs
TektBukgWTG0lEoHui9Bm1flmm7XkVeGrdE+urkFva7HmGeUIY9ci6crKhzPumM8jLPHL0+zySSS
8Ev3OcEB4QcyIOcnGOMRv7PflY7sNIa+QP2+I7DcoHXhi1m7HMp9NPKTrtJ/B1G5va6QdpWr+GOH
noqa8Tp9hO1qTom1dG1qTs8hwX/8gAxirUmj8/SsmA3RPEY7KdtiAVrxIq+cp6Bx7TkXJESxhOiH
edUuwkmBhWLw4BvTLW31avxBNonh0uiuFSN4FJrdvZ1+AJ/zufGmiS+isCPTPi0cMw086VXQsaN6
/95Ot33EBeeIp8bg7Z/jd0D4ybS7ulQZuV7K1ApR0bP/cmN9kzsFygSRk5sMHBTci+tFGi8sABmm
JtLLzbvCBwK96fiWPon35MgxDphGkIOULV/egRlqRnYqj0ijgE7JUoqJYbNpEqZMTXFz/o0jiBvK
ZXfVWbmeyZEEFc/OFddekIlux6DGGG2qx1HXiC7EJMNuT1WV4u1+weuvpfyq9XEchiCRpCVXfort
HSlKM1B5kzWiAsnFdAULLpNOT5GycuuDyf78Wg0uwGRgv60RfjGjJSL1DxNuelu+xIWRAJyu7405
poVvma3OF9e5ZVt+w5abUjeNmu4IfCDCYIrlmMfHOTBlgoc4LsMobtBRmOr8OgvMzyc5degS/bSx
v/QEKqYcpn6lTKqJezNOoAfBSyhw0xiHD01JnrJXSmOvIIkxeEhZZ0Jsf0TLfSa90tT+Vt0ZknRm
1icUStUBgtLSBca1NSr26mIX35f2tipVcTNCq3OLvWGwiNYO8XE72Kg4OjytAyqUxJYMuCn80mNy
9RxAEiwVwIdKC63Tv4uGJ9FwdV9vYaP/GJFpdve9hFRpIdrrRWg8svYaKXwPBgK/XLg2Q3oWSnY7
s2pPsAlNatKxwqC752foXUcP/oD6EnjWkdDK2GQaN5dAUYa+Yh/5c2cMc+pnLqc9ELjnt2EBvknD
bWhubK4KoH4UtnJhyy/F/DgROt60d1sgKw2QUaOu2MsEkh1UybqtFeTwGXtKYDfLC8Enan8V4llo
nRefQuA3JpMiNCtRluVbUu71280fyR8RBaR07f0MyTS3lgOzD4gcRUhd/50fsPJAM0bO5Ijd8/PC
Ae5CKv0CEH+N2bOThpzj6IrTFluj6+h3X3HLgAW+hcEbo9BbdqrGXgsQePahkld9StO7ymMxRNlV
cO9TTSD5UbZ0FFINtYLTlliIGjcwDZH/Xr11ow0QMYTmDmlS9vSzC1T1VQkFuamZC2pNsZDcvUgL
8bxriQVEbTTTvWHH10Z467PvIXL17xyQsv0ewNzlwO3YBpo7SAlFu00xidDEAfJ4p527JSmkqu3H
+H+Arpz4flH+xi0cX2CI+Itb/BzfVWUour1IBc6SxIjZ7pSbtuHvNs4+pONLsNH4PjEFqdY6W2bL
SXg6tiUNXB7v4/jRJHzjeheBGddZrdnkPAGWYeQe/FD3lQt4BTZqV1DqRZ7ssPUYiE6epFPRiv4b
GhuA9267Dfj9SQBDYNP2MnuA0D6xow3c6Z5ZxedIhWo6+4teGrMSjAQ8EmPznCfl6H0vNbzwDVfO
KVrtLeavwXQPqsjl17/nzCs8XMDgG4P5J/5P3WBJhc9z4kfggMUIx39/vQWKku1LgscEZh3Hb4pz
bDcpFgL8Fuh+nMfgQ0DYGqLScXwnJGMhrYqEYHnIv9tVQs6fyJ3ZIZ4DMhbxl2ILZbY31ND9iI33
KBzipgiC7YzmP2UwUuvApeez9GLh7PYa7v8otiUn42c6Tw7qpB2zago4zIH+N3lB6ciLakpys2TZ
CcbxVIzynhug23ycaSiAUnJaLbn+4bs9OCrj+TUHOkBJboxb0WTnWykrVgLHJssbcv3tvtcM+LAJ
NxPCeDJUETLXkTqVc5k/3P/04mSeb38+06rrLUUcVpxtcNWFqHLQUYuH752ksIoF//VwKCC1pfSm
6r/re5sKwdt6hbOCoziR0wEEXPPC7uKRWF8krvQ5i2ipseACZN49afgF2OhUW944k3xP3Awu0g8R
NJtARyEzY4cEjJhNYZKoqfM/fCnbOGbPirKLFa3uEqcbYHGZbSF0GUaDaeYD0GhJOZ7Z5dMVGQHn
I3bihI1RNPhR1CrEb/YgqSeiKYFY7xTBSMzai9ROyQbIdRj8rjC4YagxYkQWN3A8kYslPMEPOe6x
/EYkXx+0g9p4GOK7rNIIsBI7e7/tp2fSPhJONT45wbggJya0xzPxsUwIeYpd5d40Yr2CMn9GC40K
aR53bfA7A40oNOAnh3xqWd+vnOi1SkbYAOUH/AeN3WwAgGPBlxGkadeJIbHi9nllxJx3GG/JeLa6
04fhxyChI2ucjKumKBqk6djYyvHVWNjpj+HM8NxE0muInKa6SVSBNXleEtlfrvcU03xxlFvexmoK
2JBP32XbjL2qUB1ZiIUr+DhQY5SToSv1tzyWBSf5DGL4U5iHVBWD2mT6OKrZjIbBy0jZRs4coFNJ
vu2j3hKTuG6juImic5fFJGDUeKkcaF07avJRGeU9ZCIVYaCs6792raI18wDzkhNUaM6Puo1RjRfy
WCvE904tim820UgLnGTVilaffg4Uv8uglveSC2e5zwSCEPJBGJljT5AXPFdvsFg7/o6cbLOzOomn
VuDastxsFw9DrRsJvkH57C7jFJoRegFGfCfQOGTDzcTft/d6sllgQQFeosjImmFbvyT90F3VUmxx
kfuH+hGGvoah0fjpf3ePSpOATEfbOuVK0UPQ1JeeOAZipo+vnjnOSR1lvNketNtLI+BR44ifoEch
p5q1Cosl62qKqrPLYy0E14hOEEjcFfYqwQcODnmyFkfiCP104Uy2M8mHU6hJG8DE0xOwHPGujIxx
qUfviY+m2HTd9oIr/dO96ToMDwYAVGwJF1DhV0vrM6kK1El/s20rFJLiuumLFswnWT38SRpWsFYb
ZeAT5O4f/TZFiGQaQZTxA3TtTHRQYCi415oWvBJG0OVyfN3yuNanfmnGx+N3rn5RNCsUNSBXTG8r
i08nr0OJ/tM52/rK+b3DBcZe2gvYXuEV4Z2n9eN49ujmmRk6WDOfrrW0QYBOZBFWvcieOZO9Qy/a
FN6hZCl8m3mFydalV4PX36HAEl2/kyxtfAkkPp7Ne2hWig5vF4tGEmrbk49b/eWqFCkOoa+D7/bZ
8Y743YTjHxCPyxV+xNE0B75c5dt3xo1S7kco0zttYeOcYZMF++AtJQhc8WrfOViIjT6sVyyhd7pQ
GY5dE3jzuJDQors4IHEqjQz6dQunGEvVTGCcAtIqaFJ35rct5Be+4NbBHYfKWsmiWqALmAGqNMDx
U4b06WQIBbyS/Vp0p//k2SgPfq51yPpapITEreTp61VvEB2md+zwdD9BVluconvdTiJ0oTHJS0wn
0qpf33gmQ5rKSca3AxH3q3X6s93XeTkCIU0nWkzXjaElIrTIhSOs9W5nlvUBtyIS34j7TgJEIgOF
IRNPI1GPsWfNhrf1mwdmlbNih9RTOpnfxbZ2V2AGpRDgXAg90VYD2E5BP0d10A3SB7VNt7cJzbyq
HjHVPVoWXoL4TMQjUGuwiSI1t48Qi6Sa5ch6C0LtRPHbIi/AidoMEfxWoYCpbv+AvcC5fNv38HEh
SOgKPzJOCwprWuWpdCwD7E7J0AtcEx1dyRlP4sEIDhxvhW7X30ZsupdYzlw0nquVoz4jyoly8BN8
eXrL9uyP7Eq/783Dqs2vRhnxPaPD4sIXi/CiUPpey5c8mvZ7QIuzq+LEIYTj0CHcw/wV0aXcJgp4
tN2MJqx2KR9MTQ8aUGuTnT9DFTRGsGsXKOnhi8Wx/BXVu6+uoWtZcztZ8pH6l4m1KMNomiOdIQQs
lkEbyzpRYeT2hcIn/7K7OBLa8J5QcOqIwLGDjIZqrn0Ljhdc3EO10lAbaeoJbUKOp420aPC7U20n
b4Itl8XwT1ZIXF3BphVrCbaVtpja306TOEk/J5pLN1MCecdQ/bQ6OkTMMyheJvLDQ3BOlb1hkqo3
Fml8GgftjYSoUYSmIZmn+vy9UrB9owXwdCVVH4Emic+zoVuJQmDLOpRLscEEJQi8j4vD3IIK7mfQ
0XcHhGZylMW2jCxqp9Uv++ir9zqnuMqE48T8CoKO31W5e12a2KIOj50W6ukCU0DBMALEdLu0vygO
zfjoKm0j8AWMJ5eGYENHaoBNM/phVsmMJZaUvKoXee1KK5r0RgsJgN1UgXre+s8co4EWX4kJyRIJ
8DJPywS+d9SHNfc+gmAcgJ6YCz1KyGh6H6a5v2+wIwNLq7uENskOvKubGUs8RuEM1ul45F5eI10b
Wuf9doaas3ykLUaix2pe1m28Z+YokexwszGxDIgNXkbnTuj10ynF8dgBMHQnOUkCn2YXxfKnMp7P
aUXcCDE2M9dBcTXwDQQrPy1Q/de0C0Z53nys58DTTPkH5JvPNJN2U9yAvYJAPEksnZBx+OqOtlXI
cav9qnWEv617DcyZWXb94OyozptrdTZ4k3I1v0f1TwB+3D2jR9byy1RsKNvP3uKFTBFPXzKle/lw
T+DqqAgYBwD/zvRAWOrxE4kFah4eKHUrH9NxYsJmM//flftQvrbiiRi7SApdqZj/cIheM5ANHvVd
pXGIO5uDHXo6oRNDATrK4ii5+uIOD4Ft5pnfyOXaJCt7t0BgFUuCJ3RvykiBOn7MTZApbwg6lob3
S26saeE9uAc2vI7vov+UzP1jOkOQieO4yIBzvUZJKVetKILMk676gC+SaVGRL240Fbi/mpNFcPZW
J9DgDSQE4HTHLxcUTwnmDpxiU35PwRGBCX7PsOkHHTJ4086OHkh/tEz9+C6aXRa855G0EV1RSGXc
5GJARZO0Z0qUTAgtPZm6/izg4RPoQKFvdprhfUB0R72W3gbtwk4u0YgWr75rSv/QXUN85cd8avXu
L/kHwt5SUquyzWu9u8the+wWaSn5Eh2csBIlcWZeu2Rv7uF5s0CefsOzWgKfZBCln75V/ilZkU4X
UXUBUuPB1fsoKwly4JxIILgY9NbK7feGBP75/jsKugY/LkY+py3fGQqYauReijCz8k5H7N74VhEn
1O/OAraWjNBd0+171HyPIBNfo/B62B9Q5RjgKwxxRKoXdpS969NFZt63O9CjWbWCeUrpW2GB4Kys
60s6ltt44+2EI1DYVxbcWsZo+Cd757Ns0rxNwlpTo7T03/gvjcWAY+71aMZh59Pzp2eZGNGqDwZO
+HLT38Yw+rXUT+cJcPXQPc/5ABgWDR8Kgfagn3tHfpwX5x+ZvjFma0iCDQ5ouoAv+IDQhITl3tK7
NyGoTqCqlw5rv5mxJmEfrzbWsXpFqh7f9tOEaK2B+YCuFAvr5pdcEkhSNvgHuODuzsPRZU6OIpRD
ThkHLFY+jJiNS2REtwLlg79fFf4N+FJwcHTfW9RZEtg2nxkDCtDuld3KeX+zoaSinu0m+boaBwO/
P04ZT+L346dT7LbR18vCZ7DA+fo+E7r5UrX0WGWixQW/7mazCBPQIyiE/xdirxgIVxMvZSCFzQM7
KSdUKbvgnrTE6DCeOFilonZJkid+S2w6BI8SpcbFxysJdXrC4UDe86BVgvKSuubWFU3G/rGhx16/
AiKorrCkQvumwzgEZKXjodAuxOVf312+dNBi1RKwpDf6DNHj0zKIE5hUVZP23KDUBO+4OlyNQ2Tf
9D0u4vvcTsc/WS0dY8786xGFBFiZC5vMp7GarUOe+DehywROm6wQ8wMEJqAG+wjBAH98rn1MC+BG
29MeAzEyzV6spQLqx5QMobHwhzmMuIAK0/uRmxQ/RuRSgK8YNOLdqnIVnadw4goNggC69SqatpyH
ojCbmXTX6NHqlvVEZrgHmL14cX0gqI9xBCx0PRGnOKvHsqYIy5wK1QXbKftFh6PBimkXdF1OEglQ
EZ+jdaYEomxSnOfFRhijBgXaq+WlSXy1L/5N/NPerwp5sTipXsXGjH5aKjm//oNKsVKACWNtKRWo
1bFGmgtk9oc4n446ctf1F7m1q9GeQlz7YYo7IVLOtJpkgcuPsgKObDOXUEHwFUGuiXKK5U/KqTRQ
dzFZvQts15mGDbLZQpih1FYdbuBhEFMBgntQg1ZeZFiVcgb0AyDa2xgHqhZHEJVhmkUPlwKtIWA+
/Q/Tj952au7AwWIrR7s9/zccRMjqe5MQM4YNhoCdj+CgcSJ2dB/YHDYDRwBprmDpJkqR4diN38vQ
mJ7vJQN06C1EqEWGqtAr+HDoouwy1FGCJ4FrTFTQmYfi8GINGgaHgNFMfohH/V7qDK1kAGxWyt7B
UieLdVRrQLe5qMi5t/yniWXrGt/u7urMcs4+ElII00h5VrN9mvxeUZkP5QY7QEbU2Me2pBVs0fAJ
FN3lS3kgcOalJJ2XaDVMShF1n0POc+nOkQMLyVbJY9AaxR0eS8eQB3pYrcXPaxHMMPuAFhH1Tvqs
LNs5AUHrzvXQiguQ4LA3o/LlMS7AsbUkeDWX7fyMlx22VMQlpi+m2z6p5XE+w9P2wv4zqFMngCuY
K4wOsMTk+ONygzGvH63ZkP+Pgf3Kobweb3JzOuHCRwcAzQqznPOLZvFvT1Vw+rwVDUn6bM4Sh1jg
M5UwtktFdtipvB+BOKb8AuEe1Qa9RL/Sng77qLG2orBoG+ufJZQdk81arAKsdJ1FMRSUCGyKQlvZ
0lg3kq0CODo9qEKVofZN7GXhZm3gbh+A0zd26aYB/6FfL813ilX6DpZggMcnq0a3ehNO3tUnibkI
3Wa7T78UVcMQ3VAJnc/RunGCWlLzjyLUBxN+ArV+6i74Ic+LVdhhPuCnv2IXe5fGPBM5beaLJNFG
Arz8W4o4XGubHFdZ8q6TeNOTxLXpD6uKxRWqNRP0YlrP97zl4z/R8bEwyBo5rbd0GWBnB6h52l8x
GgBZpim/WrjGlNd7d2uHOCsAr5nqol23yMZU9n8FtMpsO4CvINpALLOYsb8zgLpPnsNe/eWJraLo
00w/Nh8VCCaVJxPXhN43omY3LtApRrG7d3G/vqCCnBuEzZDADQLPKM3UPsSEwJDhD8qL+1SEdDfF
NJQWGQOOcdjJgmYIMtUTl8/IJ4c/zKea3fsBBb80IWmEvryR/1zjJwJ+IB5t/zVrqMpdcthyRWTc
DWY7ykSTYR2UphZosYa0a00Hyxpk5N/+4T7fl0GnRE4kU9ZKq+i6j/4zk3qgHID0NIiQWDH3Pj+4
yGcuy+7W0vi/L+bQ3/qMQqoaIXTef6CvU7ALTFlVPj+xq9fTi+3esIPxyeEzXnNe2gfgfnsoME6i
43mxFwFPMfV9BtRKo+u8cjnAM5E/b8rXDJ4nQpofyVAS0WaYU13afRs75JF+s89TYLJd2jVMLPNo
OmNXFBNfUCoU14C1SI/sdZ+Wy+npYlYLyfO2WW9BTUqOKl5aIcDkIWMQXE6ezn5LrM413UoiqeLY
4/7bI6YAqYP5MEsaWyn5ZT1q51O1JVJXXFwFh4+GvZoknGVutl/NZ2F/8XvRWq6x6abCue6QC+Xi
JFSuzTSqCINnwQKRZNfPqzQ2cetPh2pEiODdn9z24AbJElxotHN0JtRb355Y+th1i4S39JmazDwd
61b1HCB7at16rQF2kTBIzM/LHsfm6Zunz0KzBiQel2z7ht40oRwApEIT767p2jRnZ5WG7RSCp6PR
NM6NwNCTxOW4rgRGZml5hBqVwSEFdJOYd+AFxiut1wooCEKagqBrPCf68Tbg6uUI59whIXLJilQR
B91T13TlFA8hIEpzx6KHrjuNuOo65SmUdMfWQdkuK5eQ1K3be9qpy2ZUaS/v5Wi/7gfDZq1Nd9Bl
iJ+jr4yuvBcTkAEpSFZH+PzjDX5XFOioy7IaZ0S7QXV4sV7VRrxnXzPAbv8vQkFUrfUIvk7mPXR7
4ULfo+Wcg+3yvoyTjM6HNLYLVwtw2xjmjDGTuJ+DNqpp0umQI/k69XfTDSkEYnjsQR8ehfSvKkCw
lV/JJ3aTP0ZbLDxfFdrXpFML8fNiVFn2yjeamWAq2gIdaXeou9xZ16VnYuDCb+46+nJX5mAwiuPk
mmgIZ1r/AkknW+wLav/4pA6ajsdpoOSKevuBkle0SNSOp+U0gn+mbmaedAgNIRMpwXHcHL3/SPnm
zm7YhguMKGfU72PNJV98oyv6rWH126jZ6W1kCoXQX6S0UKzRJmTXqkXsj5cs84g4welaeAQXztBW
KHtAiTcGLNW0IOdgAuMLzyUVQCwJtaLC58OQGnWENiNL37dOvMQ5VHpfIdaG4jsTdNlMdmmaLM9L
4hh8X3XcAWsJJn6jMPaovcHR441StlqgFHL3flJRlxNtUAjBzF/yE4tStdh/1rkUNe7tt/XfP437
PrvfIlGj+Y1WG7buZq2ZU9P4/Q+epjBz4eqYnx7c47l0SFwtB4Ro4tCRrYl/WxRM2m51RUh4qHI5
gP1XsKwxeeoHR4YKTDXKM35mU+F92OaceAOdk7aNfOxyudO3X9y9CQqSFBD9gHImXRGV2g+JTj2K
KyK5fzNqNAur3lxXSTq6Y1x3xvdbKiY4XP6Q+unmBfrFMTYBymj2kxBLCrhLlX6SI/er5wJExC2q
MqKTkJZ14qi0eYnVLgjy3ll2eMWjS/hVqQiFg2AsXh3QKx2bxnTQ7e4RWkEgbKBKSNHrxBa3U5MH
/Fhg7e0t0g8sZfeVDR8u3DnHB4kS9J4+V44RNhwfGRPx4xfbowkZZK61vTz4xQSluPT/nMFXeypm
rPoKVhh2kS+XphsXLVCLKvZTg6m3uUFytzgZDxCRF82kAUSjQUqSwsNrPTMuf896reuUBuADcStE
J2G57OMjK1Yp+D6JWjXK/w3aB6FDZITDs2nUGn64ahDtuDg4IYJZeRHC9mdwPVPdVFb4GLBOOfMx
tEVg2bYulQDWgABbJCknlmLBSYvJgln5Bz/YRYCS7Zq+mxswJj0oV8zUv8/G263lxq+ju+sqfbAP
vEV5gixS9cL95dsEN6ijTovs+ANpLMjvsiDzJeYIqtG6zcegx/iBN+zmaiziDlqy8F1D4kFGWemm
ewMRFiacezxdDNys4wCZZ6KNqJTUf05+MLN9g1PISiWh5df5qQz6NnKXBx6FoGaqzDKWqAcse3a4
qtrMrOEFzT/t6syLuM0dlj1yLuB1hyNGuDdAhoPjp2QC7i2rPQW+W1JibfNrapXdsIQNpE5rqX0b
UwoybEd+8sINqkgcQNJaQ8TWrD9n2uXAGScikQ2D3Jg/ttwN+1N5c5WQeZqGC/Ub6gNT2IzLbCfi
rsbcsww2JXd+U8RqKI99doebaKOWxAzygvtp7OGsuQ71WBwLWQW9fz4xH+FqWSZMyKDPz5rq+/1m
lrWdbtaSUUzCA15bzEP2cYxBheR5uWFNjn456Xq6nHrDI+brbPqY1xKlxsaGxKOpvpeVFRW4EmZZ
kT9rcantNC0hMRox7gQ9n/MPmCgrRCm/z5Yp1dxMG0XkxPlWENxtvH3EOqXooHF6VHjW9wfKXydt
ZrOZ8v7Wg3NHu5LG4LPOFQ3cnnQPWXWWZqXoHW59sMLLVz7znakFS6J6X+lwMD18FfiYzhH84cOY
yYEPJshWEfc0MVqwdPW4mwDX/QzCuLw0olg7JHxp/XbN6Os3uvNnArzJq7avqyNTGOuPyavSmizh
EZw1FsxA5/awV2En0jjaGpJdBVrN7CVWef5gLGRyDPJNPQmk9vS0JqYyL8kVUxHtGu/GNHoXQaBb
DbC6/Jx7XiB7wD8MuUGUGHsBFptFw+h0VdYmcxpSxr4/Cn+YhWTZ0weXQYV5ntbaEztUjOQpAAgd
9SQ8J/FJhE340D8EtA/Vmt20vZsr33Cn0kApC8DF2GQswgpLk8B0/tSu1jnask+k64HiV2lDBGjo
v9kIQl91Z7dklCHyU+fz2vmCIMUoxGCG8EpDfOPUgNbt+USzjv/zeIXVHZtFamCJ/y+IQdVTUAB6
RFxqhTL87U6tpIYiyUNVwqyRw3dzuPg0/8BCgMqUE9i1cDlLaj6W5U4jikbiTgPF+MOy7e2r0TIV
Bu/sYNkpWb+ErDbm9/HoLd8UvTikPcOysyVM9QRw32A+daRF/emEHO2WfW0Nl0eRSCrfYq/SOLw2
0S4VlimSCrtUfFjopDu/ZPcX6rAEry59cJa8Y1b2/Ob7Yp4btjnNN0+euyLL2M67BsbbRs3M1TjU
fuFtGTrHM3K7ieuyOMLKAn/VFoG32BOZ+FcqomZOB9/FUP5WWqm7oOxHCgfhohCTFrSqqbJXoMPw
ihnHkDqaB7khIQ2/Wpve2ww/hj+IQVhffw+OH3eZlIIK6SGHduGvhhR85ConezCvyw81I/yTRY39
b8Ak5ddH/CSs9Wh+rIkJ7WNGkoqEyPPRrtKB94T1DvSC+/c98cGP3d5q5UhIkSJgXdDqEO6St+Sh
QIN7Q6QEJv6v3puDjMM9psEulWl+afszJyeYQochabGVOd99CMW+5d0gM9xtb0WCxuaGv86x51mh
eTc6uzJ56VqHtq0FQ1TZqKMjnAnAf+iMw7mNQj54/lvwsqku7cvMc4NEjr5NIEOAkExLX+YA8IyQ
H3QGOa//YyJd2AfN1sceeYiVM9NByqoQqPDMnQFT5O5qk9XWHsvq0GK9r9NI6ZO1gPJn2+bBJz4q
AhrGniOm3lfjR0SxcfODfvqwk55at5wCRhLMSbCvmvTFpDs08ynYNisp62G4UmP/ed2QnEO3yAK4
nGBY6s3iChyJCz1q+FFCGICNEN+U9046okFL2Pc8DEp/U4blK0isiC8q9k6yChLUg5SJqats5AiP
THP71LV2KbDbKH8g70HNLLM/rVl8gncaa9rcRNvck6JtHVDXardt5kHkEdGfP7pJSc6A4v1v3BZq
sJIOk9FQ+BZoLngzoe+0VUtBBXoQcAt5My+0uw0wAd6UluKOZ4VlkDx4bB8UoLyICOtHqd5xGD1h
JD6fO7C1PlO+gUYVoLxEW3lInDybYhelE63CM1pDCrSFjcWHZYjCccbZjp3JeZd0mzpFJhRT3cV9
55DjvIEN/+4JRuZUSP9/zBdJbcKCrx4WxeIn08tDhv5Zv7HeFzfcR4ePb4/0xu8aRVpPaVItbaNl
BoUuSAKcZIOQq4TwTZK0ySQZnuA2eTv8a2M/NDJO7jgUWLDL6rNmQ7/lTzDY23YwvUHE2eQuDh7H
6T+EhE544stTnBgZROIG5agwg8oFYwznjm1Lge0uuLfcqSf5aNqlGESk9Lwj/Dh/Wg6FAkmwQmrr
qkvW5kvRUJPkuGLxGT8x+RCs5NRtNlmkgsOYzwDbZz/gFgTjLitD4GNHcrLoGX0shlzTcyO/gaAr
PXy7IN3K10expRujqPDx9GZDu34GOgHgrz9QD6fggpedcK7oZcGbaGpIcY41WH/f0M1B9thAlv4p
mMmX2csl8zixtweSYeSwEYVu5uCiY8tFAXSkKv7icwZQSFaO90oWnWsGp58T9WJJGLczMhA0gxKH
IaRkfZN+n0pI+hh7HM6uOzUXfeYlXcSulXkwfIjTf8f6es5GQjkHpUlUp1y+oLvzOcKbYpcfAZ1K
2871/0QgIGyYuztRf8r+Q1wwpSFRyR0sBq89gYniLkSnu4BH5vAa0HI+Y0qUpjzQv2ctITrH3il4
fsQxJ6TMjeVRKNkTLLR2ysIq3c63T3WlG78llD7aCMgCH+qCDuxmtiY8U3c6WdsRUNEpVlSLgAk3
pfNK51BBU/fjfxJRCZ3gYdox3osjpveAR1A7Se6nGgfGrEQa7Ud9aWNAO+1sdONcZ+I9hfdtXByA
2GfiHk6Gl/0QPRN06R67v18xoKTaSOJQqNX6I0bnDxcOtLoX6xwaso8J43xJoDWvjdA2x1xxl7BE
fLBn0/LP85Y/8W5AkuLcmyR9zBr7DI3ty7Q8hzxrBVCSnl5XR0dx4yYAc9d2PdXnshmg35aQjayZ
wVNPPvg2EmFwHJMMaFgNrcsjz3e/1iYvKTi05LI6KvpZDQdxlTbMdAeEiWqRMXM1tmCRO86QKq//
oKNdO4fSGzio47MsRn3g+t1f+lYH71pZhk4usUY/gPWTmHxkeWPe0jeNPrblJaVR6ZhBvyk6km83
Ly3pHNLyykd+4DJzEWl/1+mIxHXSVe2vt9mNczUnQ/+zu/xbbQibQ/TZqeRMkUUp5HYRTyzFsc1x
bhOqmHHwLTLBZWE1bHjxivgDEUkcqQfCwV1Q5VML/STbvY7ekePAQw2VP8+X/pE6R4mXIc8TPpNq
D/MEiL0IvHbi8KkB+p2SbputgboZxfmJO64GfMgni0kHwEki3hREwyAcN8XnsuQQIYzDsQGbXboW
009tuLUItCbfou38KjXarkNbMDovM9yWhr1irKd7xHYm3ks5S5UjL9Pn3w+cTzcf+X7YngXq2YAV
ZGwYWJTBnZwsbgeh+k2sNBWZFNX8sh9QyDusS8D1LyQO2q6PJKowukQi/b5xF4zdtQWmlG1rNWXp
m9DqJY1PzRf5yxVV8hCCwT3TtoSA9+AEl1Jxl5B0BMaWMUuCFk8oiq6o+KuSFAanypFHi49t4vft
clsxYwWTJg5ybc4EuAzFKPgeGSr6ysnQ8lD1v9z4DYoifnr5RkfQPQL4mVywRNNgZkx8z6OgyFG4
qyUDeceUBG+UQ7zG4JMVQwDo9G8rawb3elSGmqicCKYciWaToZpIOR2Gb9wBS0XraOeFoNuBoYUB
WBVn3nD+MkvpEc/kJISSNsVyyx+YugRjjhOAnRHtzdxEsjHL/DnTdZkCS1/vDZxnpo+Rpy2t0bRj
pKgEoZsRNLQPoRnJBJSG41G7BlMkwY9S76aN9q8z2emmfLcg8ebT2NuAHGShXlmBr6o5ZkKDtVQJ
7Fd8UPlr6B8bdZxfbRa+lK4JIpZfK4t3x+OPBDNJo8v+hIn9dks12Tm8PJGVhWXR+n4eQRyX31Fp
88AVabKlXbrj2sXb0rZtgDV5EmTuIKKx2nlxO4cFLf9L7bJTGG9er6l5dYlqpRdC9c5y7kKZFBrP
wC6ssDcGe+Drdj5F0TRva4IYgChx90UiAQ3+5hrR1K3rCGbD/0IH2jGVxhCC7ppbsjqxWIx3jFHG
gWP/TiCJkWXksrngjvVt6nbMZ9zTCJ4GDyNrRDUzMARrphUBHJJI1eE1lndQPDluh/8MMWULoybt
fnHRWZdxlyCx30UdCLvK7V0Tx6AmAQAgf8cv0rXo02h4NpituhYFVyowtXnfY0/iMPaWOQiZ542s
4nCSUqebs8wnrIIxKKY2gi4v9MtE1JACPKqdVIxglG4nKWGIkjM4/0bsceLyPcyRwTjdOhgVP/EX
pCDSs63sXcOQGLURmdLPlG15H8sMHBh1bPxj6fJoko+UCSXXjA5k/g0Z+/23VzAXlX1+pffsEpJa
Hj/TFLGA9VUCORPPlu5aaI2kV/bMDapeypRyaed/UMSx6fG69wnJ3YRYwd/LtCEOoolgPsZM87pK
Am7M2FOJZz6SvJJldozWx6y7XOjmQXSfkRD/LsA2uqUajwh5Qh4lH8Vm73ILPtxGTM5FzHE7yVdX
Py6+qGUmTV2U+cgH/MAXbI9bFBfG5EeoStTz9U68Ik7ibJJkoshERdx+FbfT+s6W+FoTgMQbNDAr
n+trVxa/QtIOHbuTWDuqybyAUQwRsSSDBUZKensyQRldtCbTfKgjBkEM2Vfg4KlpP61oCiCkj/4q
2P3eDCzbu5bYr2KicbuJGlRVhQiNzCe2AVrNJVRheLBDOZ5zrpeCFzBWyusROPlfJV6XFWgx+dSd
krL2rXs9UnkwajdBGYXuLuOiMGL3uMzY1rlNpjDiEr4rVQWQYPXcIGAS83HHvivitBUo3EWCh+OZ
/EvtaJnvd5B0/aKYlv7JORdRvUhoh3XgB6fyn2KCuyjWEbUltykRn6y1Me5M/pWS6IHQOl2EWttl
cbSfVIjALhyhoElr1LSly6ptOI4O71Ja13ZJHWQVoAaY0i8NoKZ2IypdR+1cT1JI+7sAG1maxsLc
gAV1F/CTHgH+2xZjQniHjLys3I4LXpnGX7+39WOZ5xdB9tIhPrpvCfkmbxkdQ0dmqYsG5J8NGwxE
ZRc9BmypO0/Mvc9K+7YR8U2Alngu0LdMQ5VFoTLFTVHhP/SITEl9YZzonysXnezbbLzEnz2CTpD6
71COKy5m1JGOQpkG3KZ2pBh4lwnrncQOZ7kMTIHfe1kEciEQFr93mZiYUjQ7te+tjSwisUwaFr3D
Xb/uZMkG3QwrE2d46CEA5GYv5LXuulIY7z9G8yr1t2xEsQT+AwLR/tE0wjfThrkJa/3zQqK6BDjv
YRYzrev8I224Jmj4Iyb/LHjtJBKP+wtuJeFUC5KI5KRtrpf7/tgrT1A2fxDJS4lQOCWXLycElZo8
HF5rC2fkPYQXxrh9c1dRQBKxFLSL/tpsiWoKkOjNJFV8j9xgO9YmGcJv2DmbUd6VxY1RHhHdd5bN
nPHiYV97ZM8O5ZCQxNUp1g6eBZhLFlfCyatgp9Zt9Z/i8+VI5ugEL6KkIxefHNoalCODAhFX9lYn
035lStA/AjB7emXU1JvGYXH6P6kWYNy/np3FxS8HFotz18ZR+a176EXR8hhvrM/tcnrSjAyzaeqS
dfciIAG6S5lyk9fJq6dp+p5luresSFofOE/9kjttRrTYGBwUiXjRqaEWZG92chpUsFqxxqQBrVoz
D0yJDiTV/2TVKQafnYGL3bDmR8KtI24ZvnNU47TgXq6UK9N5UupzprxLy7eCzCGQuvoPjUp1jHlL
AQKJsyN6jJ9ATS+RWb9bsklwvLYa9SY9tYDnTSPfb9KVgVCH1P3mF2kJ2Oi3QWe9Z9dBysBuH11D
xaG86aU1vKql9W1/upukvfDra4L3HieHePwILp7IC7Hz+buMZREqzzmMWnFAQooya8FMtojJmbXJ
apqmJKpihkmJov08lJte3FthiIDgHIKJseQOLq8j2b/pAyxgYmDMk9U1uJyMx5dOLGHaW12oe1l8
GTgrlJ8BK7WkGyO8n3jIthuepi3GlMJOg0UFnB2s7ytpuUgUVnzWaotZdWMSU+GZiDMehz/X9Gyl
P+uvxfu9u4XZ1AXCQ6vtrZuWJ16wZttkZM/1XGjdOcIR4EAdwloj0ayslI3L3TKEwClOv2dFI0Xu
ALS4OUb+G6sDyTIKoyyaWdsuQAQHEZcQxIC7OSTpRrIcbGwahHGjnZ8AGnAEsmoieNsfP9Lst0sZ
c3sBGQ5cWwCxNaCL4WygbuJ2iGUb9ppTedB64Rz5GhkNw1etjcjHrq9/L32x11XEG6IjO43r0Ef4
9Tdn7tf0aTznt//suF5xl/OjYXRPRM9XXIRZQhs4EwkSC+ACGOSqBXcgjrg0Q8p3jQ3LH3v4Qyx2
+PVMkiXDWK3AHIXZwKbAxVbDf5KyFdqOBm294sr7PiWGFhHCL+NDdCfl7Og+8vw1IEmNgxvpBrAh
qSc+8b32pn5v8XrM1looD51R26ZAAHyeyREib1mbWBKdT7Vq+J/LIzs48I1TQ68NhgF70gTJlhJL
4+bIFMOCCPWIKh8jUauXybm5/TvzUYyaylzgMO7Q192wQK36rTt/qCZfaNDedGx9zq76pRFYcEDp
vcvr1pKi5rlOCM4VvmweaGva/9ZnEV6Frzqfm1CBwHycw/7V2djFF+gI9dGb7dw5zExrAVANyhpp
JaUqVhlCtiu1aJKVFiv5lgHR4sW0QgIdoXegA+HiKujDc++0Ov8J9C2FWQCC5OKbY5z3Oe5vxfmR
qZhCkGtG8i5ikwn9E2ft87ARRNQG8HhBROeIj4L/iHWxowSaNObiiBqoqlf3HVHmSKUHEAvSJNVo
XpZ7MP1ILbgl0V/P55euH5MdTr4G8NpgIpi6XUrNOLpGAUK4r54dVmBZn9dmbgh/uZpDErMlKR5N
9UB1Sy1TzlVeUWHpOl7FJuQFDJSsL64mdOZ8I277KeDdXpOGKLoO0xUWhhBDYDOpbkJUI17reMUb
g3a/Du/lqex//eARTWLQ1qgU0v8BQDX4oHDzXDn1I1SgN86ZY8YFaCUkQgAaexyHiqjYm8voYg2K
Z78O6gWWf5uSABhcbr/qNmDGD2A2Q7jjhG2osTv7cYVtBRrKcjWf0KQogPHZ29asYEjDuzgJDiQB
y6/lWrGORunYqFEhx91ylRivtjBn+qPB3nhO7PPIv0KemvBc9ELguDdFYqL94jguWpwxaA834ZrZ
5eNu2rs3u8ZjB0zvMITk8cXm9h3Rpt3VqToDo2gR5Lkhxdwe64uGlvlHlfLHwikxhG2h1MRmsN9n
ihcOLOWaSQ7913+/MDp9nJjIsC1I/cHzfVcVo2anHUIWK2FOiA4PzhQXDDbejO4EJhCyx9bVsLGf
JajerejBjSb4QC0x3kjAqdShjR7C/wDKgTVSIPWBq7dhqboGOWC0Gd7Cp1gwSN6OOEfx7UCEn7o0
UvWKExFQHHCxf3BNWh2K2SLGPJNjIgI+fwbs/yGqwXsq8p5D6YXyy3KWWjUV4E10vDy8nnIIA4PY
G4a+XGdcTG8UiNfGPmuY22S5cdsKc89SoW991G4XfyWyfVH2CuLrFXL9lsmkNzE7zI8PKifzr4C/
YE6PwfFdUANxfNz5BfAB4qG9z5MgtNPK/qsBOB7bK8OWeKX/AlT1Tcc4PVPlsQPrWwojq6Mmv90M
aay3opRebKuD53sGUu8jTwkMbpplxiIVLYBlFJiNOPMypfcDqv5RjGHAEX38qz7lolY1TaU3ze3D
0eP920Og66kCIXxg7xMZVxYHEd282nLQIBjq1bZKgRP9ZW9IPTVA1Itdh/hkt5PWd8ZMTTAAjSfp
NrmfdiEmpHsXtuDeBHwMPz0CUoVIgQnTvLrF9uRQmn4JYmvDE0GLz1eJZ0r73X6sfAKtV5sBWSyg
z/uX9M8OvqJx+f12+I+SIhbXxD6yG1O+rSft6v5kqNx07UgPxS+YCgi9Qjhugx5YB1PiAabmzI3R
TReq8AqIh0zDv7YEPKAr72mRi9wASMpM9FOf8Xyd27n0AO9L4kAND257Foun4V48o71rDf+oJ4I8
DrQlpYed/npcNvI2JpgF3s7gGGNkJOrLfsP6yya5cXHeRLX8UKIcbdXaYlVANPjkGNi5XM9oAxDM
QX76kw2YLZL+lOh9/6yOxQxZ51FGdP1sHuviWvGqRCnWIShHSK1Mk6G0NLe21utJWZkV3w6yLX9B
PzkTuEnWoKjwH1bYFxCN7O9t8ZGT3kHhXG5nzc+Yjbi9uYDMJXFdI5CR+rrxoeks11Vnywf1OyOC
vEbwnsXg5JHHll6843f55FqFIbh4q4odfiY5YcxIR87CQYDgQNyslBI1exqeQ8ZV24oJ5qT0fehO
Q2FPVbpV7x2kyF+mjXcAX+AVyIzW3yQsrn9cOxdEoHBeYOIaOc1Nu+jBYGtaece1FHEt7dbaATvW
b0lCSodw7Fak9abwwXuFUo4YtjVyx3agDVjgRtn7eek9hkvvVWKRTNubxcYhiJTMLPfasF32xBXY
zCdqUHaOBufhwivF9P6wYkP8jMv+dt7gy1nNeVl22l7UKxVPmcBO/wwBg1x2LFAr8NFtZHN41Kw3
LcBOrrf3EzCCcwxITWXnEQO6QRXvvbQLGSdxEawLJTXKHk36XzHELns2lm9Gmw7TlMEPlA1o3m/4
hRJpnVdTdCuW72EwKRfobGpMWgbL2ECi3hWCc8djXyaYPT1EC3ZCm8zDyXtVC0Sfu40MJIQpWM1b
5DJXh+s407iJzPhmhWz+SUhzIYchelgM+hRp8eikFwDH0p6/oifLpcnEB9iClOlg9bPRr5xCxwrv
4hD3FPwCEtR2in0MMC+J4DWm9dtkZgJk0djGjbz8b2x2ZhfXhohbUhnHML03XgdG6J+dcYNWGxEU
2ag86liG2dgaZmlCvEzHCOn6UufmFShrPLjObKYmovHPS0ebCF2NuowVcPiYfJ7Cv1MVKUp393pV
Hu/QE2gXMa1BxU54prft3HTfVDExvFZIalibof+Vv6fJXgyF75NSc1lVKxZj8u8efN9xjaLccc/U
7eRXQ5fn3VXsCIgKW8O9pcACWnjlomRlRQj40+8tTfZFBvPSbQENBFB9BALUbi8jx9K0jmtp186A
3x30/Qox3t71U4lhMtYVlUSKzbELgeNBaGzm8R63w2zLtE4gfac2Lwc4jJOZcWo6ki9MVhRp4l14
eZ09tc//hZKtRABQT7EAK51SvRuFXSX6/l9NnuMf7ljmKq/EWYkm0FYg9Go83LSXb9c4idqwHHip
wLWqE3iIY154lVlRSFL9+AHn0fswBC9V+iNtkSIbfXBV/8NQxSOVKPNxbt05DEseDwQfMyJNLyKl
2ZdM8O81winhT8CR+p0M0J5D3Q5iijNpeHGookxcJstpLkcIUDyW+yZ9f+KcZytdiGcIj7t/TAIX
IopFpj0IHtuKx3KDBF2Y56O1XODJsixbDW2MNhyVBrinjZgeExAbVEwxdjKIDRLmNeI1ixNdh/Lk
jMzH5yhruyuhFMKJo5u+ci3xh/Qlod7mfg+duwyPfyvRxldVxRAh72o3lMowptg9yiHt39xmykh3
PE+uaz/JkI7X6eGM4LevtrsNHqvzvYjg922J2uSeglSr3LU0NJHIZWwh8UPN5owRpZxkt+Mqzq0a
K04QXpDxnQHSvayVGMBYh84SaxKLYgnudn/b6eVey0cKXSwwC587/u8tiBIUl5R+Uro6xyrpy9IV
1kevBqayx8YN1eDExA2SW5AbIFVRccoxCk1EDHe2dfN4xMRNbehBBdhUWknso9OX5aNL0/9vHbJA
89oG8wvNsK74DdvpK9c++5V9cAPar6V6iJ6TY1I86xI7g/nzP7ot6kV9OhhConurBSfJoEI9h8xT
YRuGYHvlMtyLXG/+lH5tE26ILEYirsnQt4rwXU3Dahe2bIxV53uw0UPf4dPwR9yxYEpCDPpfYBD1
x9q7bpZ4sRRVZBIHncqeNif+cU8Xb1OowUVi7eD3uciutTTwbxApllinnSypmJz9YOJSTKAiDKv3
0AzeYkEzUU2YUdMZe9AqIWXXWCA8x7x5iHx1RWuZ6vCKtzPSOHGCg/UKkX4BMn19xBQnw/jOyCk7
Lj3XvoqZHQGOjcA9KWqZukfpWwr3N2ClHVS/M142ooCSH6x3qfljBO4JGfjEjes4M0l1UhTf1WLn
pTOoGWlG/jcyjXlsWXHXwgQeeOuvXX1K86MBSrwxykRYeZR85lljOF5J3XLvmDpZvxIyc7H1r777
CcJdC42I4TLavMVdl/5NDgSUXgSCcak7AoUs7BAoEOXaOKHw6ls+K2vrE/XjO4ivEMzQ1n3vknnf
qnPzNP8asR3vEEHm0sv6Nrx0hQb52dCeB9oLHt7v8xQQIiMQuhAmjOuhQ5lHWW0YtuRHhXIZzglA
g9WUghORCVmo66+Y5j5WD2dXeGn6Qkp5FMx8tABZY4j6WkD4bl3Gujyk6nW7ESPBu0hxqBTfBnW4
QXxLUBaklLCHv6qCo/8Px5JCnb4/FGzHAKxd6rGDppGeF9k5cjelnCbCxVv2sZvmCdBaAXVPoVLT
RxPh5KVBGxjurnrcP4KU0oJZqfSrNjhcU0B5SedjbFmXoLaYotulinAvQT+XYcePNINEEyv8CoCM
3qAKTmGCGHugNpHfL9AjFp0L17DNVLNslAJ7RvUG4JtXSQ1a2FUc2+rlTeynVMffYGHove60/dKU
C6wuQ+miRGdABtxkXno/vt57ma/xOT/W0kgU2mpDHaKWAQOkyMbIJl6gN+q5PO4LcUaXPKvrMv5k
Q+Eer9aW14ZfcrJBNdUWgUh/T1aUf8FJsw/ICXAFon5Yd+KXvtakrTnTpLdb1rTN1mguCvGvOTOR
jpQiTDf8aZToBd++YePvjXBJLAbPMSgxhGB/R9QDdnCYU79T/9QLY+EPAK5vtW0QE/9fvvZ2CSgT
KOtWCEAlrYPPLo3ADmTevppSxzmT7PUByI64m8laJ7e+SL/7QmfC/YCy6vL0CGUN31bC9IExIrSJ
f9dgUYJOAkomX3yDgvJ8dZfR9VwmvmJjzhyIjfUmGpr06WArkQu88UFm2ZqNmksc2DZHTcUijPNG
f0/HZC2uAXuoUhFM9Lr0ZX7HpjQ0raX4KQMdoM0oNg1aa9ALjWZArGlyyQkGiqZbwbqaQJ2Rw/As
S2Eus8WVN3P857+jJ29JKSAojJHBODEJ8hppvRIo40jH1gLv6OiW1lApVek/IpY1OBOtYQc9WAUo
lxlPdsEuPaq3hXmGDAaGxeE81f0bNkCKgiulzMSzplaYdf++uFoDX2qtqI4t0VpTPrEksfz+YSlC
ATRUuM18H/vg1ZzZicXS1i/DE0D2jPDXRr+ZvvDWkl2A2GKJnS8X5gunpBLX80YenJU7pPjn3mME
QUD7g5K5cGwlP5n/8fEbu1FeaI30ctS9RAEAdOmDLw0ykC8IviIeFAVii2MCRPMsQsGbu/VGBAVi
rAm6x0Pgz4tlP+eqVIB15XAJCR5Jc0/xAieQax3pqBLMeNxMveiIaoLpeE3/LhdMj+lW2vvX3yK4
eWq0v9hYPFDfe86O0Jujj/R453uaMdp/UPMixMquUtknUAXM1ZpXSpvxAhsBbkIiinRymw5CFQbr
qO8wSnOLuazCSUE3G3Nz9NBYU5Iy37vOmOvONSHFjQJZuA3L61vDqmINvK5jbpEnDRuuMm0RypmB
NIA2e+c1/QQMn29a/OK4TMlV2V+YpHKMunKo82WhVLkOoAh80NDAfmpOiGbuuKHmWCMbxjBREWS5
B4hrsDzetiA0WilWACUF0SNwlN/U9tBi8L+cF5+CbKyt20y0mJsbo4bLxWkFYtK525GvOl0l7YOa
KQOc6UJhnK/kwr3z58LJxwxHu5Kl4yOGb4oDeYT0js+oZ+8ugYg7HgNZ6X6oSsDd8H7xZSUGDPYa
CvIansA7XHH3mu7/gE53Tm8KotYR7DgqGE9EARs7kNuYErflhHWkb0T/VrIobFcw5VZ4p2mEaUam
HFnuI3miAap21LP/IU7v+hl38ktNSsJA+BrZyj1XtGEOwE59hRK93XEyTc6qQquO148PG8g8aU4L
JR/EWxfEzAfBa25XqgJiVPu90zempHbmEjVRIAdQWKlp4tKrG21zCpFG7Vy2x1+aYqA7g71jWEYp
dN/D0h5Zf5SMWJsIgXF/dTWcTXyPyQHdNHEwTCGYVVlZaap7oenzLPCY1VdHf98XpAvVfVISBXkd
BnfxGLHdcLJCJDOEL5lroPdOJlfrGJLTr0q640c03u/OnBOZhWwqaWBS1V8d/n7oRpiBI6DcPLLD
WdJGKalEQ3E5oF7DMhad2ditwP1aKkTFD6jiIf6suqis5EdfUqMdvqrKdlhJA63nGYIEUR+dy1PT
ueUrRHu2qtHqR4nt7QE+xNInbUEDHw5/udKODNuI4ECDiRCWIAMdlqMaCn6p2Ni0nqy97e7hcy0X
i7lCfkWHssojqO3r/bfUj5zc+riY6Vu8RcDbNKSsyHQPjER6/dJ8HL1lXoKz9BmPrqOWwPiLHyr3
MjB95X/k96UWVvNFWAbjvSbLLjTMWvkx7u5NHOEe5SAJoTQhw3ObIwcdEnAlXmzz6tUMoWfg2B7e
smf2mvKrY8Fd3zlZ7Uz+vKPFpYFT/lrHn1tyUJRg1r/AIRRdxCqE6XBdHQLMdnaJkUFK/ScVklQS
D2aV+4Lo/c9saSgDTY78r5Sp6MmURnIpnuAVBTObg9CpvpCwAuQxrKTqHaAnEWNZO8fNlAma2uBe
oIPce3a5Z/H6EHPLhfMMYf0D51HdJW+br0gMqzjtFAn8q3LjJ1R6JT+C/nKVFMnWo3grfZ1S91zh
AZ321S1/BPhUyKCU7H0PL0imLcxOkgHLAoOjXRjVswPatDj4Phb+SRfr2ABdbO90Y/A8u/ZoaGNN
pjj+zKKGnuQkKlxDb8Jb/eeRycQcOMVTBbX6Hk50pFUfxCa36Mxoq6D7azXA7B4zQVZGop+RsyjA
ZonD0HGF5dMoprGNl8+dMVjCAeqKhRDVryDgS/hHjMppRYV30ul5EM7C80LGQ0O8tjPfQc9nM3vb
lkpOfnNBd4AaAGUbf7SGw7cOgGgX/pQgQcHtnPbmzgMtSMQqtMf0UbL/1ba1McZxAAUnVJ8gmZ8f
8JFTW7KAHTLk3XfFEE31zXd3BmuAvSGdfEYtwEnFVbWvRMm+5HWsDw796GoOFFI4+AkIRZ2k9SLW
Ka3pITjAbJsqPBO+WnlfUwywClzdWFc13RHjgBJRElZwZy6mhi6gJPi8/upN5wLHZ7Y4B67aCrLF
tak38C6vqqGRNvuHAct60ODhbAHbF1Q59nUSRQ+2bcpmw7+u5TzsCsw0EqNSAVNfFJc0R6mBSA/e
RQoTOy5jC8YzJEcOhW9xsMu6xy1vflSD2IbO4hdYB79G28EMZ7HRvxe+g2fiHNFMP+NuPFiBb9wP
4TMWi7HvM2+vsOMUraGiVB/cJKFQSgyw40fWmAELGFQPUla0+ZA9Ql/oEPHbmms5uzA+T4QF62eg
+yqKzOBrxKumDcSR1k/k638o5BckNJdW57pM8tk3T8HkSVEyWK7176aMbrq5+87ZESsOuhkSKgY1
Do1+Db93hpLnJ15YRlBE9d8irDF15+nYfuLpGamEAjf1O8UvN7adp8QNi88hqt0ZU9tQhGnoQF/j
kTMKefFQ2LEAERrdVOtPvvoWocM1w8P0LlC4CxMsb3ivkaom+UqvkA97fSlPGNQAHXAyFPDDWkWL
n9OVO9V8QR10KF8qfIq0WKoOA8jiGCz2eWFiwOeEMGWjbfSHJ4iaCYAndKqrirUwpLjUYHeuyWKq
EDJVFRTr0NjfnMCEAS6bU9fHUpzppEasE5ZiIwPbLV5d3+xvZBVjMgk7LInUUTUNeuWHWyovy2m7
JC2/aU3ft9oY4mbKm3+t2iumMO0HfmH5cA9YiJC8I0BSfGz0Awyhqmxr5fvmkjz3sB8kgukLf6kR
9/oIsejo7sKlnsvbSxd0P6vZCI16GAl4kwlFtsvqAeNUvbEb6pLFaeZWUHJbkehhQlVVROe7+q+f
iQQAVVeoXTlFu0TvhX3EmK5l6YLGlfvrbQxHmuXIC6xx+UiJZPmH6jrppQ55n5jR7OTXXHEzIIkx
GK4TuEA+xIs7HsnA4/asn8aUo7PD2PZm6zML3q85yYdLW6QZi4rXvxPFKTGzCSZRn3zafX5Xzuxx
HvTiTsMzzv19v2Ag8PMHdBH+3bH4fSlyBrcphGbC7fzxf0Cq5LtcKz+4IE0nJLrwjQ8QKMK6Bs7J
0WTJc/0fzs+vqTOL4ain7OFGphwSTNx4D4lUqA5oEr+iBxPAzETBhQGu9KF+0G//4kb2Z+iZWJ1h
+KN7kJkk7tD5oEg2JZtE4XbY+6Hv+VJkHSaFQFtW6uZ+NQda0eZBGWM5HSdUajJM9/xdRMt1rn9G
NJ84LQ2YR68gAInaj3JWOpqPpgbG307FC4+0R7yZQHn+a9DVEnWNgGe4uDBjQkbUh4UoybigTA6d
DBvqk8wq1Pg3arLelqzLoRt8oMuUg4mNW583I1k5MXFARgILLNswd2mtCM3QCIHl4GZ600rZEEGW
D/Ig9+kjQu/cQM4PeMcOkhBg10cX0R6Xg7IidoQRgAVbN0mV8j2EDF0QdNsIkiwk2BP+sjRfWDG1
5Qi9BiUz/VWZMNhTmmXk/+TOPN5k2q/cliHqQvYQUzhAhp3E5V7L41X+A/jER+pUVyHJeCi2OeEU
ehlZKgGkC+bvzQ3STOshBvfzRB1m47enljJWnOhN84X7J1Y0cjATL579bctcH4ex3fKZZwgx6e9q
bPixspClas14wjP3GtZyp5OzXRDtdk9SbhEPd/4UCy9p6Lbsm2L0+pnicY+qIoQpHixO7n+EU4Gq
b0NUp2WdDezgYV9Kc16tcivVaaBaDiwLLQFIhl5AkuwoyLKPvGToQxALgPkEAbZkrCiC3CTcQPNg
66hqQRZIIH/0DU0NyeHaZhNIHSijpIz53YjP2RfLECYld7IiOlZQPVjkMQZHbtw4aEkIIwlXBe+I
lVnwcVrxm96tPiZ90EabIrowBZiofpboKbe42ZeojtRMQR6zntvCVORulZtMfNg0+4TqLxHaTVHE
r9pxlgFrbuS04kBmmK66DOtPhUFoYdxDhp0gqvw8LjCuWLb3/+aFkpHQ/42oWmrWT5ubLbb7nXv8
Lba5cfUZ/G3eyHimSmxeqS9i3f9FvqsHxUJLOMziY2nNQYnU65fkcscJhGwD5LMIeB7wjZduxn2g
n/Xu6pt//vkSIUjJ2UDj0SLCVrkaU8Qxx9row+VbDUCQvj1qAuAaZXD+kkYQ0ed2yLWu/lkp5MNV
RvBuzc006Lpt2+5bvi9rRxdyFp/tw8Fa2t1MYXwmwViHES/CceJlngrqIUv2dD3gItAFgaRRchJD
97sttdfd9DmcYhAhFu2hgOHX4oX7G2SyjMCX2Wi7e+q+Jl158CWjQOh4g14r3qxsEa5fTuLjj+HA
Mk6QMPuBgCNld6h0ns1x4OnekHzPGCQuDONu31Q+2wb58W9rSfR160piW4AQ4J+aRvEqqNen1sLu
1xC7FgI8cReBdQSEhUkBRxAYRedoKzRIafio0WJPoYYmsULF6ciwxwoN1CMrxMqz58wihPzqz2gS
Ro/4Vd3+OLzvvcj35ZclsZVJ9/u3ef0mfm7VTYGPM1d0rsZtFYsqOgpGL5TvVNBBbZivtaS2cJcK
A1KXJ27UUZOIqnDgesP2H+i/BkcupHGs5wVJaqQ+BIgX7N4C+twE0HXfqB9Db5Ayf2lnQOshzyL5
vMG5GxiX78XhU+xK3SyxAVC6e62u9XgWnLHyvAGolar+BA1FCoL6uwjeUPTYD323LzH0o6CEtsBZ
uNAQegzb1UarwvXbXdqsAA4rivUSEd+XD3Ih6LYWbqvEDdZ8rb/iSeZ4/dRjRuWrifjLIWHEDgyf
R9VV4O7ZbaeUdOR+fBu8ZPgapzhVeJXMr44FipD3lWFa98+nx8LMgPGxM6/lLlVm4xKy5/tB8FR/
uL9Jl+yOR+lJW9bm4Tl3NQddW2W5A31UeoSV4ftNDzb5KOrQNF9uN4CY8cI53fc0nIPR1VL75Sfq
HdwhTsgw4Zr736ShWtjys2JutxtGePaMc/qW5NVu0pKbTelA21Oyyx1LdOoaYdwz5mc9UzfebbFQ
wYqqtttad8oQ6/HwPd7/vP19dzws1awW4z66KjSElVWZkldBsUAJ65Hd/lvxu1slofhdHzYBuT/S
oyTFPjUF5OWDLkxXJk2ArrOWH/g/l0hdaRkBKgjqPcu2i553bW1nEyGV11/B2Fcq4vuanm6MAyVn
L+xWr5ejwdw93So0XRSrE/mNeviFKciDGPyPI5NfAQoaRpxJjzJpQVEL4Nt0W877DChA/0vvqqbj
VKQiquXAMN683Oj+g3hpamKiLmi/QQdccnlOMaoJTBdNJi8FBSHSZoZI4l+WkUnwV1i5F25p9ero
l1kgD+d312y14uK3hJCvIn1PkBTBcT4/pEG9ipfFc4SUjviCmK0nVzHpk04DLiVzMw6QW5lmddIT
7gWLG4n8Eu6gG6a6sgORbMpFdrp/weLXmPBzOaD2eeqRfQMiWlhQ1brfKeUrsvSNu9ZhA82MUhyI
EIg3Ax7vmOdgkZ2LTbtNT8TGuR3HdLNZQHsKjndvC9QlKHHCWyuVuPPiOsIKcvxJBgHl/o0hAYjA
/EOG5b5qIa7CQJ/aYOXAUIiCwkIyYxRqVCkBJs+oABMOLSpOtfwE3b7BMUWwAvbPXs9cghA175Jg
oQJK1levC+nL+IzRHz7b7Evq2vRBrwS29St9HObJSz/MC3/B5GvIbFQqLYe2oGTJRmS4tWsLdwew
D4KL9jzCWxYpZUtRfaZ4IVQo5Vo+jOrA+JqZ8NpFJPIPC23b69HwsJqayzdF31EVxZdKyJ660ppA
g4dVz5ypu5abwVjhyrZIqnmNLsq2OGCI4GxMt/ZPG5pnQIUA90nCPm0EA/mHGPkMjYkgNm6mQdbl
Zw9K8oJXpKtt1VtqcHg1xnMxpx5fSTNs3fLDk+FN/IwsllSupkhhz78NNy3CrohyepojUBLTY7Mv
CidMmSqyqIEuuBx0DPBI5aVAlLdXaPd92Iq4xJmzOht6ppCzzAClHMc7ypnmsqnWnP1XTFIiTC/6
wS+yBTcIJUPzXUXkWQql8HHJC7wtX/sPQLshvOxX2j8pIN8mmranQcCh2MTvVXwa9lw0QG6dXXi+
xdRSW5dnKOhAgZYMsW+AShpAkLk/endF3VsDv2DthgQ7CoeiNQRWwxcw89tPUEUPx48V/EMvLW3e
/0qUxCSRst82Y+21IILViuZGF6Mi7JaKlG3d8I+jT4HpdBzBlhNoGQZtS7QHAzY3edL7F/gksVjk
y+p3amznRIaI9Rtyv6sKOuL6UV2Maxn+ni/uQ8bhiKNyJi+Re3OzVM/6RIpHwIKBCoczQIFRfPry
ftqeXrUIgop5nzBbLOnojwJaA7LBeHtwRUxjUsBIwkR3xPP/VamRpnt7UthTtE1ny6kEbnfF/rx+
B74bpFNrETFcIZTP83q7MSU635x97a/tcW1StQKSYdi99+U/jy/Gpgw2Yt7h0zgKsgq1na004Jkg
+4mAiR6s2Nz6zrinRTJfVyWkItL5xbkybTebzqaxFBHfl35tJKLn4NxtxZBZYvsUErP12YI0tOnS
T0xbrv/HewYsoLzlOA+SJR/Uf2IyQ5Sd3SWN9MjghRJYpsJKt1xDcB87JwoT0INT3f4K2PIkcun7
noseoA7pFv9xpD57J6ia7F1lr27KZgjxKz4PBhZOmbJop3K+HGq9rBRzJY5sK7TXib2exdIZdExe
PRvPc8MqRUg2dtMR0sMaMkOHZKBZ3OMQzkJZo1RAg7ljhDV9i4veRgN5DPLyZbb2mKbAOo3Eg1QK
b361gCqQOjbB1SRfgMeXljiYDl2XM/enQTPlV6upRbBPSTrV5OFG+TPw+jIUsT6SorOeNii/Ga1W
yrBT7tKRMUtTxHa1rLo5ZJwNRo7Vw01Env3na1OsUibnMGu2ftwj/R6hAlTPj37luIn6x6VfMx8F
hH1m59+i2FNAd2m/tY1r/jukFXZWtANL5Nk3gVgiot9dBrFS8/fBlqEO7xpO7yu+DdW1EOHh9LBR
JBOFmLDrPehkTXXKGReS5K3EQXhyRemjymHRlDfVeCETjmKnh/LXkf0WwVsOLT3Rp+kTF/GX4qlW
8qD5ZRxPfoesgCfIw29x2Cje9eevVXuxVlFn2JTeh/eLii+YvrZBw9PkQa07lZHvP5ZipWa959lJ
Wm6MVJEaxmb61G7f2tkw69P+jKk+LV+yGbxj/6/A9ynA0E+399hGLpKteJohrjeldSEE8ouLTpoC
PuaqfStE8FnV730KyPSRBXm3clJWB+hnBa2o0UWDDHhAfqHFyFAvdg8a4mbl+DYtURQDtQIaCmUd
TZwgjfMa3pqOEfxqUKInpl1ruw2fI6xzc7dKKcrySidPDEWcCLE3JlsiRHpngNTFsnCCT9zUFGdl
8D0UVj88iI0OP6l+Kal3A6O0raWx9Il9afHJycmYer2NDewQtZWg6cI7STkZeH2EvdUDXbQGsZNJ
Ph4trTDnztgOpryUSwOwi306uVjpKr3LuB+rQHSlkZR4SPBqpar8YEs14bMEJlmhoykoJ6dTjKoz
MIYzpb7S9i0d+vfVzGRKQZT9MI5X2G6SQHnl3n4uuE4Vbc1JNscZ4LLAGj8cS+5Y7a+kCJzqnbcM
ZWl6QxyvV8KvkR9ADYdR9XyHCI2NhF9tysfZal/cmcZ5tE9T7+4aaored/KSY1xSWqxNM8Wj5Wev
gBk3E9+sP/nVUwUp+YjjMmLplhLTOOFiw8sx/Ne3ItBHR32yd0uCXsqJ3gVryV7LpG7uccJom0Q7
9eDCcCqWcauzNECA84jwET4kYO79LTWDkzNDdkUKdU8mYtimo8iRvz0MfiGFbhCH4qgv00adAaXE
Rd5xPd7ni2PW6DQNsT/5YR9p2SJ28yEzFdC0hcnlBhuL84gv/X1dK89WDE/UAGIcZ3bJltFW3r1Z
cxymt0PtAduzGvRPoNYo/9RzOV6yMbIcfNWG6ldTbtmcZyfdqz1Bx15i2KcWadfw3sY3WZ5ETEBc
p16rOsBxltE/ekszKulza8ALDAcyvvVeoOmKm5QbwZbxjkoLrxUBR3awn93Ft900vhnt09gNBq4i
ggY1DJh6UfUQOrNSIQ3rTNJir3OmHTQlKl33q3zz8rGjv7moipBS7wvPLOW4zxC+KeaU6C0pFYm5
aeDwWmn0DNyxUW8jzTwNWpKf2AYbej3D5U9f2mnLZr19hSOsj49sT8KJGt6FI+WolJ9nbADc6OgK
5FgaUlVuExRlJiygruev/EukY1EtPa0UmslbaqwPCcsxBtdEd6Bsu2cME3RKl1rVO4QHNwTglY3c
Idmxs8GJuasd7Dj0AONd007XugjHQ3cEZ1BHYl48critu4s0/EhP5CAbZW+KySB3GKlm2RydYh2J
Y1RT6B9l3SlQ4QU2MukUpwPex5ElaHFNBUWQA5kJLud8HhiTttuey699RuvHfIN+vG/WRr0Lcwc4
Gu+ERmAO14wcO3hQRSk85DMgwaj3DaLTw7NVuOWlCn24k8jUkXNxjenkqYzQGkEx74YUUiyux+Vs
Jjy+XI0ZKbAZytt52/dSfF6BZOkdJcVWhyQ3hThELfVxTSk/r8lsAxMO0OBZZMMRIRH5xkiCqtYs
EZTMyO+PEHuHhyVPY0ZXPb/Lg0GyMA3OqM4TUxOU5fOgSqj0M4DBIYNPqLmzqpGPDHZBxv3flFYa
3MbIjslumzBofPQvWbQ4ojn7TO0riM/n1T1+Prg66M/OReDMmKeSysmWrmfXYH5J7rIE9efOqDt3
WGn4qT0Nn1pil6jnfhsq16iFAT71EJfP1OHBMz1XLr7qnNaf5IcPArxecyPFIdZ3INqf6o5+hijX
5DO0TR8cb67cJkoGxppDZaogu1fWnDKgGvyffMU1WHcKOJ07+BDdfBtGIVd0rHuOyd3jO/FZ/s46
+nO9QYlzmGQLZKHnd0HIhh8kaXgBNRyhpSn3v0xtzguqazqz4U/wk9pEtYuZqEqdnjlzK16vOZfD
P1pe4PGz3Vmb2nO6GBWwvT2XcVWfFAEEWBKMxuVTjSwmv8plS/jAGT2bZdft5gpjkpXdAccfRVxv
q50u1aSpRZxffU+J3R2vOAl9THuNljDnY3Yja2r4kX5k3RuA71hVUW+iJT0D2iHZ2RNlnTWqEHeX
jhfSU0sxSqwLaEUhnbAN4Uiy1p/Zupn+DiVEz886km8WXFuF6ABGiGPWf04+W3d0vFkf+24B3Dk4
Hpde9MoY2iote4Xjb8AH94eSa2G01zmBy8Yx83qlHTRVRcT/w/pwQ2+lNJrRIu+K8TxK0KGwPpPp
ui3BVajXiGF5d4Dmf2Se6oDKaXaKadhHOwtFcwhQKvvBX36iRuct/NqauzNMd9zP7QlrBpHuD5Kx
VFK/lGNgSTWDuYjqVt2zAfT6vUazSvoyKsXRWYcCrhnM4U15ndZ4P+RB8R1DVdd+CtZG2pwZyWQu
iAMiC2SEYJup0cfn+JtUvohMDhABnt7TZ2oaadDRpUk9CAc/E5mIruyQ5cPI8+XB9uosSu6uPyKL
SbeCmlS2Z10e0NvqDE/fNStAY62cq1g2hW/YOgV19Qf+rWyNDhcGaPEDFFn5W1x2fnE3nJbyyud9
iuKClTecZuCsU1lWAgHF9wMIIYArlttcOPhnZJGGaaWiP/4xEPUfbvJyMfusPE+oXZD+z//rM5rc
HvyXsD4a/6yyuIBjKoRut7Srv/DVFCND25KCcQaEt15pR60BPuPo2E7SgSCRAClr7MZdxDoiR7De
yFcU68gJzyV8KMVjhGgNwZF51DHWXJo2B/bajZvxpuaInSm+h4UGFdrrrLbqIh0YP/zWv0M3ZCo6
/K1+IIYCo8tg2uSn7XJuGBD3UDAKPGTTIzriqLr0OVyKns/m1kgAfs6pXgazP93ZcD4cY1QoFYe0
/vhCMp9Bq2PEYeqXjif8XYcCfEZi1OswP+9GQpMqCYiv3Qd0VAD+BbQPGJFDh482oRkm9Z6o6V7r
Sa3trF3kg17W9h0X9y/hTaOkjRSUT1ZBGjptu7yVFsXj/AyhmOyLu4DT9g8ZAyW7SeBnWGqRT7NT
GLL10CmU6r3x6/pmHslrMssWqqZxRwdlwJco3FzSkBN4cVadq2+bmlYhKjw5pXyoXlr9R39zaf6g
YYnbA37N7JfiDIaoTxv3AthRAzvyE+B7JX2H7ydvqeCh+z2OA7jWoEXaYmvpJCtnQl7Y0CMKU8AW
ZTUZWc4nN6h0yYMA4Z7yotJk6ZhfJCGTQ+0vH+KvdxeCYntfM99HefOJLIf8eZ7QPNK7yxLu8tqF
44j4Pjw+hLyIfmpGsb3/BSgnVSYLnxfzZurP5oPKh79W+HzAUFz1opNGp84HtHwKHqBA/e2iaGUO
fJf65TAmWoStYdBFUxDdKAQ79P4srbOAnrAEJmJ+mOuIMfBjz+I6mTOA1aOHScf87AzV5dV2FpPX
/vHcgH3fz2/xiD5Un5r1c4tgsSQv6hAoyfei7sNfds3S2g9Lhawf3SpEWR9VvyhPDjqUIUMcH4Em
PwJwrC35B7yfBx8R416G5rTq+413a500oOdAE1Yb1D3OaRz3S1ug0HxFH6rpTWHvemQuhUY6d3Cn
VJ1lQAnkzklSmq1lJA/wpUScDuIARLg5IVDPpNUGmUXgPflBlMXQNbRvsW8UXdGMJZ0wtPM8xdx4
P9Ys0FJDf2y5j0Ko+/730u5EOq3Yr2v35xeu1DZPl21IRvNUic/5PSnBWGCIl3Rn5DUOUjACfEqf
QUVrpMzd5KSEP9/5MWf21XL8NkzJwbMQKe/HLsCTd+xzC5bn9/rn0qzEsx37RJ9p3yFNtN0ssnsJ
aunoOzbxmwUCYf1Yd9v4wwLeWSziT+wKGb6sMpy3cez9ib/Ot7H7dCjJPZCZyl6XzzGS1SBxUfNy
GCdGRRbJRiEKydJidlnHmfkBaMJ6V+mMNccPRCf+ZIhEVpQNw+rBoxzDRd8vd3UhwLbT1o0sk9/0
dmnweUzL++eBHNqdsNAf4RAYAXJ0JW8FRNViNGK4ZTz7iyZkBh9bP+ITdmhK1beMY7oj+2shxvt/
YC5PzVk+y2V0jn1hn0I08g+oAr1hkiik+EhBYRewj9XqA8ix5uQ2O76RhmVU/CejVk0AIwl/No4e
HT2zK9sNZ6xTtTsoRXdQCdDYncJDIomtZ8LnrUWWez+lVy3QqEhhCmNbiboRqnXog+7avop4T3Rt
N4U1uGCCmbmyWKe3gDE0FAIq3xyLT5FgDbezpg68/61SFgwX0VcCWR4dLOVhZb8bM5SfU4b7FwyZ
Jir8mRVEtJKs5d10HF5hBiLI1uxjp80UQQCnMCjbHU7efNUtD0iLg6GsANwJSoNZvrjznXhw+tU7
hJ5TtRopoNGhiNrt7n+Q5vL69gwbrPWPxcr0BooQJU7yS7VGPugEMglu1hdlZ6o+nVqHu3Fg/fGy
9eqfS4znv9E4HAMjFW4VdtM37Ztl9FksOwtxZjS4a4OAuTOtyoq52TUDra8bHI4crrd44EwiAMoE
hfPkaAukTz2+8InZDFjDgfnt3Q5xPMsuIvvf52U2aRzMD/RrlDKGTwes+oTFKPDDU1oLjTogTU66
eXwQ64a/Ja2f/Mf1V1pYvvszRa2viVswxHsgm/yW/Q2ysV+S0g5Uzki+6PxyM+2VOBm558WBhqzB
l6zxYLFA6u8mwrgIx45Ptk4tRswodcthkMQn3bw1W7Bwk20i49EvGONIDAlaf+tzHuWGX2jqW42A
rCGk7z9W7cb+0RMLwdYC+PL6f0iLH/7iP9mTBrBtqrVWCxjAQokhdI9L7DqFO4gZgy/qU/e8oezK
zbUN2ugXSWzaF8crjUxzhN3unGIk68WyFuv+NL5Rrof8bzfU3iIjLxri93SJLdViPgC/gobSbVGc
LTg1ShLbCJetQ97HGLo4TCYlGhbgdIkdHVQIPitClr+b1voP4PU4rXQuA2N2pCsu8PM/HZC1korv
Ry3svIjmyeLXEV1VaczY1WUDXBbjK5zpPBmFSQdGEy7iQfxYhNzpPXSmWNArEXTM+4sKyRq/6Deo
E8uRp+KMsOokubeYNucypVMVpQnw7InTASrhDxWW+VX8Bu5rgVcEj8fJie+QvonGNnJrpg7FAHMW
jI+3kxQ+gE5max7TS5WrgKDBzaG9N/By1zSRajBmsQzBcsnLGsYMNMRkHMsTBLqraX5gq/VIpElp
GB636ulSGNDnPg+GiXlNDbc3DxIhpSy5HvsDnh8EUlk3SKVFV2sCpRKGAx6MrhKMd5VJhQuCVg7u
KdcuAFGRkWT9xovKyVbN7ll68GnYYTbh1QKVqKB+QCJz3Cf1KpkEJpDjEjueEr1FxjJ8KnX5tsEY
3qEG3k5XDlaj7UlqGjoQ1fZuCPfJo3dsMuGSyDKjcf5clb0lBV6oP4ZFEEOCA3KDVz52secZLxcw
XwvNZNDiaFlo58RhDVMMaeRBogX+BmYl4qzjI3t3sQQEovhhxF21+cOVXU8nBbnYLJ/cclkzxHzk
t4KVZMDjlU1ddtuMORlmjV81pjRYlFY+da35wZo7whrz9DIjo5Z5GFikj185KIj6Y4X1gQISaZD5
83ZawtG/aws/2rnW95jWp4WFa3f8GiNisylQwfZ2CHsafJmLbYVdr3dh0EUt1tDrye51SQTb1Rnv
bN7ebZ3DElH6IE963XIgvGAhXE2h/nr1xc/ioM1F8eqTXjb6Q7AKClmf2+Bpb0P+cNsB8ElFKRuA
DxnkY14F2uABZIPsuyEpcUWrg9X+k6/fvHGp60Ey/2zk4Tu0Ni46rmBsBRtskwdATdoVz5dlzU69
ynQx2C26RRWD6IAuzcB9Dv2J2Vv8IvJNEwEfTsv1M3hRz4zi9LZ5sYD+s00XCGE4EIZJQ1LoelBN
yEUNhPG2HhoSJ9PT628PBU5uHQuu7lQAbtdJ9Oh8PaaxO5OMVg0XGhNwTB1emPrEaSh07iaX3Rqb
KQYk2msF+aDi1Toz3xiTqtEmlPpOADLUzcdC+96y6s23G37OgHFtFVG5tnydzaxE9hVNCSYH6ox5
zNda6VEcLpTqrj3L6QS49jdphTMf+9RM+nkY8uJSa3gvURKCIPcgW4dUikY4BO8ztqN13B5RQoDN
Y/sDmqhrst4QkmZsdI/dhfGCBOIRDpuG153DqUDdKGw5icZeI+X24ChL0F/iYcV3hFRZf1Pjxo9G
JSnm9gWkQTxToKGEzx4v9GqvA2eCAIyG/n53QdSdIq4PBb30nGBATI7ebxX6Cjjlw4/UZ4aotDnq
iCq75WA9jXrzwUu7tkgh2a8xzQmSTqbQF8qDdtXXs6RaYG1SkXm7/hrEk3UyDxLhf04kDiJGho75
vacu064lfMjB7N6ndDhbYnq5Ae069MiOCKu4w0IKqbHWpKTPeuE/DyiWo9hXTCd7HhaYDF9g0biQ
KpxqEG45q89g7VzujRzxQcb9AkkHqVfpXUrlfPguD1uHozdHkifyhdlh3ypf8792Z/YzHjVbUqEm
OWGGvUzBUYvQwDPpbodu7EeaL2JTzqrtTcRSu1yr+eiEpobOqPfLBGIwJZfVzGC9UMCAkWBXYWh9
K/XA61A+b7RJzbqO1JnGIeF/pp3Qe4kQXgnGHWBT8yJMjcqZciD0RZZO+WAu02Z2qIwmsa9x96gk
dVGci6o6GD8zDWN2yDD0zlfAK8jk7+jjoJflYAfVyH1kErJfEL9X01uVpame1PhDiv9kqf/kZydq
sQR1N0tqH5VYxfyvua6Aw8ZreB4xNqg2dHMCGG+WjNJxsq72N74OJ0VMUSu8gegQdEIuJclIKoqm
IwKzjJVmWG7W5oMi2wOXsaFQJIEJyWx89pqF/BKa+Os5xCGqskC3D32NdFBGOj/ad8b1YVo1Hvr/
EMCHrFw2GTfhVU2scE/27I1U4vOcZ3YB0Fd0iek8N7JyujWGJ3NAv6ebOHVqWC2j2J5iT2SPWiTK
5zEy7tOoMfGVRsIRdRAIC4J4sTz7I62e32PoWA8577FmKcu3edALZeDP0RynrlTj3LFKNA2xngYD
+ppYBCLhvWAK2UISJ8fdS5+mtEBZLZk/eXwZnQwIcHX0BzMAVKC3LGxKciDD+3cPNFgtu9P9hr8R
IX+jyCJAWgMHikUG/8HrRlghmCj5h1UiPRlJYYGnU7qzgNlbIrKpCRoKUYacDCp1ZWdp/o77Dmii
R5rxFJe9xIDsGAvHtoc74q4Dj9nVEqo8nXVMF4YqohoZYciw/WzB/skU/BNKBg/5Ktb5PkEM6zWK
jZEBACZxivj2x+AmSEm3xiEVjIUnjLcZzbbH5CC8ZYuBFafSSADSpoVBWPVaaKENPcjO503dtnq1
4paSoBSTuwnRnt67QhxcZyg+4Y7+qb75IXV/ngsWqMzNFYQRFaR0u7UcI1iEu9+eddyYTP96klKG
oq41LmXEkU0o1JJT219kDtQxj8wdQGwA3LhGLeybLCBvDduk1HCMvUMB0oT5f09Gjjc3TbOl5hmt
dJKjicEJUBSjy9rQwEAdkXeUPUrkEtvtIwcHkdrPTFnbvB4BRw5obkzwJrSz2D8AV8dMBcnHZqeU
aFueasrW/srBGLpVsKnjsiPyNnhDMchrFtEM1lU1l244Unl5FvVoLXfNdYl637sT5FVmqhJZ5/5p
qlW5X6PlC6xfiIrPGO7HFHmuPoMx1vlGC/Xi8mNQ9PkiW0MZ7yT3GCResPjcH4We/wHYJvjSYzrW
8F764ELsZt45pdNv0/Hx7LiHJu0Lz/K4bvMXu4ZduZ/cHIgwU9dLRphDazFtRQsPkyty5SIvacdO
/1OHO8Y3EU7+00f/RvAc+ew2i+/mAoKx8nekfvjGj9gLpBonICWPSoDQ3vRXzQufw3AZdqkk45g7
zmOd6JuWfuLcGq+Wt8mxHHA3FkNWp+IyTeQVnJhB9Cue3UMh+3fFuAGbDYiYNcS8qoFIcqu1Zr2u
BKVv72FBU7jBIW+zYtC8zYHMt3HL8kdHlw7BxXDcOiq2CObHKM3VGOFaEysBFfiPOonJqpMxFfSX
6+yPYa34nn+ItNkiCshhRCP3pehRHWsem6+v4CY6VTwN3wTKSD1Ia3/awTHc/qmXVHHsPsULChoK
6EX8KulEiZ2OpEcmohAAQxtcm7ew2y+J5goX0+YaRRh0+GUvb/QcZn8z8j7Peaxhz7zCeoAkdOM8
K/PPh365WJI2P4VNjFeY1sT7HFTnlRtpeiRTu2eRSS3IkmdhUPFryJM8DWH0dcS9wUkXqzg0F78+
2Lsrh0Mf1cgB/qx6YmynLQuxPJFMKUeSkT15U9p2/1bHNSWvdOv0jY3eoprtimaEu9ka+TNcd9l3
6tkvQdQTXPsW3RaWLHjxNMil0b1NTzf7VqrYl6JMDi/mgf47wkA8GAYfmtAUl8Wf851v8X8nEjoX
c2Y76qucV6IxA2CXU6w4rDByEjUpHxOg6EkMuF6mmMVbdWaTM1j3RsmpRk1nJY6sVUhHvQrqbqTD
4fazNl36f/bR6xUzBjtlFXu44G1ks/GrRaZG0VBgcKldwZNegY+32GhCTjQ9GDwblzDNOgr3mn2j
wzmbD0CCBRXPyKMlnXf7qJMBYfE0+SYwmDHWrhTT9ql3EcVxef0XGbb4qUt/0x1XBXXBQAfE11Py
xT/uOOicVJZ2I98743pHRz33ZSGm/pVT+ald8c01M4+KYV2yL8XP+m4knYnTePPNg/KBD3Cg2MmS
fM+CuPeHb3v0HV6CyfEPlkLu/jtMv+nozEB/kB4HsyWRGMWWEl7SVuelLqmcoQew5xevp0SEnKFp
ro6wv+S7brmSK6LG7iwBm0+O2eDGAy/m8EwbinRnQtCSfWy96gqsUQewpnxfdbbxhPkjYniuPxly
4+xcZMPyr05FXqJeiGlpf/uFmWHaGNCfef7zAirX4gODcQLyJrFCYRi2FCnFdm8wxVnD/WDl2hj8
QmKK2W7xUtJml7ucXO0hBZeoaVvuJ6UABBDO7e0qVCtzN2Sxvt6iKaWy8/wCtPPjARlonlMkKkun
OiLRzDnM4mnfyY2IkJpunvE2G+adivOl02dclVqvUqXnRHOueiytsdG65C5u+2aogFHM8TJm9FVO
+Uc0e4ySRPflEieSQ+wp030bdqO2WV2GYAUfEsR/ioL0waOAw3r5x9sd5Hz142KHPjOzD/Jzx464
kV0OuIw69wOrjDSSeNa1r1V1wGZBjuzEMuOmlfOchbNFWzsjZjKI3PvEj30LezfTHBrkiIjYZW/x
/MKOj61r2/IpVXwVzVat3cj2Fe8FeKOomYZGzscduEXUqQBiMRYpQ3T8H1lWqSPAhKOv1vLUwWcv
tLeoXlBkEhEpFG47MV4diQOWrRfzJN0EYa+dlxmqkMfEhyisXnNLCQLBD3Tk6qX5kI4EYDF7YdZP
faUuYVqxW2RjqrMIANpB86rU+hBvx2LagHz2RIqMmE+BLEu8dKjrXX0O6UPC25b8xG31M6pyjILj
TYXmusWGqAvxJjC4VR2LE17eqSD+10+2N8P097kNhinOKetFld86NI1qvmWAyC8JV4hg79fjD2M1
qyXGHRE4VppLutdsQlftEP2ICIZoPaXauYadeHR2RjYo54DFmpLDs7cer8fXfcURWlEHVX29ar/e
98POuQLATBQMcAgP/w/+iE7xp29wqrErbE/H0SQnUuaOP/n5exinGdw7Sg/5AjGmgzEbnIjGTV/F
2zYC4zzsO5jfUVecgpUccid+ZLqd3WiEzDJ+PSeJQFNo4GBeZLMuG15ZnMMYJBrTKE793C0XAUt5
F9yiOqoo9z4IMf9Wnexzb/+6GMuiS/vrctCwsdUu52FSiS6y9NYI637FyYYO7HhFv4TwUMFrXcAj
o1KcaLZly3CE8Vvhw4LyUUHZZKDFXoklyffiM7TrmzlCIfLdzsE1S2WSbaf0+eZbMAQMbn8Z6MIH
AkUiSoxC6qiiW8cnbsAfpxeJrddGrQbIBN/68n/RNQFib5q0+77aj28CiBODOrOwNC8XfoDXBDFe
wrPY2XbLqka1hiLHaORDxjxrOQRkhiTa4J5byvp/vdTXh+q5A1Fy8pAF6HO3MR6ileGekyjgDvIw
xEJTkRrj1WAeASIgF/h7b36rVDOhW5GqEiZUBtApP957g1zQlaeNRrpuDLD5kDsdpBa1kW3JmtFL
frX2V85HzeOrGXaZm1B88AsQud8FL5usQoG224WooLK96Exr8CKGU4Zb0szxfkQ8pZPNPsbLohig
EHoxrIOJTpiTreSc442vkCff9xNNDQ5zkwwCrbj+MQEezkfoKC8itlVUVlx2RHIkXuZ26PJwPGHh
3cD8z0qwCM18oTJUm4oL8cqi6FiXVsEvlQHXGbAK2s83TngKIzgsWjKtE+Y/oVRM2bFFEAnQTIkM
wEsbnf1TtnCmlUEI0suMThm9izcm9UQ0Ny0q3/NaTr8qpacg7St7n5iZew0I/LOhThVqTJL6HvUh
dzFJkyEF7JQwTUbLozH8Vt6OX8Vbp5lOH+SfHLzqxqqWvf0ST5H2ipaUzz/mtmlbhf7575aYSHXD
oO6wqwkf7SDPuAVQ/JvosfcRmh/4dM6fD3qK6Fcijmhe7TJ2Aalrho7mtogXs6Pj3aTYxq0cv+ch
rk1HlSJgf1vVdrWBrSTQSmoO7ONOzzyUidVz0sqEJQg7lFevzFeJlvWTmNAM8c4WZtKHfhIYYwG0
HvFWBE+B5PnwnKcVYPct1V6d6gRW4g0w3IGObTqt6gv6mNrVW7iIW3GOHP5eEpCqphBB4ZfxBDZY
u4YurHG/DccjB8/yT5ZGqZ32T5WAkVTsQFHOw49qGxd7Ep/SCUIY5PWx14RKCWD/jhd2gkuCKusr
MfScn2sXZ+3SACGccJ1oC+dIPlq28XVlMNXaT2vVorEn13Y6/TfIg7g7Mcu81ydrFC8VJgv13PlZ
n767aHpdKmmlxXF0yZsgYjC/y8B6Cr2Zcuo0gJUFu5yxIWFWMVaknbortXbe7eROpcQT86+4npIa
ZoL6H/mX8+5jiCFwlAeywj5l6Gg5B3OwaxHFq1mgay2ozwVQQvREaqV81ErgwZ8ldKvqVCuCM3R/
w2WzJc8QIxxvj7KtHKFRyPhwzU6MxeeucwW+PaEzGB41N57mjGCNkeNhYKTxKgfKCkXJoQl7LaNz
7sfCjNQ1HAhFY7vT67BaV6/WGMoRKHpvulLFG5TQ+HwW7geuDd9WqQjvGsDCUS6ybnV6iOvir4CA
8RW6KrUC0Xi0EjBSdIPxQjavRsGytsClQlKEk4YWpUfR+3Z1B/0mcI1tIHJRh/dPhKPoQki3T/Ts
30BSXEX8mI7MayGtKo+f8VZyL7oGf8UmfxZI+WgQluoC1Qr74BqxNzFUg/CToDJPyWWKyWh9sEGz
Yo2NIsP1P/PcYf9ZNSOAwY99keynpFjKEYFguKIGpDfUNdVtsTPVEIHMxVM6bzKuZas3UDy6q2dT
J9jN46ag8EFRvD+5AIRv9+bdoVETWxeinTJ2PL9GpaWns21KNnQUngVAyUaiPEqlLIK1H7AB0pL1
3gyCBu6RzuOVeku8ff1ort7KyXs4F33dt6LQQXxtu73OGhAXPR/IBSnOFXujBbD0pH1pF5T8Q9WH
A9vyDYreX573zZvQyQfkhAP/LGHo3ed8EMe4xE6pxm1wQjWAQ7Bw7lJ6JcOw01uxBkdidlGOir7C
lU7Tn9edf1Od2W2q0lXroJZYbQtw0FJCTckpQcXnuE3JIrVhD5vHVwF8rQayVzTKLb/JOhySNoZl
GlDadL2+pllUCnqM6u66uz7DWSOXr8XZhDj9xisen3/uQ1SN6s6Gv9uEOLB5y3zlgoKUT/maMvmw
uudhwg2ZPSw+Grjb82FZoCxVZiehxkg7pvJrLB8EK9T5c/JeJatPZXFs8JrrqM/ZOUozqiniH9oW
mFctg9f3V1PxCgfUewdrISFlH8/4yeK1Yz6p9oImVzuJcLJZHhyAzXg4IC38MMBE6J42qPfA53q7
QJE5TGt4BIARjeRDNm6bvu0xE3r8gsDxcKGa1i3qiB3SlowWM+xEZ08xj8gDwNrkSWXVwXiKmlz/
uIwWhGpcToDZZdmOEn905SC6MXmOeB92lJXFr+dLuHHjQNVpXPljD5qUlDI2W/7+ucVGNjH/AHEY
Jbm6yTCxYQd2X84eM5TXK8Hr+lrK3+fL5TPg7wNj1VpRbAyGgF21LfX9DTP31dQpEbzMUXuIKMhR
EZPlZCMN4cJbwhPh6f9xxXsFZqiCVqMQuOwpC3YIpUcSi0wkxkxkR2SOsRwV0qS+69mqFgzmVJjq
CfqRHDnPUofFi0h90wudD/S63NIsq96bhWHMu0TRTpL3Byz1+l5eK+V5cqCaIhv9qFK9udNW6dxx
c1pOjG2Ep/m8bJ+npcqYv1mNGNFxQ56C6s/R0d1wU0lUfCliT4m3sdzjdT00E7fic1o+22j5jhly
2xh/QDLgnMlVZ/ExADGaNfmsQFmNCoHEi/E+sBS2iLMCvgU8lS0tLFX6ZBD5FizfCQN8wUbCNB2e
EJLb+BsXcAzC6iNrcLAPIPVis+sjOnDBvNtVAMc297AxuAYl8dFkostBJsV4t0U5/5f/sX6ct68K
gVAsqpj+GgET8ILJBujH84R42WMymkMULxJITm5WKAte5WSwkRrZwojCGyd6JxNo+imCGMWJUvyq
eZZ2i0GIEPngPP9xrBkDwV+gk26AwvOVogrVg3i3T5bnp8DqcF532ZZB+mkkPouDow2/NXidejyJ
Ojq2gLiPeEWhmkn/WynWG3/OUiGmTdKQTbQvjlBnlxOUFA76gvri1si/m88xvbjTL47Ex3X/0aYp
K+bTE1jWBhvY9SJngpg/OAStLSwx+M66VMiTPoyOEa75/zrNsmXirduA1nV54GOTJjY5jSbGNmKL
1UE0u46YrR88wJCRls3xwJf/sYLaxpnZt7ONEL8lqSpjGIbB3fmDp27NpaKESHjFh3zuzXFUKdyU
acwlc5c0RJwzbNAuH37QsDETke/nlWAO0uLH0Bw4u2/acJOsmibF/IHgZKl25wlExU4vZD9CFnQa
i257ohNjvsdiYm9NYbzjPfc8ea0uNif59ohlBoArfaKUHawNHDE1gHbOsgJJuDord39og73PIjel
EMRoPGN9KDpp45tEBh1QH0Ami7CnTL/keWVSnorxyz3P8zDP0Zm/YoceihyCOEBKqlIy5ywVrOnc
wEjCzcA6Tocb4xhUx1BYMP6Fu5HFMEe9PonFYIOAamg0Y4Nx5z24Fz8eaYnnRf01ZpJMpC1rJX8F
YJBpyQNV/njyjbstZAgdCwKthDEPp+6IioMw5hbWT92DRZJ1E8RjE4cmFXxomWpb6wqCJPL7nhvy
VAPPAH5IeO1Ebvff/+CcOSG226qN9+shh7uc+lyYAw+lL+SeWHnoIIVZfpQ3SbXebYYOn6HAOnRc
ZyVwhT62FWj9bbrbQnI25+3QFTzCTJeYchHO5BpPVhHUzu1BYYDTi7B2utsesm7UgDAkFTLnWFgj
2m933cKmEfbmE6WdDzJB6sou4uc8A0EGwkbYBu2uCIu/XuaEyBNtQ+k1/s4YF91BVXCqsITJqN1R
E6HaymReDBH9TH9NN/AgjhHu08+kRLeRjxwq/5m4nHmnsc1e8UP7RNB5NqSiNMageatgFO+wk3OU
oqy5jvKugmSJJ8JdG5kfwFvTHxcCKMZA2wDzs28qzyRkY2cRRNdPDEM2FZvRADknuw8rXATKVgxL
KDxVw8i6wxgs0JTYJLRoB0LPQdUjUYU29LQNhLPngaX+Z9P0NtNmq4q365x6pZ3ZeNw57musdDdy
e/SCiqsbt6sB6FLDu87GB98wRnLEbz0sOIUMCeJMBbkf7vHNDDCVzE6ew8Xi31oFwn3kDlnBvc3q
oMnD9GwmonLo/X+ONJKCuJgYNbioFPogoq8996KVg9at7QdRv+AS/IqXv/eqCedm5jPaUZHe7Rxg
m5KT+6UbhX4+XQSueHKeBq/RI+mEMEIlh4tkMpVmFNaPIJ69xygneG8ID09s6GfTsWpfpzx54qXK
rdILh0p7NMU46GcHurrZaQJk+x9KcONwn17NE5xhc3hCu9nopnyBm8UkORdEJLHDs2hVEyxOIW3L
czW8fmNE5RJeSmY1fiQNmCZQgO7NMgc9efV9A563lKLt7238HD48QlyugbgcLot2UBGZHLFlmv+O
SEMpI29+55iJYgbw7u+p/hYAJoIXX+e7gc+4PwcGiDe2FuNEuGXLsEMEDUZhFwfXU7Ll+gRCUhxI
lQOtDRpQrZSqbIFaY1Ez/HUMREbl2IDqN+R6RMj0RU54yzQKhaf9pSKelvJUu1AmLybOvOj7r1xB
qTFwkgUYyk3cx8JTzvLzPONfdnH93ZCQDD4Hngp/rtFQ0APD17Id0buMf/GZpl6hvD3yuaw+hdNj
9TU1VwaDQZtK3WEqw8U5Ke3z/XTdnYvjEXB6LHXRsoLU7U1buTDIm8XR+HAdG7Mw/rv/p3GLC9qG
sLpAJr19U9+vevf/7D5xfQEz8hvwdq9wp/a9uJY36yDKLhUuGAVX2szQ6iXM2QaukO9kUVqinnzy
CMxeB9G1bBxQtkwpukFUQi8KT+hYUZf19gllpePcq0t0VaOnjsQLkrKGqx1XuZoXIakQ8kR0IgCx
cw61ZK7T2wj9pbFstl8xt2Oo/AGJyZYigUeEIyqpdGLNq5gl6/MxOtSf6NZSxt6TDeKkTVZq8D+Y
/LN9c3qPn6S4p0r33wdKNAdTYqXfJ/VsCDKb+o7QSKw5HmaoSvaNwqTKNrCQl/jcqc7i39VdPsK3
3g99CAYwTWr+AA5XlkRyRNdNUwnwOBbtpAfMhQ7GQryw6tEBrou0I+3qrmbWoLWvsMxuMKHiNNsR
oLQB9EFOqvj+1aB1GQUI2a1z00oKPNOSfg5hCF04UclvcL+W8rRtl1EmU5/nAMAEoInX+7zIBWex
Oht7GDKT9atFWHPjBuk8LiqKnk8nhJ3H5+JGSe82qLO3XiMAot8PfBp+p3UxsXQD3JBpcZFq5Btj
34q5zhA2lTr5ILpgwMc34GdbAyApLH2J6X0VJfC4A4WCyH6yoaFJFkj2edPlvCKDrMrNtA06dPu/
J0DoPzGXanU7hydBzHv7KxXHWorNQ4ranyFhN8PmUW0xFXyAq3KhnyOMV3LGYqaOY45xwAsrSldQ
PLvC7y0LF+AmihdkZHIuJIDiwvokpivKp9mBPsqDFU7+KOBbdwUSPVj2ZTA57YCMfxQ9h1LL6V2f
/DlgWFe9uXUQMUkDwipgJuOxsykYvnuF44bWMlYwH9U+jUn15H8LBt7TKb1ugNEIVnbGq+EwkDE5
Fa+bGUOua4ivlm4MLEFFDgmVWcK8yrENeb2lsz0ySFqGH+YNehAjzw7pWtdm+nZSwHtMLg8pBher
5Diw10jJpZ4cTUJtFi1cQxTwtR9TM9zYfbdG4Q3WDo4Km5pfIHXlFR2lvwGcWOXZHG6TolaYRquF
qyCE3hMHv0ePu/Fn8Vya6Zft2dlJKyQddPKKkuM3BDptANHW7f4/mr8J6wLYPYrsFMrGvTSrq3ap
mxQIPOH+fzmr/mWn9o8/wY1b5YIhVUkXXWDShus1t8bPeD9/TkXdTkWVQb0mak4V2DejfWoLsb4Q
ZEjZElUBzVX6LN2z66DS9+0E4QNZX5nKfMONjYFSkwxJ8oqwV382CKPKeOrpBZukgnb7YgNbNyfx
e8UF0SfoNnSQKK/woVc78eW50PZEKxFNw4dzDLZOL+83Cn9UEX+OlrUKG1OqDM2OefZusVKkYuHO
mn1+kIXLV49acO3gJvhqtumE/QBAiYqjwrEVSnwPwntQCJCd1fVwo7K+AbY6nPrFBi3/haAYVXhr
n0arrD0eE2BqLqAgPso66DZ8opDzmUqTv/FmCkyVqdQo+nl6DNopCgPDmsGZTRqqwbBWAIr8afsS
WKi2rsvMHCjWVbbcbuvkztil0LpWwCMwx+rG1VPN0rqDajyXLjH9GCaQNBdx2nKdKrQ0sdOfstu2
Vr+ERnWrzbK3gKPx++SVmJ30sfu9xbxvvT68kfD7YAXvKLn+5aqUJxSXMA9vZp1N9X0ui1OSXlYw
8h7uune4cXLPCjMvwXl+8/nrJGzQ6jF0M9GQ5M4M8+ZOMKTAObJ/313/fmW3vlHR9jUEZtzAQgHN
hB3zAg3qsltCcM0l6ntiMqSZVBZqhWju0UJc+/5gqYi0yTHsd9nTPDx78/sE/PZkWhQGpmsO02J4
T0aFzK6zZHXhaBm9llgqERBa5CsGzAXEtw4JF6/l2ifKHHVl0LSR8SagUFxXJhZ3GnPIXf02gs40
Gkyv4G6seOedPxB5yx59i9KBYaTtWkwzC7cSY106DxsUOKdWlWuM31TGFpyDFYIxhPOQcriHsSnS
6dFbPbIUumJP1iUPQrb42LeNNDcf5798cV4xGc+/wpnj+EJHUfo8bYzgz1i6s5vkNTezpx60ebs8
clj8yJjLyDAt/124q5iKKG62kXR/zQ7NCHRy9K+x+EdxDhxAu3k2xiljV3ROKayg4gqvFCXMaT6g
D4tbeU0DKL9S2k5BMU3CqCLjkTitqChqBYhqiIOaCaiqIjMSCfS6KlIbRsgpQZbCPYroQEia78KZ
yxJECBPLVrS70uSQhm/ROSANBEba1XNrB6IxoHHg9K3j8bDGa4ONDSWdY+K+gLGelYktfJ0y6ac5
8JQ43B29gMQDAUVpYDuWKRzlKtnxWYvezoKnK8Kb5kZV8oPCawcmlUGCnzXOeq1N++cyFQFsUiKR
gEsqBmMKLeCmHUfO5OMWynDK7yM/ied/8/5UADoL3uTEY4XQ8CQRpZPb+kPTPPRmGLvurcbrL+rg
UJAaKVPonA+Z3k0lXaDefyHRJcQ3X0XGGY999ZdeLhlw379jAUXcRhsrbePMHR1TSgMY0L+GrUaJ
VHY5xexi949oLTvt0V8MhwryiBvlel47owVeUF1BryD4Wy0hxMP6YVkhJAA3K+wtnT3J63+7D9YE
IWcp6SVMJquKPtPZwPRkxFCeYmgvnO+z8QJU3tWSBrazEzrNiADPsw0rzL997Ss5XH6zgBdbOU4n
+V+Jd7HNdPl5kw26GBeOjbORf+D8+8PmTunDyD66HRy/DYKjdc0KnSC6xKrL6bVdbgGL0ANdJ5mc
TxU7pf5Sw/BgPWGyB65LT+3Qda8RV4zugxq+RFXy0EtHIuygBC5YBdKMz8ChA8N90Tal6JFNs6iO
WkaEcCn3OQ88PWIjPZSWuheRP7u6j3LlKMesJSzccBmcLM5YcI+fbuRkimqB+6m3TsoEOxkK0PQW
0sel3R0gbdxFyYO6aUWnfTdR19lB8JMqAquGYKK5XXdb2aCtGSonbgwN30V9x9QGA836hS8R9VBt
SAvzA85B3/qRWTOSuCHb+SVzVSpUVePf6PDjtReBiLjO1O4Wfqi3zH8VBtFPAYzqOehc0L+rZc5W
ReDKcxQv7nWGHszrPxsU7/fxjCJY2oMKsxLNFkZZwjUWX/t0K98fuVOZbVN/lj7g9WzHF1r5zDg8
Nz17OO2Fuo2CmvWoZjFdQ+kModTaa844RQHWJLYt/RzLXAZ2LFkDFhvbx+4sYKldOOkzA8LIQkIc
zWLbyzQsKhiuD4gfveuuoGxK8sPmdXd+OBjGWJz/GPiPc/5mD2U/kjltwr0p5fUyijh0EAxVWiQS
nOZouLqWRwIpJIknXVQkCCyJ0gyX7muuNbE+ovXkMkRO58QeDppaePTGXLdWAI6JSlQvuAPZxPcy
u5o57NUhXahk+w6O+2rEObK6mLTpZulqe+A1Ubz5jmdfiI9M0n/RlgaIzqeU/lI/cyBDoXaMGgzV
5PrSgxAqhC3Klg/5svRuo7PbjDpLp6Z7eJ2RAnQHmyOauwpnsI+mtjvXDkCjcPwVnncuQKE7vxrt
Hq7vkE/MeoPhU1nkxJmrlIaSFIATUmmkoPNpSNvfA6g2OOTrTvvDhxa2/y9awT7i5Yu0KFCW1L0K
X8E1nrWn2Yz6dpVmgJAfph/vKQ0lVLYcxJBR6gY9rSsM9GC73xR0aChKrd44HBBoOEhs18dEwb3t
GvupJlQO+35cH7KWxks7EuT6x7TR5HxXj2Md4LiHixyBB3mN/YHxp1SiqYR9COKYASsqNAQ2H7mH
4tn/eS1hGfS6jZ4dtQHZ+UNRH65rWi/8vMcWKvaiaJhOkabQ2CCJSfSv3IPnDMB/2976JOtlw3KJ
lVv9ASub46C7YJldr6PC8F6QJu4tvG+d4UJzAypYMYrq9y8FVban9yCJcRFhU29X9vfU7rHBCcgT
lTNy3lU8EqlwhdO1uIx/RuTQ5R3U5lKO3lLW+QHsdQHRRwdR046FlJ/Y0nqW087LYNxcPBG/xLAY
O8VgIb0y6whokZwu4Ef8eBPsU+8Zmwse1YFw4tXn9z06oEcYY2tXKetdm97nd0jjNg3q2eC6BBFu
TAKbZ4NaJPxQnY5AnQ1DQ+yAGCDVn+Qk/ga+nIoK6oj5ZmsBRxZU8iXx1ExJ2zc+9BXU/xIbRQ+f
Y32jU5iocB6pQwtwn2vYF91XQWsjYQ1zvP5fTiaSBkojGIUsAOUdOFPtFRIAnZRC2UL42/ISiqdk
xgvRS1uk71gpmFrzQIqmAypHtYQOSWPfzN+67825wAqcJx/oUAQBl8GOptwHKLLCCR9mXFWDg+kO
Kl5ro3Y2bUfhHNTkQPS5EzEogq29DSwgiwJxrBKCJUsvVwFPtOpRzyW4bzo7m6d6Zefb28eeEd9f
s/XWqls7MK2mvAtZZF7pmhYe0MI2gsSRz20yJsn4OZO/R3wXW7qMyg/qDkvOTv78JdOMr0M9Vvnl
06jSv7tET7WynaBVmIOtMlUUaOqJeAc80Aqpirial4Cqrv31HwZ2BZ1RikJhy7OWJeX3QHIHX31u
/cx3+9Ai0SO7tqrxNjsO+LMEAYuq2OUt0UvGnWIM1qFeQCqyV7ZlNb5wTfD+VowkFdzCepJHXbWe
rh42FX3n6a8uJrgQ7yOgDvtjlED5BGMNmvK1NSlyuPfTE0txxam9hdosqOnYcygObBoaz5Xnim2N
I98TsuLcU1nyr7jfMIkDu4UFY//pv6Qoe3edUkEmQTM7suC+/XyMZd0Rjv2wQpGO84Lvv4ONVCXr
G9pd9+4W5fV/NNv0Ftw0CvFBHHLf4lmlUMr+rxCk0m/kFVq46tz2cDNt51it0vP9vMaroDJoLGiu
f9goAHzpjozX4ZCW6GwZuykvlCQ5/YT1s3S9Q8V4YakAzofPYK7g6fXwaopV+2sPu31pdshAaQT2
oxQhvBVb5p2fsnJGQY6HLIq7iXvVzlmzcUqG95hCDdpj+hCslXoQxIYv7Cdo/JQ2mjm3l0pw6dOT
W1kWL/5e6a4RBeJAJcbRqtl6UBBX6cycrkREBOJUQS9QHwWNyvRqhID2k3KuIkA0cr60/Lmqqfs5
UGTHBchf++Xbdg5kVbjvcGttJjHoXzL5GOwA83BcmtqIAT11yismOEK/FKkgEONymwSSl9KELNzf
NFxjEMrnSTnaOUGnHuPyX8yO90iDILNRO9iAQZd4gWUOQ2s9P7P34sIjnZ9UBkh/VsE5FV+mKWgk
Qii8B+6QzL7/tb5EMfmX0BbUdSGmCw7/L9CrVYK/iNqm9C0UbJh4R0S9NwrPc3MF3D6S82Dd0khd
+a5naQWlRoPMpxTpqeA4V5MZ+qrOsYsx7cwJJO1HLGUbC8ut19wioDTqRO2hyJPknDBSqMXdjTKe
X5QTWtYU3AojF9olx9JfUoIf9iDPjff301F9g4CDd3kvP9JlJszM79c8ZfytfieMrfJOyeDnki9+
mDAGpEkvaz5tP+Rb5XLZJ9tfVlmlq/+0xOdTazzJVZ8FY4Lz/y16OKX6wH1Ip2tafp0B92J1i9cC
xbE/8bHT0Q3kRP5XIj23loXsv5QhyFfMrL/MdtcI7515vaRdVQbYDpRdPoc783p4426TCfvHk720
r3957pGbQrPJTjTDZwz+MXNFZ2iYU884Kw3wYKlxSZE6khA3FmJ7usHI+33ki7lQLnTVBzatKNkW
9haN2vO8qHybiI0Qwy2y6tVohkYzhBqhotXhEm3KrYCFJkprCgB/+SvV3wKhYtrKHkbL5VNknphJ
y9Mx0wL3nnOUuYO5kV+XlBfvsr37Ecjn+od68OzQ1kx5CDkju4HKOIM124qTNdcdALAwvQgrpQxt
8pTf/5Yr+dnuEde3EiL4wXjLPfPhngkvgBO3k2yvKN1mGTvtUgiY6TiN5KPLOjdQu02il4AyD7s4
Z0gHfjTaIegjkaeBedMlQPY20Q2QU7A9JzmmOg5J8W10VK9Q19iDqym241j3nuW6+ZttqjLCoDQ/
2kP99w/pFYpNQnSvnJslet2YrCXdf1M2bdyuNu0z+q0py6uBQKbZUpkSQXHQhIFWAWX0bbtDzWw/
ztFsqPD1aP7kAaBGa+tcMJ1j+JeXK8BtFR4kVFZxaESYaSTIz+pLKrYRbtbiGP11wC5vpDEh7fF2
wVN3TKgjRsQ6injHjwm+d+jaFCB7DZr9G0yzdsS4p48bk4Cn/Z0LFnfE7iUsKUXcua3JkJpisLUM
zA9IkTaSIjiNfMF6Cc5sE6mRBfWK5vnCCuvaAlP6LyF3f9teMPK6BIZ6SEU4J8hUtu+PCxJdSISW
PxYiQfpIbkd6tmaN67HFCsxZrdUYbef73GYmJdTeYAGvHwaD1mVayKSDGHYQ9NN9oL56nixnP+M0
qUqp+Qs5wqgc36YGaLdCZb58b6pnS0v5V3NO18cv7g2URJCwEWsBnO7o/F3rQHj2FFb60TGAEqix
c8fs1r3+g3YUWQz5jvL5ce0AB9p8OK2FiK2h4DYgONV6SS3R3hFvHXcbOgH3SSnK03guEEFteA/R
XwUqUmvCIfx1ESm9a+kU4bU7BFGFwudF6bB2n7dK7cgtrDHHT2E/C4ci/tFt5yD8MCmvGU9RyGk3
pbCttL95TTpnm4n5NEQgWKvDJ47z/aiAM8W5GGtqp/EB3pvPymEswqEdsFxHJlcy9KhuONG7lUcV
jNKja/8EjULUwbTmZyc+cEd2psSAKPxwrI7h6FtcgFa5xKSAjrPgKrVLPFWoyQGSI7WE31h91bEf
5TvyFE7NcmA9L+pd+H89oVFdv3dzzK3pEzxRXOrLhGmsSoEwefNCZbdpqERq8ZcZbpA0EmnCdkiK
Sv1mq5cKCL3IYLpeWKbyiCVWnPbZr7TQKi+1fDigmMxpbv9UYIkGt4XrfGbhH1ZZskfaZzidlu8K
fT7WXCZipXO/RvNOrt5TkXZrrmd6buBSTSYKLwKmPkI5c15oODl2C6OwHRI/fhyws8K0n5SSfeEe
aHyOXF2OG7xr8NdJkuTKnevzhoghMcbL9U9iZfT4dljYaQZlXtIYZtCp+/Bf8OOwzrsEnD7qtT1v
HapGW5xxEwRVfln87e2nY5S7hkWqFABUcfgqVqSLGXIRG6Yxx6ySUp5cZWXboBlYHyGxu+2dkZgk
itemii2AqiHuOoj0G3rPTFf+nHf8mteQ8Eazs2XR0qxF/X9l072MRymjrI7ciKYG0IkptY/78cra
ijpoe4gkRPMQuzNLQXCjDlLiYeJyaYeC2Lcm5SJ44F+Mkk76/nu3QcCikbmxxRZFP664hpbu48tZ
QlwavnABt5jqO+BKFJfy4KKfdpfAQlLz8EO6/ueeCx0JCvREF0mklvC+whIyiFl67H69cXAiygEv
zyLkwQaXTSrYy5AA+Y5bxqquxUGKs/9BwwGDPq1Idmk9ohOEVHzGIcTS1OZa21P0FCroXGF6s8V7
eEv03ZHeinb1NkhpjyASe7ZKsNSAoBFJECqphwGxbVKVYpK3K063hRuCJuQ90WAVCMhqZv/d3Aa5
gNervlzREFUjH4z7VvOCH/rMzMqH5fthK+eNwzsS5mOaHi9WSxF+YDgYQYqX1/VHg3Nwoj4j9fRt
h2tXa3Ibmn4tUiBHqp4AkzBLH9Ya5IuSQcHF4QNpsN2sWmn8OAoVaEL5OkYCmZQdZwfNXf+Nz/6R
BYheK1A5E7U477uZOPHI0bvUbuOeuf9mxGrhf6/3tsrHoyJsr1aZuzVmCWbk0cQpCNNIsN76mQn3
RA58OFdL0nJ/vXnVtBAzWFZTRR40uQzZZrut8rFh37HqwTcPAtctqytkdqFUX2KJJf8SkTRx1ZXU
O3MxkrQmFQuBRaVtZOqQ1uU34CC6cR2aYLPDhhjrfKV0RhF+i5E5D7LzGH8zJff3hHtWaIHZob2R
DUgLytHRjuMNHIxGU7Rw1urQEevN/cZKAhGWeg3BL7vBdO7+9Ce/QfuOBC3yBRnt6S14NtaQJ5Hh
+oidzfSaPC3suNZL9HdlNMQwQBAsuY1DahvrWHZTGGmTUmHNex9GJE26yi/plchtdTz6VtGr217Z
t6Sxm1755UZ4sGE9Tu9KGUhBrhBienrs9EEWxkKCB8jeQ7qQ3YH0Y62Thg/0IzjNptLDgoYQqqpf
zqJGoAQfXGegiyb6pqmUKPoMuKUo1nY/VuyAP2JkktgcvpLxH4T3+159Glcp62AKjLaZ3szAlSy9
gN39vgjsRZumxzPEu1CK544fjbKqYIGM7QKMAQeMR7ZsdlmcbuYOEQb+uvrJkl0t0hWMLa6rWJ5+
rV3NlXjaJ1kyXnu9y3MIzTRwKCd2NdPH3ZEB9VXSRRsnBYUH56oC68xag/2Uv/NBok3wneFPQErh
2Pzu5YcCuJzofVGAZHNezM+tl0eB/PZmHt5hhNAY7aBNEaA6aIrC0NfMemKUPhmTpX6SuyXPEVhO
HO1KKoau/lZcWhs+Ma3hnGnpRL+8fr/EP4sRV1rKMoqlBVX5hQmULW3/6Df/EhreRmMiRxdhbvbJ
FVh1J9Rk5g/vAr1pOZPxo+1fNSaphYTtjjqmoPaizxpKZD/CQGj+aNpe+bsU9JBq2EA6m2aT2NMq
qj3esagWb+mbAcZFj2/iCJWwPmtzTDF+Ku2vb57/kvlRGdEHnGlcTjtfm5ERpyP7KqiGN/43fp73
mSi6uCHg6SAsr1Xcp6Yi/ICntsdN5hpTQRFF0I8s0jz3Zf6qB6ngCYhRBtdqkAyg61APjK6VcAtP
3NAvOSlK+eX+iCrRyOJmvsIyw8TPzEU+MXfZ91FZ4wdTrA/fG76ToYG3gX5zB2J3t0KpRsC4OEuj
HzMDSaoIdh11VYZU3LN2F0NgVz0lD78MmOgPMYNYIKytycxrdZZU3TEOlwjG4chD8cdGWp0NwrI1
moTgAb7PVwe6uL/VuzfUzEGk9I69ScRQ72VonccdTGdRAtwAeFnDN/BQRIiXYqtkRulyBWqxd+Ts
/dV+jF9PSH9x+XqQIbkV3qOkcnyvaQu3ZQfZ7hiClV6wIaU/Re8Tj5qo3twlJffYcvu6nB2CQZcb
oINw8lT6BWiXz88frU6UJfryeVZkSEwfKO4hKg39rY+Mplg/TTUhni945KJ+r1FNw/O59vl6rSBw
vUb5bWQFlDh+KK/Jwf4Va8OFvW6Zfe+Y6AQTr2kWchS6vZGwuBxKSBH+LEezaKLohyzeccyIuSBX
fMUWXKLMn73Dy9XDGLQ5GmF0Bp2S4Ye5IVMTuvWaD5xdtY0r2j6Bb0r+t/PKrD3w1Ti+MWkI8h5W
L+7SzY07dTBWKvyPyiRkiTEmBWVRIQoo7rSmI0URUcEklokg9IvEMmlKJprFhqUI3fZPYnVOHhXp
tvDHnRnzfCkEf13pDcCmYUGbrANLi6EpQP24Lna0AXdZyvK8svyIfSEFp5LaixtXiSRY6bBR9REG
0AXwNL+9I++92cLyzkdS+5A0GzVgzK4ktJg9wuMwc0w+ALQY+/TdhsFhH3ghXhVmWhKGZ1LzBLmI
SnA+5sXIB+Obns0y7Hq8Ri2VxELG8jtuFoQpWN6HrZyMQY6i0A9cmZjFtaLDZRMAJSbgR16xrus5
8h1h56VZlCz8jyjS9R/r4JZZYtRTMigIqGN0mv3r2gZuExh8Y5V6GJs+QcdpTHfLZA34yIsShfxV
MNsr560kh1OwpA/65Tp7bb6Ebn5AUe/ApotlYHsG0FIlFFW4LSAcuANq37zqD5awoBeGCb5nbsYp
boWdc67fJmeqKbsxNIMc9UDBVJ8nQs2F1E9kN9UX2fIbzTsLxA8q39s6iZwzYZl6D63jlL3aScDh
0e2vKBN7pHGLXQb3na7jvKX4uEAWbRvjl5ex2vGm3iYqLbMD+T4C81ew4h2Le/U09Q46wtTZmZ11
DvSXAD9Ff315Xu3Hp1AAVYSrF+bahZ75qCEhv5JOILeVQFLvfa2FB6faZLJK2aoJ4nO2TcgYkOtW
QRvWXmzY2cN9Qv08NWzUgq93uAEDMqecvMYnEOzFn2oSfG/BVkDsjwkUanl2fEHoR49LA84rIk4k
tX/mzfnCgTBo2cno99GoYve0GIX91To8KAU7qWfl6HPQ9Vt4BXjsMB1crx1we0quCD1oquUJmNej
Aues6W4riCH9q9oZLJIvulN1nKSPpi1LPUSCHQEL3itL8xfvzsE1y5hQx6+k4j/+/pG5G7bsdQDV
4d32U9rlSu7Qejf65gKcKvb5gN2IKv3u6WOoc1FkXGUrow6C6uFzOzHeSFZAGRYb2DfperwNqZHP
cTvyU201Y5jU2WrKnFVladkcgwKrwBFo+yzmNhOzVTslZqPNT4wrOZ+Ki/dvT8UgeDIwy8NK3pUv
ZR/X9rFhqyBbg0hdRNAqopaMgp1k3dBv6jJfuImsg71bBvT5kobbvc7/ndJykk76QolhLKzj7wuW
JEEHHskjHoggOpF9oJQ3sqsEaanP8U16qpbeU+A5DKki+iu2xFX7pEHWwX3gVFqq5I5yc8h77fHv
cwsgqk3xavFqDlyIVOso/sWnRYgOs0PjGKVos8ESjBn81sPhi2qEPvVjkvUOJsyGZeu6TkDREwrb
BBrDmRV8EliONMJMS1TaCGSMeaPyux5Oh87yyxx2GWd+upkO+l/zL4kpIsFvpFHu3fK/S1Wn0e6O
imENZJw1835Vojo/FmSVEHsKHUInWWl6padgyiSBLo6e2Ad/dEEHwVuUTSXept5rq0k56sqAAgBs
lh0gFucMB6nQ0SrhaL6XNlAXrvvpIiwyglQcBvq7RMrRPal17XHp3rj1DDNq9p1R+4yBokJvRJzm
MDfz0MX629T/UV/WWokT5EI0axUZRPh69KpTslwY91/fiekDmWkDQabyj5lpN7n6zlvwUF7CefFd
G0YTbLg7CZX36JCKMiVB7M+y3rWU1kPwagrHka/quVVtBNU48rFrji5T4Z9DnoMkGHMI92WckL2J
dHvzD2s0/58Xns/Lw8PJQ775JSMluSFtHFqAaIicJmqixr06uFK8p6CLc+Cn2Yfua930P6j+OaMV
uZd0uuMpdfwHX/3hCNVRuNimAjdXx1SKn559opGtGpKg9hMEciIHbzldmhF3Nr908sAoXw1wVW6b
FDI04KKVqoC/jZQUsmPyy9eNiPuoOWXyqgwcoQOvFbdujaBLnj9r6rHh0++lgFqUlbhuSm/oA/UB
uX/XqD6AFakgKV2mFR16DQxigd96ISW70yPAkE90I2u+EXbaHCC9MZ0c2LpI+tylaja/XUpUZjIp
8QjDJRnXzVBsnfFNWfczcyI9hQNijpD6nWflql7njsYx8txuCBLrNU6xm0rj3IBiOSC+nLOCJc8q
z9p/tNOY4fhJgST6mOxd0MNdMh9GxdNX3kVrv74Za8cHvOveLLNPipciuYqmJnbsUZ4AIbrViw2B
rg2p7YYmVXsOEFPBTC8w3LbWeOKXTL0uOf7SH+GQRqbhgAYu2Hrtpj0+qYRHIVf3MMy3wj97Il/N
eRgTkxvKdNQnl8KcN7z0EyipqUJfiE1HPVM0cHHRYlnCMrs8ldCvIwir9uaW/ob4YcMVfinNbOds
CETZTmR9jGkrmblvbELEWr17PTJYWpzhCr2NrkE/g5vTvHdf2+M9BugC0CbMWL3ZPvOBFOFtMOPA
vMnrKQ0aXXtu/abOhXR6n8wF+m0qvyfER8v6HA+zC8EuFTguSxj3Yks3UisIvJBtNql0adPPJOh8
g1qZan7pz/mJmQU8CHg/A411vaPxyuZtLQiL1fJBFcS8Xs95S3PZuw5IDXBzieNpiih2rP18UJdo
J7X+20PA/76LEqmzaTtSnBFwsQncDVRb2/IAdbYPjsVRs0E3fyBtvS5nkAJMx6mDmhjQiJx6zy7M
CPyrOLsDGwGC8I7zLAiCQQmh+kN2CwEBGHzlKChTKp2GyMpphaWEx1Kbjavgh3637uBdSsKJB/nE
evAL/8Yg9tihO0Tq4S83Zhfi7iYG/tniqANS291FtxfTpsA1KMdYkoty+gdyjYXwNvK2i5slgFTi
5+WKwDptGROuEVajhFiL8csMcmcBY2hgD0jwEoADNQMi1WELTBmZTjuivSKLSCv0OSxyCroFfm16
NldY1mvsqNBv1lXp8zHxXEQjFeGkSpXlcYTB+v3A5CQ4XM7AX9JgTxoG16EKnbl3udjW2yLs9ud9
eUug/VWhCo1XAGkbLGU5lgaJvG2ocjxHoA/K5N8U1w8cznn016C/PJK3Sl7ThGWVIfpJ5fociyDu
+JJ73gn340Vjr+4cueLC9x5meS8UUKTygk0BkeF4BZFTtF7GRuGH0pVKuQD9lwXcxB75kIdWYk1y
zmtPiTuRxml8s91UI3MAZ9rVSEBnYzcBgVd3b1zizGhhnrkkEZeqktlYkW7xaXe2u/PGgaRzIL+L
X/HccWo0b2lsV++yDvW38eTUHFC5JqBiLWvg4YuiCc0OUo+XItZMLIYHHogPsWefQJp4ETU65XxX
sJgjpGk39aWSbaldUVGwJ3hVztqo1uHMN7MOWvgCYvIUW/K/XQuOsEg//EKID9k1YxLVAma6tbWc
AYlPabxK9OuDlLsyZ/FdUewZjbuqshO2HstT7vM7H6Bnai/P9D30lQxU3euvJ3OJRq5BfihKnCwV
W2vMNXEzX9UaSZO5lVQ90koPi0tDScKhCZ4eqj8xojgA3v/fzfNfGGppwfcumOGl4WxNSVTedkoB
b/A8GH73gWS5mQE8Oqu03229IVSFtB1hGubHGzQefwVghsS79dVbF1jvUvzLFYIP59dVM2PlVAdc
N5nlSZS6iAF2wTuWt6WI4JUnO4sYFyDwvU0rWILMWFB+phrFf1UC+ZAkypsTVG/y4M+JBMDeDlnO
1MCH1DuXweBUEVQUji6muyWbLbDyTOTYHcg8VocKsHlycXn72BZ7mtGT0OfBBy7hCB0/zQ2JGbpE
JhLUWZFZqVgecge4YRpmrm9uw0LaiXi0W8fOzRJmuEs2rueijV3/8TDhxunAWTMAaedvFopjBfFx
chF/vCHasINm+RtEdI16p6Dgw3lodpj5An/fLiSPhk6w+KFyWDjjFozz++trMZRUz6YTln2Mh/B+
Eo64O9SPN5IK6eY7xM9jBlFMIA3Qeb0DRdScRyS8MYHcVFGEm0id84c5Jb69gPf/0/6t0EQkW3tl
7RvjSdjShGgSZoaMUNJfp0y2He9zOKGmngRSXg0L87rkQ9DMx+B6TaVcp/E1lm+KrotUc9fhtc7B
v3MJcVnAJjCP11K88w7i3qIOZUYHjohcxSc0xKjIawzYzCD4nOiIhY9jue+uoRgn/qtU2BKuIqdC
N+8IxxafSy2AUeyJZtGpWQjuTGpuw+XeFUt3MvT0AmtxAMH7ZkXgGfvk/B+fdB1C+gg+frBwGlx+
iSfvA5fD+/C4i9DSB9PfOmVkB288DlSQ5Chmos83EE9wOoFxwvVBLTlGeHTWEVvbjaEcXYZYTgEx
ajm32H6zujYzpsqQqCiVGbjw3e43lvDbH3IPBi0w0yLkPSRRmiZ8ORDR/8TCAoa5eENgzcYVaNok
WSritHphZ+2FcCymVg3Rbzh9eGh9ixRVhnt7wRifDUBrmQaqJFrhpyH/4zxpJx9OTsjezKI4i4x8
ncn8CYBMuJdPfX6i+9vgjLXWuEoMMWIoi+wWYzXk/1BZSmbJnYvxM/SivNFBAYDRtFY1pVljQGAo
sOA1qytba8v/W9QRcS6Xfh2EftvcBymg8CRMQKB3lOztr1UhNHG+1LKYf8qRtH6v6dLfmq1jMafi
eMiNf00In6rrZFqFh6ALFdXkxmSCrsyvvr95OcHsCy4CTUVL1XP2JvgLfKdirZShUsvSROLCHQIj
oydhilkR+6PrqyTxqYeITyTrmPaxHV1CbQ1ZyqsUqyRlC5Wbo86m25BJQL1UT+6F8S5RgBSStWFV
hPtsM+kpoxYG7pDDGeydr4rkTOssFUZBbV1h57AOqy0JrIr3EaDF/Zl67yatfr8w5rJP9xoYWN/9
8wofQ0X31gTg6lJ8/HmNqOOHr0Jv3JSGG2xE44nPRkp6+ts+nRwssK/wtApZv8izwmxgGk3ffPbl
MNs1z3OuDI9qfkLmHqwH27NSdlMb+lc0OC+udA4IW/+34fDIGDoIl4PtR+jHYVnvjZvHQenONle5
tXrv2Uk9IBb6DcVGEWN0SWfwqO4rvXKLmVgYJeJ0+kyB667E/5cCrqFk6/RU7HIaaKSUXVekshio
HcO1t5Z9Lj/jc4mc3YR5zaAsR0h5lq98/QXEHwLtli7rLyACaR9oTk6udylxD4b+UtetmG4f0kht
1WX5j2UIdw2pm62aMjNH2iuWrz2qG2mJzYY+2cwMVGuaOHpOGfbcVycORyilX7fVYnmrI+xaFcH9
CxwVM3bK9gwT//yEe7+pbuKtL3WnkpMBbppSEByT0Zu5nP7pJ2ToM3Do33suOIOLGc+knGagv8D6
7WKRt0nk2VKNJEg4VgjnsuNxNdws9c9aSyEN1BDqyD/J2J0k5UiQm1zjQ9qg+IVGwnEo2Qa6zosO
PHO+/6sb7nodU7E0ABip+Q0S8AYhetezVBjYpED5NT7t7reR6c+PFsiIF3Xg187nVPO0kFsRqO0e
4SGDrZho2PI9qz7nVSqjFIOOYhotK1uXqQOi0xVNsrZQOYaqQr/KJ0FIYMNXptTc03xLC2Dv3X2h
uBumEhZMXFMEXmNVLBv7QVSo3ILU8eR31/vW0Pg/5Fp2HtA7qwOt87tOcZ003ApKNUUo/wQB1b07
9eHDNn2nVvRXj6N+MzyLb5iN0VecYaa4HFvBWmZtGHRmQlR2876SRgv8tZD2CNMpqzcLbu21bXsE
xUZBgEg4ND/gLskuxS6AUhSYQdBQWz2xa9us1mm6BVYr3CKLpzpickYeAgOs5E0ozJKbeediXbaq
n/1HUUG5cuGlgLIiwETI2R2gzEZKIBuUrC+ka9k5nYnIupI9JDgtb7ZdXTe0FltfjGV4daMNnfKX
SdZsrrRjeGeld7VsEV9fuuECasaGLFDva/chv8r5yJ6WuG6dz2JFcSczYqht37mDgV1C+ahpoaIy
o8myck0odk5/jR5SAlTSAdhb7RlciNxW8hlC5yWDvpdwGd0EEoFa0wa8vADA3Be7jmcOrBDJgCW1
Eq4tboMlS8Qc9NMUVClotOhT4ntFlsotFrks2QtfLiUJAA8nvecc3wFi7JYm3hjbxheHCFaQD+ss
xh/Xh3JiqX63IDMQP3WXPtPC8OeKzKtW64oebEzL+TTzxs6iH/xCnR3HRvaW6EGW7qWuY0jO/ODZ
5Z6Zap4jBLAXwQ0oeInFjFcgNtbDJGeGF84bJCvDfNQGxhpD/fjAEMvOz/mqIZYcE4BgOOWOPUgB
U0xXRwv4b2SogctrLMc2t7Yqvs6lJtc5abepcC+lLmImOOXpNBtagaBTIfi2S7R5378r2AKadFmd
gkcgohyId9KU2tDfdZM5/PEkExefM5cHZbpJ3mlkrLrZHIChrkFraXCmt47BpbPiFQUGTkuCZGDi
p5TKI7UauDUIvTWd59UvmySDp/RY/YLU24g2RyAJrhreP4NskvZ9BfcS+vur0JPoLqRbhECAmcLc
A28OjvnTtfBs7jSHm+RYFKjkmEZXpbGFIKFrAAZgLJWnEQXRYcrCJX3vFZ8xaMJOmGcwYykumieU
Q7+XgAKQ5/8mx1CPaQ7K7mWdBUI307/hG7uT1ug6TituHGT6HkVPpBotYFubX5qog3e1mqJuLwPA
3QEvetNp1u2pHypCg6vuj+ynbEL49D57Qe6yX7UxZhjFsUxjEH1ZIm26IvgZWnjwTrrXsqwbLEiM
gNnLw1N0Z18Zs6xh82hGk4U0NkHsrRR8HC/DLgLzg7+ZdWfACEDjqSk66ml86IsBt902F27IC/ju
iAGo1OT6/hP8Um43prTa/ZchxknA/8bMHtW9TYw2WjIC9+jZcj7pJeyMB+dKO4GzvW4G4EvrwT9R
lMnj7b3CbX/2XgfWilPA1y2XhER45nnjl+BMn5m3qf0nBP0bj5f27396XxpRHdX4d0cP/4njHQxM
Boahi3dwcyP5xvYFpm6PUGeyF3vwY3k1Kd7HjJdD38dzpBsK/i/59kaf/hajHYwkYI3445ULMH5Y
8a2X8aQzIxPPdsSblSTCXRpkCpauGUBnjrJvY/XANxyRX8GW85XACGNWuKMx4KFNe2q7PU6+OUAw
Rs9e7DjNHq9TPogmqHVT/E4TShPSex4nJnWjauE682J4e0g09f+v9rFy4FrnkMeltezTaAxvYn3Y
ILCIS/tBuTYYQ01AXDXb54C/oFS6g/1lQHDUfhw6jzA4V00aD/9qmwihoebQILvYFsJhWl5z44g/
s8Mr/bkshkgViEf5Zc8xM3QbVDmNT/vEUkH9fyULlxKmArQaoQ3jW7SdpXJmbbn/xLTMh635RXtH
fWsBzEp3hGhoBAmmDHjakspzzFvY0XcaKUH3oLFLyxNRj1gV3PiZN9BlcsSAfyyqxAsDFrsbGsSB
oVKZjRYqLNytsi7VLzN39Vt8/1N/02YGb7oSS43L+usEVcybSvCjzCDWNJ6wdLu8aO8JfaIKpy5x
mE/1pL1LcpsHj+sKCVMIKfXZC108FxOLArGw5KdZXkW1dygMsxcY45IB24WRqKFdysr9cvrNWb7B
FslWbZBtMB66/JDk/9b0+TftzSyAlAIbGgfRugULhZBu+vcxi80w6laI42Ghn+ebOSPEYA19Cv18
fIyWrTmzBWZLef+zaOhrb4wyUT9STyw4NN+m+WUbGGOYmE9ZsamxzhYQ/JpIgCw6xNdNGjcXiVC/
SmkgE49Te1xvWQ6/D4qcW7rKoV7OGrHLrnWvH8JBCgijHylpka6KHZtYC0Tg/6CD8v6unZiqpwsE
Gk8xH90/GeGjRKtbXN4IrsAJp6bCAkkUjuVp9SrQ5Dv5VQzQFmt5U6E3UKkWAUXzmaeAVlQI97R3
Ae24gHHFZgIJPxh4gobJBVVL5KWjyQlUbeq1LdsVHfLwjAc/V+CW0+aa9HRsIDU4lk7UxcN8nR/l
hdUez7Xsm1yO+u+rjdW0wmQWyn2oqekIemOhqz7vwancXkGPH44fIEcbX41NtIuUPvzBQ/Tu8o+s
Jwq/nHYN0WNIqICoMCPicN7sE8LD54u/CZinL6GACiXhnKN7FeY0FXza8De391ba6AIf3Wtl6LVh
s6j3dj7N+8/M3ZALAKrdmT3qJH1tkp5nE8Yzx9an1JYoIT1FN6TLujD3eayN5SHXV/ebXvyLCAUv
I0HJLo1W6jDrztEMTCNRv8SoiMgk+IPRR5YNzVFxFWGIjmUDwqHfIp3fVcCArk2uEowdpZLkN+ou
of8qEANTBlNWPovG+wvDYB3ceIwEBTO6TdZRgSbiIB7MJ7hIHS37uu3iUDIivKDrDlj+7ycdIJNx
k+Xk9DMIEABpX18H+gUecD30GARxcCELI2eZTTNSpiayW7Ucn2CFt+NEK7fPV0bQu1SCXMpcySkU
hvbP+Mafsj4cu837XQgdqt/yNQ0qX+WUF/bbIpgtf2xH+jh8kwoNiazYoKfktL44rbSafS0X8mC3
AjPhub/RAI5gTAZN1KuZgzZv+bVMG90LBvyzSeuu57LmoD+cLXXVOKkfO7HaVreiFuPuysgik8x6
K/S7YBlsQ4R9138r8ruYakgSCb6YBPSorYloCCXmnQfHvEAbm/LZvnXQ1lYOVT+yLFW08qbaSKB3
FXVwSlmJXQKeCS2vWWdpWsPAJE+Vl3QiRDKIx8tf8g2qeWBim9E8Mz7ivqQRtLrOYdLlQhZH4LbR
fIr0vrXh2LQWb7EvVa4C+p8yLxjFeltZlf3JasidtXAKJmlCTsclNMkwbvZ2Fo2hMGvKJHQUiUnp
H4xrpqbdairXFTJIQPqYJKlJSeclNRgRKWlgX/dyH+5O4+wzYj2U/wTNiN0gQ4H23/MnPsyYNGCL
qTSGgnV0G5vmad6BCgh+ZeXhi8BDM3ZUBvoTMSg0JJKOFSJH0lzKTJBiIIuPyd3ObRqyw5RIANBh
udeYaQJ/LFowuJCD/2U8SmoGTtl8ywqSyv7YjGYdTeNm5AYKZBXpeCeDq+7+npjdzjyaXeoW8TM1
Ek93LbCYctG5cWB639PTu3U/JGEoQbeMj7XG9oAPh9yzs3+wDxqBCrWPcBdGh9T0I/Ek68WXOAeo
v5twYPr6iCqcQdJBhgrK1opQFdaZLjO8Rsm3maxDNaUh4hhi0YA0JBqvb5GLD8FlDbJ2vHS6C5nX
gULxuFtZuTnIh10VTXA0j+m3rEHN2IrX8V1SM25Pi7awb9pfYEqVRMSBV4HdCt+wSJNrabwVN4gV
RWHCqI3IOTCgWlDt4bVxkyJ3Telf2qi/ik/3SujO0Ov4kOvtyQpVVJtd3djde/CMGbsCsV5T4DNS
o/K5vTApNIMRG+EsxJAx72pp8MqFU8k12Mj6LDkgRqVJL6yzk24zsE46/vQKITr8g0nWBtGH85/8
+1hTsCO5AR3iPr4grnV4r8P8PzxgTAcDYK80TEYgq130//WOhv/Fs4v91kZfE/xAygWkdTh+MVkY
2XqXji8xzfbDRBtpjZh+QupWawvsImdV3PABruSwiB5tDcKGlsTA3yETKatY5zuqzPTPNrIJ4+zv
PSSho3NRgaYtSiFdRS+bunyRdO3nIT9PMnDHtG3EkFtwS6npLRqi/zccaWzlk0MKmyyMuHkOInrS
2k5/+qrKWx3ORRiJvqedgmntcsnGa/pGRzE+mXKfveEqgYJHFtXvVOvwONv7p8IVv5IjuucRGb+r
u3+6/Ma5dJJXtUvySKedBA3EBpheGWFYC4LqAXOviQE4X3+UJkjIAPkgVWn25DSn9ICgrbq6rIbv
AedNh87Z6TvTXecnT2dIsU6A8dOT3aDf/UI0Y+on96YI30jiUVbbPa0p7W+zSVyX4xhMbVphZcOP
4lvJJFmmG6OE24o4g2iRuol2UqqxyWRm3enQB8+Wjqx8VlMCsygtbxjYlTB8ky0EuxJFETbTJ7TS
FqjwlWcqXf1Y4HwyFEv4aiLSAL87cO6L6XLA0iuf3yEhxEJSYhqjKqmGVH6iCar8KQLv5CKlW7Aj
AZKv8Fa0lgghXEUUA5yY7QQixAOkOfarWInUOa30GNRL6iMUpy0dLZlP5zalEsA3c6ogybktLyJY
Y1k5empk1qb4251A63ilul615q7Pjr4bNZafb8UP1VSvJGlN2uOYb996KWnP3ugT31g3LStMtuGV
QdPnCo2BMA8pQd23FEkhmZv9JFrG9bJfCcRfusxgG/9bGCvH5A0YulEABZxGS/uVG1synTq18uL7
bXG4Jo0nAbDfHa5Y/1YVoP3gA6ISPPoFSW1cUiURYv5F8oathM2lyaq3fOchrO1egAHqqnSl35+A
8uAz9ze+93Fe11gmCV477kxkWyexjl+QnTE0d5UU1LTBaCYpNDoobV3KgVLswRtFBgtp8P2UnvHw
C7ZX/Jt3/G8Sv9J2UQiamDuJyAhM2aQTHNW0p4Rp25Fr6qUp5MTa9BykTTamx06JCdZz6p7dusTj
4jWtsjxDR0b1RE/D6sfCHfx8f7Kp7BNTJPds4DVscXBEWh3GSL5EXWuK+ZYtikCKMCmbAca11SmZ
MOmRu4zqhan6O5zn5wg9bwm3uG1x3sNv6wE/p9rlN7Ho9m2OLFNrsR2xIMgtc+huRQg1MgBHe5ZX
du0bS1H90BDb+uskUbHcRMiMebAuRA/sTeD4Ot2KqBKLQN7CXNyVAhhKYglvNh9+wKXo6vz/knQ+
xHTgCimDewlrgzz3Co56XN9TQ8fKeBNe5PpiN22kudTGD97+YwIp1IpkFAraghX6fEiflmCbpTJu
aSv7bpccRnZD+wytxM18tpetRFA3HC5fooT+t9X59dX8gz3zHpuUKAEaeDckQmOpIYd0rYw+3lIN
TRX9aS4FtGSU0yKBnsKDMj2/WCD0noC8nLILSQn1vMBurkadDZ6/ArVUztGX6hvbWyWzEMOYmTR8
f9srHnL8HoFQe0jOMelLcqVx5aGFP8VvW8ypO6RLNUGs0IGtX7Y17bvXtTLrmmbK3e6t4zf7Qmvh
1XRX0vmsGZB/ovxGtKhEE0GFa5U93CuLfbAa8mSH3n3MueTwgKccw408i25Vuh71HKUf/2galxXu
1EHAdR51W6J/yPxsdoJAndzGtRmJBrnKXX55iZ+S589cvnhL44h/OzXcGuv/fcUu88n+Yx7Hp3Kz
N9ZmC/cRHnMkJD7a9Ck3NR1aGGl3zQuysPPtY3QnPgtDWWDdWbFVqCcyaaZHKjeL/BLeweg1mN1H
8813dMIc+egFm08JSeJO5bz6rTEylA7Wcq3UMbpcDZzml5Yze7DP2gN5DMum+Bm83Ms4M/OkuI4j
Piy1nfT/Iwn1c1INepxvQ5ry2UqB3JFBTKHPKsXAwrEzAitx50BpQYhUPw/48N0i+MbLHiA4RVXc
TvKd4Nb/PtXYJA4zVu8VIxTxwIYFSj8n3HOyGmSknpO8qWIAp9ZQrkWx76j1wbJHOZUcZ1yViGZd
ZOM8Dy1YDgLw4UHgArKwZNmkQaeP/1UVAHy/08k3vp5zSi2icgdsKbMrh4dcskzVVY6THzPzF8QX
5ytjNpogyLaYsv4Vh5ctDocPsOkOb+YMvt14QOTA5n+8Z+Zlebl3tEryjB1Q4F7kPBKa/5Lr0mNn
T+64ApPCT8gnD77xjyZkVFsf7sRIiQHy9jwKi1ZaJSbdZjxOBfrl14BiAsfNaQBIDMY/zFkUVCiZ
o/4VB4X9IABmtcHqs1i1DcnNLh/Z8lQlxJSS6ndly4r5YjlJtLHKDNBeuTlVc77UMf5BvIT/V/wl
B/Hh0wyXXtlYmFrjR0aqmzoNwxcvOVw7cgIblh9Avw8jh6GvUBn7LTFEhJTk03mEH/xd0yyBH1Ah
W0eQdh2W2fZvbL55/1m8fh7F+Lz6waG4RZgyZ0IJC1Lq9wguOInDDoi/ekYVGgkT48L91Y4MfbR1
rydXrdIKsZvEe//Ol2YwxQsR2LJ5Dj53mqWprnkWH5N0JXGTI0wQaoWIyiLlIQMZWLvKFiUTKyTa
0JN7lee/AzRukZGjHm8VF3I1r8csHMuJU/f39fVD9Xgnfvcblnld0wQv9W3CC04UrMAfhPJBU1/6
9oZZzO7D2fDarLOKfr3AD8QKHob3i0d46gabj/naslRELpB4mPULv2YUqL/GTYINSnNXfTfJkgj5
7ea0/6DhQfDnJkEC42d6rvNWRa/U12BO+ERL8jmlOgElFWGuivptZ5NPdkjdgnQeBxDE5GdobP8r
aUKt9Axlr0764+Wx8TPd6FFAWejFUKKEC6bol1l0jrA/I3Rxglnl4cA/gS1M5dCbgo7c8dMjLGfA
3DUC+CPqNqXqy1JvJDpzsqK7Z5nyn7FHuFsg2BiT2cJv+k1555dJK3jaEq9dHMlTnov0BjztaU0A
SvMwLSHH51LN4uplknJ9WwdDJeV6NpNZlLFAUrBDRBe/tRdHo06gtxHXiSKz1jFnG3/c7CTkxcsk
oCdJsa1cb/7Ee9mvPk7/LqNykw8nXBeJbFJHt0mhJqq22BGe0pLWaQcYClDG2nwTncS0dz/3qHRj
bSfk/q22Lw5JDNpoNbdz50D2D2ASNIdbsndYfU5TznzEpJZPgaDPYVxsxK3f8nvqkHzNOU3ReaBJ
UBvur0Rl2zRWRtWaT+oPuqvnCf1VfGgN/1kkM5iJJAbLe4HS/0kKJU4G5sguesAEa8rXHz73tizN
t5MzDYBl9otZAcq18N+3EWenhCzscdx7HIZ7hbjuNq7sQwyKWBo9kOaKpRjF9epon+lZTJqQsG7+
99MHN2BlXleyi7EATAgrrrDZhiH9gDOHDl8Sy3hcVzPZROqolwv3vxqwksGp3VlnWzfb0B2OB1Zo
jZqQ2NidEOljxftd+OH2N0+rcDh8qlsi/TwvZn1Yle1CReftPWXVjuudO93Efi9IzUV7ErvpHRxN
bC01CwUjJ0zcH7QZr0F0S3TFNihlbUnHc1RSBEboErNSTI7yR7JBn3+iLhMf1nXPRAJDOSU6TNQt
rnSXfpxt3qbhpl6ybaQRwxsX5AQ9cq1aM9byy1Q3RvWduqT6dkl5UwOv0hvFNcguADsz9b3kDmpE
sxPD5/+zA0Jtjb2fAcchkGvKyOqApoxh3dl4rOUMwATcvl09wCUTxUDl6sqhDH2DRiqf5Twv4mWw
QAanFst1c6cQxjyeDtV/PvL3rLLBn1yoCRQahaz/iOksZFbN1d+GLMSuhoOPVPDe9E/bgn/wRgF0
XJR0t4OSl6f5soDQQnDQKCb7dZLXwCDAqsbZ+cRXtd/9S4o1G6HHTaBrsjVkpULCivJ584InoaCp
i/Wf6yqFJ/55YNrYRQ0+sklXZ5uP/cFrx1xVkgKjgr8o74WWwb5KoJL69Fd9kodCPyiH14x08LOb
083YKFv/KeyQ8pyatFuIsiYJzo9UwZjh34Ox8HDsVd0I/pDVIgSp7FcdeqyzEcu/muP4fVamVPu5
dmmqW0A4CQExMRHCHMtSdTMzXPS6fOJB7K6z6XIYnPfghZxhKs43zs9s92DbKf5rgZIqx5xK/Rl5
FWKEvXOnUXXQJgy3TyJqYyzh4MA4MY5r63aqcW3vcU9PdkE8E/ktcl9MadcFP9MdtwMoaQd+XCcP
Yn0ap+p5atF0y3cx9SOaviTKTEpE0XzGWjJ5Wff3synzsE8+i1Nb2oylhUO3cDqpBlBxOSbRX9wn
WeTV7SIV/CUu3upW31FFsI6w7F2VpqAA4vlK3h+UjgtVcxHeRXe/RtgRzL8JRbqlhfLlCifbinL+
lGpEYEOb7D9INPdvjMiSk52CLNdTHAKkbXHJwzku8B+Z2JN/SPKI6MBoSwovCfG0zSTA8w3tDgPf
ituRoRkEUNoSxD6Bgwm0xOcDsqnViZJe8yk0uvtmwO0aaoXjkh78GWR5xm7igqVfRY3z26UFGg4D
r0wPCfg+32I8SGCOGoSHRNRWJPgEk3eWORzuewOKE2ykcVhXZMxuk8wa02MBzOcR2oL46g/sWDGp
NmO3BTwP5oLlxSbqAvo+FkleqgcwQGPvDMbRGEYgm/Q4NKA+bEKvzPtUupYJYBPDrmM9gSzviLCT
ZAMbi63dfszXkxy8vA6QPVOrH8ju++a8paghzvV+7tluvhHM3uzJugO8UVIvtIfADf8DLOHXBSmk
ZRUTjYyayZpWyktKG+WKXlECG9gjubTjRic3VvZD6JC5cwmjgni0F1Pcx4bsWw+ZSdlKw7zFahku
+wix2h0wIX3Gyyge7ABRQY85F80SE4Wv1PZMlHhKMvwIt5bk9IZSo3gcyNNaWQ4hslcOsmQ29nH4
xuIXxFmtp6vdNqaI/6P5ITybzhl7UwSkq2ClKAj/cpD7d0MDRTDOdotDR2KLzYpIf0qAVAEkwHZ3
F/Wj7YuIar6K+hb+M/FLJ1GS6uXV1Se0dUDkERLbCUbmasRdN93BsIXVEqCfvH04F9P4xEek+rB3
qibCghYXJynJBo7vqXwl7jKVZjdmN5ZcuHZv9lkBGVLNKJhjuz5HUNX2xo97QPZl/bfwlZzLqQhk
wi42Ofxzmz3wxCG1L5EIdzaOCmZv/IResQp8rbKeEsOLdmju1fTFE45eo3hb3bL88PnjwuGKej2y
3K/zM4VbPXKGsp555gX6bKpu96owE7ALJDjErWVyP5Kt48hp/cEhuqA1HKF52acFUcbbHx+6UREj
G3nydwwE/q/iOLFd5TorjbqWVPSwRniXdD9KNt/XYJlRH56COQquTimF856ektlymNpDKIi2lJts
9W6yTHN3+PL34r2F6yMvBFjh7OcxNkdoyoMNHcwAe3SVy6oiRtm/O/VBY+Ei4KIbDao+dBWkDGV3
U8IcvGOvr07yK7j69+K5MyVVPBnDF2npO0/N0PfN5MORD/NR95KRDCd4xmyFGqnTImGHyLibZSjy
rhJrdkB3zotGSk+g0RFYBqd3EhWjF7bbPZJhxaekZlkRGeVC6Ezfzr/wO4y+yVwAH7mpd0pLubpU
oGnuPD4li4rYpwhHD5aWKKdiEvkE+UbrPd7z3PiLnhrIPC2j7OI0vDF9BHjm0MPWRN1ts9OFCyqk
vHrNSqh3AM0kUg2XC+paxhyYq+DeAwSCDIMQQ563jE0qwt9RYuIR65pRFp7R1Cy+RlC9PEjmLYci
jX5mIhwWkogNnRLgAcMFN+dqqORqMUxnD2Y6W3ZNYd5ryFQwqeyAlwrTsJesIfcTZR/F6unsvflu
TmwLe0/fOzh6KXsrbiVuSNEdD1G8AQbjMGev4lfd4yH3jNZ2XJS3BITaHS4PcH+ZXsHdgLnSOiBd
OhWsf8WcYQ53LYi6iRx0z0bm02LCjG46rDp5ig/G13h9TQ/FTib61QMkWZvxfammn6IgVUofO67w
DtdpOLUqBg6ETpNXt2yoso4MMZkJjACmJppazDg/2VE8bNE1dk0yPjTjoAAl++aOAkTvHGwQEKNb
apQdk8t61HucdTnPiOMPKNBEiu9938kt1IjuFq8B8bzxhdLc3LQsLSsavmujeiKTy8sxkbf9i8Hv
rlBzXkI28u4mmV4+Rdl0p8Idfxvikm/13DS+WF0/RJ/dFr2bx3edGdsEVv+8H66AOKwUyks1N7w3
jxqbL55Hu1cda9IG78URdRWaQk/Kd7RqNP7Di9eQlaJwKdRDlndxJ1/MMGe4ke2eie5s1znJhd5V
GFDi6MLEPHA8IAOqHvB62gHH8vTxLX39O3IH09fRQCzrG4qadbSy2LN4gYS6Pj7vy3IpvI9NZV6w
NsLnKlL93ZDMqCNSp2H4HapztMv6DTogSCY94Zskw5xUciKHSLZOfW7mbrwZtXITD9GR6UxD2lDa
nlZy+qatH4AO6p5A2bATIA2TYIVECNKvGvC0BH/2Ar8a06g8AtGOJYmmGLym2F8pXmAtJN0X3JzF
VYKO4RUfO5H5L+5tFYLAxEzIRAOEgugr9qY+2Dp/Ss2U/FjnOSO+cv2mx6epmD0x2D34zgokhZVB
piiBO33ojHTdQav5DSBlJi7sgqvW4ZQnzEqks0El7BaKNHP8HvRbQ4gG2Pe/l6E4+fwUJEJ4c71a
i1LHuirWHA/bGOXkAobizNvZ/Nv1S8cpRh47kFpbdKESHrZoYu9Qc/gMcYOenfMH0B7bTekCbEWH
Eejhp8EyGHYfev7wBFPMiCdwniWuL39dT4i39/m2kEIsT6NA7cPKYFr6iOn5virTOMWSsVA0PhPm
ngfKQrjLroN8Dv0ShqPIEIrJC+QFEZtDuXFkBk3gMsZDPJ/rgVI39w5wgldYAi6InhnicwO0p0Eg
kqnjdbOIjQWr1LIvzKX8nd7/nRtFKTzdxXSAH7BHUJepvSIJLK3jMq69sDmggoyIFKWy6F4KakYt
fZE7mPQZ9c3KTz4+4zA1QdOebokpqoWnr3TQuh2p3g2VuKsrtuyZen7T73s3ljzlut2sQyxrHAHG
cPOuIGyteuhdRIQ5lDqOvtsdKip74ZCbxsW+zaVy78zXhp7RNKseqV3XpMKWSOoNhxKNKR7ls5Rx
WTNCyEh9aHYJBendgW8nsJXsVzeRsI4Q2JaET8iJfPu9HuE4FcpHOdZb1p8htkf6DTuwAdj3+Lnb
OlIIg/x7cs7wo/n1Acky3maetO3xoi7TkrITHAYaGrMxcEimFu+oymbxZp6mRj+aQ7SL4dz2uEeA
BZbksDXvAeofcSlRG2iG3l6T/1Nb7MjSXk8A8uClyRfBKutE25aBAUud+EgrK/m74jh9tm6g5bsn
Sgl4i040dRLdmc4TrCLe047iCqAqt2ed29TkkBL3U5Z/o5vT8HDdaYi0uE0aY7beshic4J2WZmyQ
qWy2Dwu8RhmWLIAjGRhWUIhw1DdCzRiSC7b7vo5xaFUw1gSS/iuJnuCtpH3NRq9OvohZ8wR+ms15
52yv8tNThs4Xy81kPne4s6Oj4vrMYOOZlFjFe61yixxIrvLv/3ZpHnDKbx//ABTnEk8aduxIgcqE
y39RYswIXJuIs9wQ2Q74GKf43VY2MMQ5eyVbzKV71POBB5BAGqkpIMXgDfa1ERC6QaVr4ZDp3Osb
8WnbBhzZcwm8TyaIde/lJal+ejl8+jfe+esXx9FFEs94xMdi47WEVSu3Z6vlVxRR6xqK0Hyso8up
ulGeg1ea/FRgKjuYruAffi7hcLLDFPvmbgQWQL6hOusmisfR8pIG0SJ71NFq/Qx0Kj0I6oiZWxsX
lAshOxyPfggaNtqzK6f5NcTgJNKhg+hjCp8nkoCQs6R0kqgIqBRZZhZA+1Adz3bzpalOkyxBt+i1
0E9XK3DIcm+Xv8G2HreEZyicDtN6/1rwz3tJWwhPhppucbBypGm/evFzqbjGeUO3sOYfhgrxycs3
bG41LEBvlESJlDQ7el9SPTaE4QwIYK9VrI0is8Bm5YkT41ootTU3Nd+yo9dMFL5pNX4G+AFYMDBM
J7wPLUSxEKEQZLdqIo6kR6/5LzEdYAHHhKBvALg3uWLktn9pVdWYyRvDaQW0AlHfxClbd80gQR8y
9Mipfu4Gsg2sr9UvIik2cbP6Ss0Elbaof0lIMq5FwYjzWFxphcSF/2VY5luZeldvWIhwV7SJDA6D
xlEbrZIWOa+U8DefiZid+fF7O1paaPta+JKqPq3WImlX3wsCZPtV2ImMTYEnjb6cRNOxQTKqrWsH
RCdh/uwAurLdLbl0HPGM/yN+CGi+KoqufiwyflFQ467ae9fxZ5zPrwI3zvLMA6tvwTRCBy32NjLL
+1zLM3WNVmwB4waN+CN3blzNnaCryfqaCHFO+qsQqSdTJrQ/db8eLPh452eVo3szHnjg6qsDKdJD
TeHCfHZkme2jJZWQVrlHYozm6L1UiPh+bf3tx/5DsTsdO/v4n5fllznDkCJJnnzT/BcjxXKuWuok
5yz6tj/85LVX6yIa4occKDTfHW4NeSBqDVB1r3+MgRdH7nKEvVLj6YlwXzbVKNGX31XMjty5a70Z
jtJOPO4mtxISjTFXrM99qpkCRS9BHXycNy/TZsRegtbpXzF53A5CUQpcM1OaER0fcDXmnApPOIdX
aqah5ml/cVOFEnJRKBdX+BdRXIHaQHDiLEut77pEpieiGNtdw1wSNZ0xoXM92cfi3FC+rNTMMbz5
zI5MaP7hkbSpE9uy6IdtiKcP1KWiK5W3+ZzmLAZbEtToBqNQeFp3x3Smyx0BrTto9sA2kx21KCW1
nRP4dTu0Sn3ORkQwQpfKDrjgm3GuJ+Svja1Pzm4LrCVD/aqnb48ObRgq7wmSA9X2aZOM67a+BoFL
3Z7Gldv5BBnaXsuot1+Uz/+0jFg7+lvitNDkC98GtEe7uMDyqUrF6DBNKCVcDDJa+tLCNJQdVOpR
OvvmmJDyaHe8l6ireqgzG2TeCjOGxKEX09aBwmGUo/4dq+yX8rDWR43SA65oKOVxavRTuZL6wBMg
QuBzVAxusk+YTi5uI5bLq1wJTce4AZA6Zh7mubmyNX8mr2LIq6YaK+g09wtQmW1ScBhP2ZH5udB/
GuM0b/i/5aVKJLTtr8QyRZJZ4B7XEu6l7aVJpQZt7CkpFlA+LRmypqLSECDc4/T1J6F8yTX7sjpJ
9tiZCOr3A/kV0qye7s2gW7tahfeR/ffPhKC3utuUNbmCKOWGJ8SyHGhK501br9KgaQjTiGl99nMm
5jyCp8Xa1ZX3fgD3Sm3EAyFUZifYn+y2T9tQp0rfyMcPsAABGXgHv/bXU8DdmtZj1cOh8izMKO7a
JIJwxvHXcYGY7oIrTuhIYoNKus8KoiGpr4Py4NkGPOMi260Y3A4fLL8XU2kf2+GUAoLVijc1njbv
hGrdsGiX9w0XLFVqcvsdpzo/f4u8hlwbRz+5r698AjRKSeKIcT7jyNC2QzAQfa6IkEu14R+oO4Lc
Yw49MxyBLJso2HN9hNr1cSLvqFcbn+SHsZgF6EbDC8YHaIpsRiaGTLpLOefE+5psWN05FqJdc5K0
vBfLDUo1tpZrYtjjJPQ9eREWfp5sCnXBSL8W397CsROklnKnvKl+eRt8jovmGVO1R3MFPtOPTY6U
97UNYEnf4L6DZAcpczAuYKZcrCYHkn9oeExSvUvntPQuMij/aNiLBd3Hp1s2UhaQw2cGQJOOBDzy
lYiNSByzOddVPhDaruXN/r0P+z/52V1tN6dVFKkkqWr3glY+18e5q/+u+0wPtEK9gUkEDNPJyI4a
/rNC3BTbLZOgmmyGeWwMjOYL7jWdA4lzXyMVk+UNuz66jGjUL1bospxWVBV2Soq0mCDiQRHXOvPJ
9fHuode368KFs1M0A+VC8mCAfJdukY/0W7uiWbqGZIeTdNadkuAEUt/HfwpXQsWAY8dyJWpmsFDw
VV4LE5PxQGfBqtkcKpcUHAWrTkre3pkP2q6uVoYo8VZrGyskz7BarA8ILqiwdApPjWPKdeFgyjgv
tksn5LiagnDCztUXkPIl/1e8UOXw17PP/grQb0fObDPUABBAxQy+P1+yDjbZi+8RjgWZcx0Iz+t9
UcwxQCjzUAidW4xAY1zkgbzEx6rNy+tZsN3h19xs4FZKzSqU5CDL+Cbw3jh48RCL1mE5BQYIMynW
WPgqDZJdSFa+6x97LqN7P3LkbVhkFB7nIEF28hQysZwwF8YVVjIt2DCpjPl/8uSsgpv8T2PwFxV9
jS1GYNemvDFPXnn5ueNVlAcZyrQMNR/5WaSugdtr/XFHeNjQb6ft16lbldBvTy37m/SLtqnffg7r
LADcW1YeYbZFQXo37W1qcY9sU9WbaBawhHMndZ6B9PQsISOEQzVtHw2RH8b3fOw644OCw+CVVjsW
9jUptDVU+vNoYO/fROaKIbIQ1gXNRW139zp3OtHIrJgi7qX4Icmr/pUuDGPbL1RIekfbH++bznzs
ghcVytuPZg63SQVf3xntgP116bXEr5HuZZtkWxGdGmjAt7rtQQpUYw6XnclNzuQnToWaDLr0l9As
myr7fGICPOdKy2lOKkzwn8Ra7hzTvizieukiwmJi0O3auqPTBNC8z3Osz2JkeGfbBsD0cDgHtF5h
0CkXs34UEAw9IfVNkXXa5IfhdygmANtRZ3iOm/GeJf1Xil7Y83H3xfal4Ia4iPIGbndDOOt/ChOC
R30ruxnXc9ekIqBySD5m5uus7MVXZSaijyOAGFkgfRUaXUdLu7ZLnZYIyesWnZN5jS+n5Afy9ScX
xvHHYXUI2c0tHNnROck96chYbwIJ96SlnSN3fmkj+gYCQammZAqoK4vMNrRFCBftA6h4J4sgQe98
48UWfdW7N04k+1WIVI4L2w54UU/DKhkNEDIDC33CP2DAIoDGPTAvUrs6UUE/UfX7R8PhbCktR/mm
us6c+WjYfZ01toC4WhnABruFvpLIdu9yIHjjwSmLQtpV/FsnEMomTJM9y3gu3+ITgu1Lys5VIUBD
FgFROB4rFxHV5DfhmiPCff80j3O0ESePRwOJVNTULj4ylV05mRvD+enMviJXzDE7iMw7qpw0Y6cG
WJ6W1b/kYLjyef/hoSTgAcWmHEKOZba0MCpgC1x0G1mWJsSOQnvMkoURaJmhixXM6Wy5rU5B1/7w
nRJtdZYAWXe53bjxxtXia0k0sECtop8c4ceZRKGXQl8hYNZgpuQYFjpv8H3CrL2uCojuuWPKCo6b
UGqfueyWyx5NGWmFSmP5HCYrZklL1YQDBXjD4BcLamJQ9VkMiQ+xbNEMi8P36EH3IUCo5w8UCRDR
6hE5+gFy0VaESgI8LYHUFIMdmABn8+AkRJ0EXBwolpmGKPBOEohh/faOgIBmOIvB/IXLHtVwX431
bz/F606IQfXiK9vn5l/nhKst3PQ7ueAXU7KUY/WaLEK+C9uIuCJQMMg6OurpiI+dBdsDHW3+Eyfa
7bnm11HTZ9kaGWwbTRuX33+TpeYeb/qD6mKk3prslpWok5ebv3Zzle2EtYeXkQSkZLBhp1Cmch7Q
MesVtMY7akLUw5F1bXx7P8FiYaLQ4u1c39CiOpfWfm++ItEu7IyhpeWuWnWJ/yH7i9k+r62JI5vD
72PaCKVo5XU7pOwi/IYymWSeuNdvrjFHjBHZOCMvyMk493fIyImyGeSh+y7kkDET0y/WLSIx4tyw
5XsaBbPXV+lMH+vBdKLiQPs63ImunO0YX9HP0QuLkfwGxpnGqT8c7pNFNCliqMlTujaN0oB2yR7l
t8SOeYWbfya+YKR+Y1cmgZ0yc1TyWss5WwSM23MMtJX7CXwkTckkuSXE+mOCJlleDLAVeZM6VEOm
NNPbe/Nu+/22BKnyKS3fVDAxdNIezcTY0LTnOobXb/FnIn1186T+6AZa0Qu1UA3A9tvcwcw1e7Nu
8Zk16oB5d2KsQG7y1/sfTF6P5ir57zOlxFAfUI6cULpwJmofV9Lr0cQEDR1F17JbL1jG8KTR8cr0
pcQLlFLafZmb1voOZ54H2symihyascTysJ8cYoGOMWuY8zXhJGZbBhohEtM6DPVtQkPeLnd1gndn
PZBHY9YFikmGw5+ZKjnupC6b8dP0WXec3DleVf1C+r5DL4k9Po7HoUlXUrLS0zBepD/sUO42Ztip
4BbPOHm90VAXyroJl5WLSbF6YWKkWlHgaleMclH6r/AA+3jT8P9y2fuzY5VqRMrmbCNZA24JhOTV
uMe2m16Kz9bxPY6xPzv4H8lokG12+EXyNiYR3py0Rd+kqiPAtLwGMYg1JJjFbN7NQvd0DiBjdOnK
Vnk1rGdW5i7awOOjhzhiu33PVH2407s/Kt/XGSACjwriOacWTUMZvGJCzDzg3JsYLPNn5j5qSYYv
wBp8qZzHPB8Qpg9j1OxPUd8D0N+csc9ym0A2PUWsOzW/hJYM23uZN2ZSdSm9yZKhNq3zZ8GoIqsu
ybhkkt/SAJeq+15wJQIGpW9j1bro4A5MisW3MBzV1Leknzg2b/6zrmuEe8HCsSZFd3zT/53X7suu
tyFklb3hj/PAL+ZmZnfWpkm2G7+veQeN4phwMhPnIx/+pV2hQ1WX03RBWEcQBgZf6YnWuNs2hv5q
mtYn96Uo+z8JmPlwi3gytaIWV/5MQSqKiOPtsS4Wmkw4kdnoRWPn1x7ERkMmyQhFKBYZmFx8YkOF
tFyi/03pu3hn4md9Njlb7ASWL5WOi8kQvkZaxv/9XzqSRiQKYAqnMhGtNIjsMLzUIPvbYrIpzi+h
z0v8CsXIWeMyaTBE/fb+qoZ1AnEatBoKQebjM6yywyaJJhlJNxFtvYAa7Ft9qunkQhaAH+cPDlY6
D/59sWsEIvkMSRZR52dJPIvUJqjt1B0Nqvx4x+0RIu5AOkJwBqyBDgSMCAWzXF5VgwHw3aqtzdIa
Tkn7Z/BOWmpnKmApV7TvXbNQCYGdrjy1OkkmSDuUPsKn8tep88HuHQDmVfqf2UVtuahLpYe9igkP
RaRa2dOsRJT8tVIdl37XxInEe1nSYl0ON5p1noOAQYmfH40jpSvrvDp+B6/DXoSJsf4MA8vhkuvf
SU6Fie+sIXuuQxHpQ48vXRL2Cv7LfCy3oDCkosFKviYNjbhrRM2hyLWMyFsJaVrIhl3T1i415Q/q
s+TQrFkVz+XkvuVxffy4dlDrKmcb/mJ3qtImVmFncY+XCH7aJ94zmYeWu4MGDrCApXn6ERdZT5Qs
jWFCikVv+eg8cWDiXU+pvUgQBTEfNcxhMvS1sWMPXsBGWP9ngTItu/aHqE/trb01WGfu+MAnELHu
cO4Nq/Cv8IiZJlEud4bRH9jIL1woovuNzrL3QEB96QnPwSSuuj7qLepQZ6Ox+O2Uv+uCkvzZ3fS4
Xc81eHhSr3i96gxC8EwUEdHxPbfb6t7a7gYhuLABpSt4RWL9KFTdK4R6UtHpl/RSgQNyCNegDp1T
QJFK72yXtasNZOwdsMo2CksQWFSuUtN6JHwrltuG4//drwA6xQCqBMd8zpnVvf1BD6ayF6S+Foai
20XtVLmtwMzjfWaWHIrmB6HsGsqMQBbikvYPg2uC0+bNhKZKiqufLUIDL06W60zQyPG44xnLE86S
jVJaKjt7bw2dxFL8+cjoFdTksS/Cnaw2Zhd7uRnC2vqFZ/eSvHt5DBwcLqiiwqM6d+A8XpjuvTYO
8a+6Y3m8xUxuBuln8NfdPSA1mtRgN39cYKYC4IFW8x7DDxSWuNarxHTFMo2Rz4aUASL5gLxGiOxY
ehpgSUtOjO1fO1dd5rBnjgaPiBTepwwEu/egv8/BrwCIzh3i5xCNihn2H7z/B8Dt4KgQ5tqikjYQ
0Ck4IRXqqMxBeORdaZgOAI/B1ZmC2BmIfYcCHNj7hxk71GAp842TSzFnF7248psH3GarpFPIdZjP
qe2nEXR5daCcJnfhKPlR3sXaDiSabmFfT3wz43TjTPgFacrbbewbPwJVNDy7GKVB+aTtkePyPyMy
4KK+Ym19cM8yFv/8fnJIccmmcxQlZ2BBxJFbAfw89raVufgn66RSlUedWs3etkbUwrToi5G0EfJN
h+O4o201o84aEqx0W5vjl+woBL3VOhY6pns0ykJAF3ge+B7IgQqUVwNevgl9vrsgQaUPMzLM5RLd
+yLKeWpyuRdWYkD58AEd1Xv6o1nhSRVf1hOJSh7aijSSYWWfebf6VbzPQRFJAU2dM66dDW55H0w6
a2GKJaOrqJ/rHnuIz5a0WQMZ+OI+IWQMjkRRGvhCBmG2NmghDf7Pwkkmfm4qKYckqaOu/E/0PqZr
DrJahb4EyuNSPNPfDMxKuYOxlnutc1elwXI09loLNwJpViI/9kMChKNlxARWmFJFeWvZKaB85ig5
GH0wk2d+mMJ8ZwwFU1W0Y5hOokaFIzRFg4/cJgPg5eADpi9+5WlntfRuX45zUnuY3NBsjxDM0tFk
PkSP1uPINuJuFPJYh3+YwZT8zjxjeYt8C9Pew37bbPXH1IQPgHQFSA4G0v1mVFh8NfHcoIQddPbo
zhiCavGxLxFK8RteoIt65pFJuXd7vIX6BIip+LIILiOPMEUESgjqsMBYjU+6w6z3vTSgVHPOtD91
hJcwgQckRuN5d6vONXoseixsT2mpUA4YW38apLYNCy8Z96YZBZz+shLY17P5MxkHbicx6tP4u8fL
Xgp7mfBGeDUIsu4GGXfhslrsA2BE56HmWJg9N6Siq1MnPxJI+B4AT7Dww2FAs3BfyN4E4SGgqcQ0
RMPeGYlSR5Zwfryc7jUH+JUBwnTc1khXFk6qsY5haH0EL0oUsObwSLe62oplzkICW0fnF7duvNiM
wyfncxk/3HvkXNXACo0UzYsMjjsln8UU0BqjbZ7zXpH4x9oPCcFMPRVrumm3H5zWtyiD/A8k6IQJ
9jt/g1zvkf39vlAVuskIL5qsw5wp2xA5v2hQpGPTaYeYOD38QdbxntVffMPT7QRvGsPsk2s6aPUN
208Bqe49AXH2VaUaF9KPB8Q8emWhTl9NBwlT78IT5x0omdWbPbdW1VXYFcqupTdSIzWcQ2MgFudw
dWIK8s0AyCIBITzH6pKxjo58XtzucKi7LR5JVV58/kpD8T/mm5afBs4JhT3ZdoG8THjJG6aYfftr
OaS9cxDTzeCxOeDKMNMlLgsCPjHUNj27RtZzHoe4USeIvldtsPAuGtVoJHrr1+e8uDiV6gi9gQb5
J7at0vUsK/0IHyo7viRqg3Ngj5G1F7X/ceqS3BP9cCh8j22j6ksBq95mUJfdYUKLBiCIzI+WxXgy
qStCRwINK9i/saj6jYbK3u84PuvxjzwUsRUyUUodtOxvpmmAGKl5N79ZKz2QAvHIhLJKcMbAwVrx
8j4bcp3mzZku0I/3NOeVB+aJxhCA1x/yJiwXIUl1J9f329DRGiqBR0nFMpcPPD5DzbTVyzDfjSNG
ns5/pFapp+SnCd5t3HOvAc+TPNg6F1lhShidxkEN2rku+wntma4o347TmsP2lJWiNP0B8zWlyCH6
FVMeOTD4DIy5OJKEFUgBJPItwx/CG/SthJgl13rg2TRkbrlaBNJ4NFLC6+mVR1rtqHXzdJuk3foB
pdQmr7sJWF+UcgT0ifXM0k8BFPwmU3tBKYPXXJrl07CRvkwdNpglX0YYfalhghK9Jm7uZqKUHQwt
rksiCbJPmZn/tUR/LSoftqsDrFsPhKCdN1VwIdS7v6Lq9UIK8Sa189NeC5ugQET7A4SnNTiWgmxM
aQK91cCcORHcKOpBAu6k6WI2kB7c5wEEMl4GQ4ztvWxMqS0yMp485IUYKyvJbUDuAqDbtX4HYOeJ
u850Ffud7fBChTcPAcckNcYHEMTrOHjBYSY58bz39oFuhN+0oZ0cCEurwT5eosjrMyLnhuR7df/p
iO3r6to9RNUzcSwZ2ze0FXh48RwOWUTInyQYRm1VgTjLyZ6fS6AoKTdzPVpWaZOyV0YafF2/VBrk
3W++HOpZ/linzd0Eu06gOIed4pFQGzdip5ccyCZGht/18Lnk5OyPkI2hQAbO+TpftQKTRh9cw1yO
e1Sc9tCUz0P823jvmo/Q2GOaDJGyKGZHMSOfjC+fDcrxjXS3tGVlyJQgNo+QxeEDg8BniFC7dm6w
iQa0MjFhnb/I9s5+wFQB6WJZjok9k03/bcxBxq9Z63rLY8bqIw0JK3ArTm7CfEK4NAEb4TGN+m5A
rBm/BYxqX5Bt1Yj8yFa7IG0uQj2AxKPEnwDLEwsp7ZRZgtH0kb5z0elykLhMzl5/C4OtJgNZIEdA
ko7MzIxJqTWrtgqo5EJkn+AVYyHZ/JVOcsEnFTpcSk71VJD5J3fqysA18/jitqsklhSVqE/v2fh1
5lS5qSDJUt34f3rypF/a6IXvECF1GJcwVe9bjeWW0iogi0fLxub4Gz0KNfrRwVtnLNmCMaKFZ7tH
I1+nkBdsR6F0MFvVUCto0cLiIMr8rqECaAzTkq2yK0sC6M/ocI79G2eFmGtZTB8kZn8D2WYSYXdK
OQKx/SJfNXyuNanDg12h6m2P2lh2qda1qYQr0y0kWzZ8fOZ3iQIaK0bwDy6kOeEafr0w+scRZtv9
CvJVN4JHewdkCZJvPDadmtsXFGw1K0tCdl2UugerxF44CR8WF7nwWjyfG9hlMO/47EbvkKGa9Pqi
fa6BT1OnDZDu437k5jR5BmJU0skcnOPYaZ7nTKorN4De+wXBrLWvSOkWA6FA5IBNkM64y5PydefE
NtVFpHbvFIHVLTQPSGD1NaXraDtaRUpuSF9MH3jVn1yxWmwlBIvp1J/o+cKLSB1ZT2WeFKZDRDDr
L2et/KR+TVS4Oia9w2gyK7RJaCbdAouW4ynpQmjXvWc4JEJeBZbXaVAVE3aEQrng7fmRCWI251UJ
DdpmkIgLX1j/EdQzMzlHClAtYBlskuIon8SDlMg3h4bUupp1YwbJexWGsDDzpoEOpTtp7wngLkBI
NZTDIkYOGYXLXLGCyQYBgxea0ZzJ1fXmMXI4J5oKO1Qn+12w0PxRon3ERZ8WW4+rumGrOBNKCQbt
fW6NOpaXwCF6nzwIaapjRmSmKr2ny2H32XJTzVWIVFq5GEvQOqw1863mieowO+fwaMyoGyZa114t
aISlvJ6XPdS/4Rr9Men/CLvlH/KI1RugtWY6t6+9TFSOHspytdtBBDL7zCWD7TLwDCGP9NtZOKwm
P4efhDAlh92bJ9Q4d3DlslOSbVQUbF0WtuLSo2qwOMZkx/1IvYHFDURiOVTB7jWetXsFSQLyzCdP
sTly2zU/VbPvSfNt3b+eRyn45tZ2xFxixxej5bLKiRyNCacGK3RW8Cy34RB+9Mgrbw/zcSYOcsSG
LJI8Lm502cekkVeY0vbu6e98BesY1WLTKNC8dZsRCt894V/XfhncLepwW00zYDGLU8pe+lx60psr
JOb2pB7/wLewdz+pS/DPvj9D7k211cAAay6suHzHQAfmrNgwkdMYcxrBVrUQJCmoi2Q8CU8x+CH7
fxwEZtxzoZLapDtOk9efpsoMf46PY1i3u5jEMxCzxB8YoPcNs/8NB7pQV0I6ck8uCIoAvfEKfPyG
AI2oQ/sXWsKOQ7SZB/YHj7bMohPDuFvgQwSJyw7mJJUpEHNtENzOZtbJUY6dL0Fde/Rl/Jmgamt0
QDlsvlx58CbyCCZN5pipeJ78FtzHgOmyzgk3VJ9jy/MhYVRwAuValsVBwzMhHO8bIGK2KRyQ00Cx
kHTIaxjvhBksm07y+suqr8M7KsKGFdb5YlErKLT8DpYHSgwzOOw1p8Sj5uL3jEBwI1SQTtiBT+sS
e9DP9ZNXuDEXt4wX/M2+kCxVlUOnri2KyE0Sq6rFSAfDzwOri1fkSMu1HvHCnqZt5b4iUVVyQCQI
iw1ZeoqDfD1y3DHpVbIvB6zhPhSFwOom8XU/c3boLBMkGgHG6blMOv7QVJJ2VqUKFXbY8UzlfA08
0U90l10PegzJEsoN5RyXq4Dp/rYGhxt4eqKLGLf8KqQtnX5ktMAomQ9dExm3ww8NCVUkU01o5FPv
RjA8UuJd4ArezUKcrPYLICAjduKeg7UPpxnp/tNswH4+b2JEnTevf+c/tK0J06QXA0HKzlIRJfq8
8PkFBmQYQOE/Gh6VgvnXUEgwbAMK50xK6pmNaaKHFok7C/Fka+T4kMgtVroXa8KWj8JzLvs+KwEL
KRRM9romkETmGtjxlo7moYDlm2qyd74XDKMApPxW8PLLpgPfgXlOomPzxkAEERRGa2lgc1o+Q7qa
pa7SS2bjhmBvvs5Rx9XGnvk44mW31qMdI82H1ksvlk0GXP5Gt/8zFopSZYIJpe/bvsk2GhtIp97d
ObFWDnK7VIi6/+bmJwPypmB0IIb1H3GMmozrmGukr2TpcC38HcKSl7WJlXBKu1hsHHdpp7YS3xUb
rOiz1zLj2Z7Fb/vhzNVAKQkGIpKPqphRQSHxKdQ3Cio4qxyz74SYajNXk85AuDE6g7SSCn7TeVxx
zi32DLw7qsXx+bhQ9rlanmt+ar6QsMJ2JL5hrSBe0g3EyRinyqrMwmNMMzPHvXF2d7bPLkK57ldO
IUOqZ3xE9i9FsjO2h+6hDo55rh8X2G4vHgmLu85rBv0VnhAbD2zifL34ruOoOOt3Rl154D24oyQS
wji0Q6pw8bZllw84X/z4hK1V54HSK0wShMtUjDlOg7v255QWZu6ka2498ZrwF+Lc1Gya1AZL8GnF
NJLvqd3httQCjbrTfC8BZTb6W/tt3JcbZDHssG/B0dCK8r+H60clFafH/RBtQKFLqOQ+fZMSlzJh
f/92DccZYJn1cQBxYCyaU4k/V0EPm4lJ5dH9nNPcKhIpttsDViaDpPs45BCSjRzmeHwdrAtEInO6
bsaXRDrAqh1N+XFF3eTqZW6HQVzL3jRD3wyuCBWLU3ckb8SxFP6yqhIP+PsKczLOPTBwjCsfnl1/
rjHdCJilRvtoNKvZOvLZlgJPH3xOEwd8IYift+Y2G9x2CmQ+ED2tfeJcpM8Z4KI0ExvjvG4dMPJ6
NfqrRU7XdLHA7w2zjAqg0/iibHklDx58KC9T1rE5Y4FN4eE7n2XKJUM4nl2z+6y180d3lWVfjQH0
1OQEUQWDzaDZNqxbBu3rY0y4nfUeaNN9w7O6UAD4Se5kcjs00nGUDhspxwOo37p2FA6sTni2XRIQ
IZAGqHLt4GijUPlqpK2/1E8EprdBMGDovMr3qVRhHMV/kbdEwKS3/G6NXCHPWPGQkFfe/xEQ5Bgu
gQrstScGdCmGNnwPHGHyQ023gKPRWk8+dgaAipJCSML3pbwal0YKsK7Oej3fPN1uCpTSJ1rsGMn+
mTTNNoJnNZApbSVnp6NiY9w/9Frz3htiGndBk2XknCMOOG6fJCSemcjT7k44scSMDcWCbm2BOM08
aGi0Z/cXqMpe9xuIMn50q9Cm7tm8x7Ny8QVgPyUoeJzRp+PNV5SnQPrbf2bQynJbfc8WvVwNk2as
EhI5AFie9BtrBmv6lolHfdsHKhBHs4PYDagsBKlbddHDTvSPMTTYOj6EXIsrBROTnts39UkCLjj/
DA3rJlFYez3B8YCHmPLPudg+R/ehfqwxboMBnsgl35QzGo6WGpRq1pMeK0jnZtVoCx0BYLMJgejT
+0Jv5PfMVRbi1ZdZDWoy6VDL4NGUKxIryk1Vmf2VxOBk19VqSwz4GlwCBavfvfMTffmgW9ubqxET
0Un8HVwTp/+8KGE/6uJSlo2CpbhMKOVkXmTFtRsNrF+4iSne9b4SMGcYUmys37PEh3yv/fgXKvMl
vtV7IovZUSDgOr7O5/ZpW7XActlB8GjT2Kw3P4Qw7zpMwLVf4V0CCFDdMdNwULJTpkqHb0kdDrbg
KYQiRHxbkJ1FfBky+4zKQHSj7l3RmRQ/+0g8PRlt5Cb6VgF5QwlM6naS3MI2NThu/Rtevw3l51i3
HIIyA6biKYYPcXG85nfZgK9pIo2ZeCv6IP6xFQ/Top536kLEzyhBNm66RSabYVcxkv+jfPS0QDaG
v4oT34E7KWwUbSvI6qaf27yemePoKvOchgSTcd/bIONa6wmn+SlAK4odmvjV4ZTcJJk0dF3lNWM4
/SSZS1LRoHaogjDZHnWbX2DU4OHsp+IV+Tk3xY1TzDaQgWYobYgfswK9svMhGzpOdJaAwkb3J+kg
7I2zN0PGrwLSbNHGLEpmsLA9hMY303q2Nfmsg4JBOYPzWQ+0BqLMXr2XsYGkb4ECvnPiMoPMiUIr
JsoWkQUxYeyensSF8carJxoGHABo5mY5IbgVbLmzxcYGSFQJQHvsWfL6IXHS7lc4VwIyKqMaKbGc
iAijElIeRrtxZ/aN1qqr5XaRT2DvQ6KVnZgkJXZ/101wGQNfFNNdZMYZHqDxF1ux8CGFgINYmElV
D2kDQzMF7Mpp/5WgkObCtks7iKTO1CZARDJCSHLt2dDr95cfRdBXQpzsyVeUvA9vz3ioOX5d1HGn
aoredAUveDSVqGMIQuQ9m4cLOpK6vu/HJraX02i1jXilIKJmWefmRLPDnw2XNmW/N0FB7uUo3dYO
mepoX++hDeEJZKjQBsgwIy4xW4RLk80r/VFcl6/5MlsHWBWrFlrpjeaFv0lF492I0B7XsvpFP+nU
JmVcxjsMMd9szzi87IsNbSsjXnYuvubeeLlbAN6EgaxvREcbCS5xZbC2O8CsKFQe18SeJ+RjvmWs
OnwW9RyGjos69X3MC07QirrHwqrHUvj/+QMmNymsqBoxQZxtrduqMyZRtFrS2UtCVSblQl772SMm
LvlSWgNhDCYupWtchuzLwlIVz4vFeNXwmBJs2v6KZH7IOO7+RtYfJ24hftBMs9GpQuTGZTCzKnIQ
lO9bUqFYlDEQZ/1y+ta67W4rwgDafgDCZugQ89xemg4AFK2UhlvLJ2D00DgGqroW56IGZyZvc+mF
n71Qfj+672OUY84ZvNVVgpHueMRX3cOtMoHXj/I9uP2750+dg0itS0faZmTLZtZ2SpHMcP+o7GeE
OOvhPrt4K/jCulKz/LSbulRHoZ817EiEFVUi8YpX3VrO2iu/63XjLjI7kkaXQdKNMXlhEeXyTa/H
bIylO5FLN0pGFXrrtvGX0LIECwta5A7ho3k1E+D38IRO3Meu9Ehmv9d2Ft+nW6iyY+wxKjE+O/qg
DU11gzBBpq93JpHd3NStOcRTGMT05/0eOCqpXR9NxSQW15XEDIhrsM6/qjKsMmziEiO7bu8EznGJ
Ewb2Bi6V9G2oqbCk4ECWIg5stfnWge1+gZzpzpU2ioly0Wd+redsVVSRb0zmCsQ7+PGF5bAiWL/e
ojcJVf+x/XTKDA72o1Rf8DCF05NEJHfU3eke3bIAK2/DOciXMDq6n3xFjYNm4mjMlsgOwfINNoC2
/b9nBfPhE2hxHwhomMHzo6RobxszRxjeeUTaDf7L/xG58XmxkQTpqqafDDfCJwwqvX8dKDMeb77f
t7IF7AGnPHyuPHr70LDrJOxYOj9QQckWNGHM03DjSnvJVlPCXypnTNlVN4gCXyOq5z282lcqwD1U
XOLA5ArV/uDn/CLdFIp3c9WzxU6o6b0GbYsZjjmuw1mbp1lxh30whlHX3IHyPOVSrrzO9T+rWFc8
d5aM2LaVbK+duAxDeOGKs85d67tVD3/0uBBv+m4/csAydkzYysivGAyJpuTjPlL3ZoJkbrbyW3KZ
b9bhMVxk9WxH+X/i2g2Jek+usruLOOfTMurR5NUKlhbCyDT60ReXHqM95OfWdvSbxj64wrGuxlUd
sMvDz+2qWcaAzjh6C7pVhkKdFC/CGL97SdABNbdYGfgJGBVoGFUlFAW8qmN74R9nnt/080BDOH0p
9rrouf/itcsOMHhc1MmfI1/0li5ZfP5CDXY9qubqUbbhijsuJS9wC1BjpvuUwdCVuqqiSwyCYz6G
3iDCUxevApVznxVFOzaZ7olnkDero/4R3LReKN8XLLNUTNVVIR6FaUSol4ryJVgT2YL05U9ekC8S
/S+3+wbtbn1r8iVZTmN+vWDRcipEfxPeyA56Qx+Lpf7R6CUeYSxAIaxdhV1DvY1WTdletPlHZ52x
zr3LmljsTVzLn4P5uqM3CYmYvSippEIVM+7wzCsfpAtskAJMe9IWZgYGIUYQGgyDVV0LYynk4A50
3rxh7YQ+1s4OKVSi8uBwAtH7nh/uPfQMIbFH2FYHsIsF+W1nb9jnrwuXMpEIuKQCwnICb87XgMQH
TrSo5soYIBOgl6Nwl8MzS347V4Eyp8rzPiNUKrTJl7i1sKfLMauEyL4s9aoFKhrCLgtRvdAzsiwy
15l8Es0bRt709euHiaGGgGeS2vt54UT8vaWWvpccSgwjBzp7RjCQTblaDRHdBtTnQ4WiC3mTR1Uq
Hhvybo7lqRGsjsy9Tn6BOIKS/lnKzmZhTOFyCRuRZyxmtpSYPoIDXy96NXQKd3JULDcYsYV3hUI9
ZRNp74FUzkeGFgiZvdxSTooKkX6H10zy1h6Adp38LHZLnneUEgoRy3NPsGsusOSPICofRoY0E+3f
1yzHs/NwrVNWhoToB862NPPRKtuKmeaTQI04qK+p69/JxLShBVFvFiS4nVJfrbqalMxVreM7TC/M
cwNyFVy5uOdzm4YTwnKT62agGGNIizgcLKMrcWBd1+TVPOcXsnfbfcBMxbtCJ7tlMIGFhedKZgdb
Fy4+OZlf1s0OrfbZE6oseydxiZB3t27+5REpNB9Lm6SiCQK11Q17DgoXnoqvakmWGmZn3Xpxax4k
+dBDuMGhrMkQITPYYRFMZAGWSORxqPjQjdmT2HpWrisVjnQsck2z2DzSIEFMHEwmXwAaHh132QNH
KN6AWaAL0QxHW6BU5eaTgir/lRnYht+zt3cXjs/xcgCQhaA5VHdMwE7qOHRkDZkAEnL3bvEFCGcU
JCy/ki2WSqRoBA5zS+1mrzobXRZ9v+AP2lAUQN8i1rOXvGAceYfczUta52cxOzF3OqFQ0LD9pTEF
Fd6rSrsq77CGM+n5OvALKLcnY12UGy23DcvSQxsxGb/fRTG/Tm7rHRNNrdnwhLLVYUcJvhpoLSFF
oMw04RFMWsDxIjGR9rOeN17JImgihRTJlWtQGS6GsZDKxXo+PraG428oxbDzOBd8s1oXe+l+qWSL
ifTtk/Wlgfem6bZdsB8pC+djAuLzA3CsOGdp2/S21MQ0U/cQw7FoHO4HAp0fUgXvbYUeF1WdqZGm
J1FRRHikRhN5lDLoFTEoHxyKHEXhKlzUGVH7zQlUwKmZzvXJ7ZyZp2fp+7xA5qR8L3QcpiE3eTrO
CVCtG5BLuIh8kdI9vNft/cgU2YE3jVJhaqo260NfVw3Z4T3w6d+SNNWnkBEmlvlEgNG5VV2xhWQL
tM72We6JbAwkfECotvapv96IKch4JBtFw0b2KE7TPtGxD76LrN7tz6jPvOTIDejE7iRcri/FV73R
j/aarUmnFhO9cMwXptde+MfObuq88muZMY0KsTQRv/nNxSuhahtLeRgt3LR6UryZ02k3oCYlMeL2
HDIbYByHfQQq35D/IuO2zziGAfZvkbQ7LC8Mp8mWHi2EE48lAcbpxCPnULZix77HYVyf68Mv/56W
Cj1+QkNG73vbbUMrSCDuE1Vtvp0tSBDtFbH0uZsZmM1fZkBiJCeIu4RpZjSBVhu0RTbi72fIj4jk
lhLWKjx1F/O5ScESYyj8d9Sm2PPVe20ipJBPavm7e4io+dqCIX2tKaP+Sd73ILK1ubYx3AXLb/Tv
PHD4BiIl+TeLIi8jUf5qkeVKCts5ivzX1EwSCBak1KhsGrAm/F0/pouDWnX+9xpGDo9ZjDXBJkHj
AJ4Namogcl6yAoIn/odEgOq/iaW/wIGLp136z0vd9EMS14H6s1wSZMJwLX6Sut2H6URA/5Tz6pFV
+F3CaEYHQwyystnPqoscGU9ij/1wsN19CNngpa2roatdzcYgskNasnRPmxVpoEdzRY+bIKKrLxJb
DudRQIGx+i1kP5qqSM+sfh1FkpOgK+Zbl+kjDyejaXGMjRgprdc5Y/dKtgbwmzD8uZLHdAj2L9xV
Rz0xalkhIJGUrutjz8VxVFW9DRrzJfQm95XUarprhq0SADCnaQ1ioQ/L12Rhm6vwcoT3B4ly3C3K
9fvt/qkxCTnXAewpSn8Pmr1N29FhpG5D1NcP3tgBaBineC9UC2n3OPl+u9ZjucNBSzzGlWxuZimb
N9RJRNpmq4waiKuEHPlxDqdhFHNfccCPlVCizu4rP0L/vNvShmWPHr2BidHZNjeBkC1ZG2R2ZEG7
IKhQ8nt2yHA4YqUcv6AsINLZggZe3Qr7fgP+nhLOIZNTs0js2hbVgWReZbepm86LJRmfsEDorXL3
i/OvrRNL5L21BAVWH3Ie90lJSrHai79mc50C7URvjlDa3juYjMWXzi/viojwNpGRC24oShsa6ISp
BXGKrJ8Mqeq66f1+7hSIA5bX0pQoZtvNLX7UH2RbTSF6Ob6p3bydNAmNWBJNwEecEN8S185y5mTq
ZJDLoSiH5hsMzMvXZYUtdK02u7iMIDG0c3WS1s7EIe2slfGOVTqqa3oUdZsL1mblwpY8DLYGEc4p
x8J2nIWU4uZwtac27p9egrd824nnjlTWossEPdorCOYCe7CqMBzjB1+gcbr/dpaqV8qHq9/RbGUP
mxW7Abvcb+cVeTB2FfxSbx1yKrrItGwzzCeJko3A5aOU8TgLUEbcYf5Iwq3JalkfGP/LpNtx7TL8
HDRSSuLJvGEkgGeSH+JuJor18XVRPH0EnBmuxWZL3GT9H/BFgfRaWAvW+YishVR3ZVPN+oxISGM7
i6bJInFzmAfajNghlm78X5QNSPMa5L6jszKy6D7XALpDCyBLJqERp9Xc0TEsPpJa3kBXtghgHgeT
2AKSTj0MK+67802NtRyRwWOTmd+e59smcovwAgCrdq6Pe+AZon8aLusi0TQ+i49n4gsuEdnVO7pv
K8SI6/tju6y0G2fZPKN3hI6nTjOTXRhU7BzQoXOBCKjr2AgNpKrm3JBDcy7i4TsNkknxMaJm9Ta5
9y1Bct7EHQti8h+XbvRHq92YLVUDXpAfkkwU9tF+dogz8/DktuIUnhLtXxxGaQoyEfrIh7MLDd18
mRo5zejKkpaaJg++dOgdybVX+qplCZkBFvx9mLg/umkr8If4+zGq+NX/j/mH3WMQKGHbsVdZ4UGD
479p/YE3fLeaCBG28t6dhsuLm/uum/QcmaUk6ZEEdYe4okCkQ9eskduUkkHqFLXvSVgkcC9v5D2V
sWlEmUcF/M5Vo7yiClXWKiSgtbWckhmuurs+8WVZWjtLRfowwQZ0/RoUWoGR07KtG/9JiPvDKr9z
WnZBDnGvguMb7BS4aLoHzNE6kcTBwBg58kkLOzPbJQNJf0x4DKFXvzzML85so8kyanYDk1qP9CtC
Ntk+4a6ipZvoL6cNdzLIRPbfCt8MclptSmOdr55efw8PkcD0ebt/cB/trpywGOYjwzCk93gY+AF4
NQMDxgDKvD8m85jrriwUIbofdR/+ih/hq++WpvmEhxxF0Ei3DYIkIKNpAwAqUDR7cAn6ClqMOCqO
R4+jG8lEhgqj3BFwBWh5UYTeSccCITzSMIvNSXdpSQgiIhXpek7v5dQ3R04smNOX02lDbs1xMCV1
zPrLrWVLWvvW3oEHID0wSgJ9wwSrt93llH4rbAd2LCyLRjVCC+8Vycx4F2b3NYFau+ZdjJ5de47T
8p0IAENmShBptdtMQtUcU3mtjrODb1EHlIALTYtmue1S+ec1Bcc4BGE285ZWQMyIf07KpulYlfrV
NnsuGctKv1/xca97fVoQrkDh2LLaP+aTErIlKY3NbvCTrUnvYVGGAwZdPlSGdff7wL3EA5qQta0K
cMLNtRTxQKLu12URN0N0q1WPw4sgaZqQ/BPg1mBvjG7Yv3mPbN4zLVe4xd9oj2IHjBfvz/prLakk
JqaaaKfEW82NXzky0GFF0cuvKKYpo0rYHo1T+S9v4e79qmHwffvFExTEXEJRvtMniLru3hV6PM2T
h97ZOHIbkkNhNu1AvnsxV14uWVlasR5gLU8DIodu5px/Mh5azoefWigJ82vPpHBjebgGcjPrdNWA
YVZaElWHbX9hv3CHEg9+EIivD1lXsic8aOiJcOGZrHL/4rIiNx7i/qMI98J01meV7IAjLw09Z74w
K59rrZrOLs+rWM4LxWerfydQLBNyqTlC2Yz2SOGIcxQ7bAEmQDKOrJ8tK/AuEHF7TCqcW9R5g5QT
nJPLK+KPhPSJWeVj2CMT4BIQZbX1GEfOvHMvoPBd0J36IiccFVrLofIzaBQ9B9p1MOCKndl5dtBp
9P0+WssVTmXd/NY9Sa7Z5MmP6AvzppbHkwzjwiTYUpnb8NJIA1Q6nX8Vj4WcwMPFeppPU5nnvhs4
9YVDNlFO6Av1R8+h1do3FY+KVZA0Ov1ar1cv8q30NXmMyDt04RKDou6nGgW6C1mRLDIfRM3i5X8E
peolCHCprpOG+SF5FdpxhuyxNeI25tmjg1qhVZzCp9BNX5T6LfCzRzPNI+WyFY8fzLnQjbD/hBuk
8OcYvLQD/ih9/E0KwDrr4iHCxE2BTa9bYUcXGa401V5K3k8C6tMq67X7KegPN6oPZ5H/KSHkrbml
KtZiBcxfOWFcHPVeDpEYNskuo1DzaGTns6fWGY+ryyfTMo3+nGAZsbR3hgB9bW0/z47BJZtN4a/N
9+x1IGYdfHRQ2TO6UTdcQaJb/Z0qBVzObMBjjIdFacf98uMG5Pz3WRkpaTEJdbZ6+/vib+MN6cmj
x56X1Ch4FtHKUYG8e2wRoccJFIhc7yfNcm1g2N93/wO/B4pY/5nj0C20IOZndtl1/orgI6OEUp+a
WrO3iiY5KQ7pwpEw1Q/AXqvTbv+VOcBVAELbITNNTzWKBiOqe5KxCXgtEDvHuNcK2eM9EF4wEiYU
D+4Z6pHi9VfgDWoca8aTuG9CtAlMAA6Hb2YhiWRCCFKzZNpb0X6OFyx6gSp9K/B0KBcyZTxcH3jQ
fHwz0vJckFF5QgtP2V6Yg8X8qTC6NMv+5hMvYiYll/WVdhvAGQZNEMGQMFOu0tEBu7+2Vg1bYKtp
zH/mijW7K4HZ6h9M8gsdnZB60EHm9YVDpbxzlDhSGzWaBPrCwPr2JviuR0LmVlYuQa4sch9TYRjO
3NVTKoP9R+aDNIx6kJTwrEkv6bwXNf+B62KcD+KsikhFEhPyQnfqBXr2bkrA3H0Y0/8vVgBvEK+r
LrdHOYP/znVX1sBS7gyLuptz5aQmI/HbF2drKhO7G8VWCPlQSlsVpHcwokU79HKAvo88MKRi3FnE
28EhtcmOioqHHdimIsMBEcldA3vX6DpyPzbdcRU6VyOlulnsiY+qsMJGUikIbXECTOhW+Z0UjMHh
q4eOQrvUIbWRvG2cGI/0hYiN38TKy9ljOg/ePrbVKcPPpwrnPFLZc/UI/3lqBnnCTnPAl2auUnt1
YyJHH4QDR/rD8r6GAKmthfWYpFzK3424DjHmIxKdfmD3fYeyQ++RjW4PQwEo7WZtog2KBsQMu2em
JqxlFg8/DAHxn4tio0IUJy3tjWNmMfOL8yNYOZHKgdfESb0OPbM3xZS4nPU72pLGDCDjaWSvkOYu
o4M22uSQjmlBgawgddUA8v4OVB0yF4afLO+KuVmurU4U7T0QIGGc7WVm7whBm+Cb4ZtCUZK5nUPx
pgCpkuCe9Rvr+9Nn6vbKyyN1EcV+Ftd4AACZDbKaN3ruvvDWLNVLk/ZBSmi/Oe0IAnE8fYIDUwsI
mUdHLtb7BdR8na1XMJIoJ9fkYsQtJ/K/ctprX4xoQPQZPcEyaGfi3MYyVevtRDI/09P7i9coBZVq
ZRau3TqFHz/pmQYH52RzL9hNi9APog8z+Ju8oLSXX+JiyUGlIEXBm+piXpRb4hqSUfAkwV/HdBlW
Z8WqcLO3l/uP9ON+p46O6zj1bMicDgphzSqgasMM4P4ynXK+/2CJvR7pIKmKZrCgwRIWOn1QYKHR
cPI0O8eSmq/p1wmWCVMbmga95GMXxloFCHWKMja40ZnShspzSTsBfd84+M1XuJAM/FQDI4MJsIK6
/QmjpPw9UGz7+oY1NkKcoxjpfKUUlTpVUuz0kS3zCR4geKwbItsugUinDeVSzqYbXpQv1xQPR6RE
tKaSbXJzcKHAZz7136Z0PNnpRSUOlT+ZPLOY15T2rzf+PyR518YWX9lX1CJlo3fkSiWpLQEkx2FS
gEAx7IAo3sIA6mRZiPYjlzonCpxg3THwcVqDFr5YyepjPie9vKdSCaNcyLHRqhjRVtzfTLYFmCeH
Gz/rAJFNgWwO0mYlwkUqKQ0H2AkuMj3svFvnIvhtdWxz47vwx07QHDgtBz9R9k3PpAk/OS2JOQus
2Ll/ZwiUN56yDT9udkiSdUjssVsRabfpMEuxgDEoGDdnYTQMotEas0hFaqWRYEavxBrMdosrc/Dr
JSEBR10EgaoYZt50orEW+VPrXMFc1PQnSoCkv6jg7Rkb0D7/HvF2HWPvahQKIigHIoVptyYcgMy4
vPx9zSnFrvntLu7mqDCwXO6zjDpdiaykOYmc429QgzkLurvoCiwvReBHE0yto/4Ti70j7m9MED8z
OEqU6Ba9e0fbtoZYj0Ro6BVZlnfK8psEoqo0IdeXcruHx4XOCX/5AKRF3HwY7/MnMvvZwMnB6Abd
mH78iSHmL/yQLC3FaFufVpxuewJe3sytFp4/fcUjUXKnvU2CA7Yyq5yP+rfJeaIkAH1uR7U1q4Wd
A0UW3r/3Qbdqv/QLx9ySd7xr8WjrlE7La+LUtag5ibujhXLe3aYgycMLCMH3vAuev+nCuFvF+/jf
qR87fIUUp+K8ti0ompmY0PM/ZvsvM9hXl8vYrJ02ZI0j4a4tAvAyRPKV+E/Cj1EsgerTAJD7V7ed
9dGaTfO7VrD91kv0tHt+WwU107ANFW8bx0ox7QL0J/5Q+0EsnI5JqCVEbLm8HjlP6WFJ96JdZoMm
c/HDa5Mhdsj/E07akhJa6q6bLu0kGXYzYUiHvSrDFfMHhCl/eRIctfbbGyaxCtm0JRNW7k47xDDl
hM2Ov8C+MZAy3xoare8DI6CJgUvOh7qmeElUbwVKDEzuqnk5vFQ8QvEgBOONNxlQRVy6mmgqIxMW
/rztoS0vki8XOEh+YTU+sbY1iOv5m6dI08QoOMBz5duZ9ruZC9GTpuBH8kXKi/09Pxe9SjqM+O8s
XkaxMblzW8JpSw7aVkBBDGyxJvSZebI/agUug6jMIpyRj5CF9+gBrjS5xOshwOlW5RIYbJytS0cD
QDs7UQZn/hWhlUdTz9Zyqe26CEMFcuhE/FyRjgrBRc66ElcJ2TiZLRTJDX6xNjC6FOChZmKWuDXW
Hp6tU70uky+nw6019tIwq9vIx3AZa03B3tNtFFwsaHXZ5N3Nm8BreyAYtfSZcFdcLst7IQmks2iD
koP2Qit/Ben8H/oXJroc6/BB7CywNMkGYCyaBGQ5Q+mG9/qx1gubXdnWRu3iIV8AtEtQ23KYgmxx
TSvILU6fsj9rXrmJSPlDXZiIzNkced8AzKqm7+trC7jHT8FamCKiStTE6EQOvFo4P8RfpJEUP5vi
pqIVzfuz6/8/7xuc/GaKeDIFi5wOyFSJfHT3MoXPiPtC1dRxU6Ngp7VF2CtJr7G/zHkTkOiq7Xev
+rQ7asEvMFwCoLEhEGwv2etupFpH4aSr/hY611kfT4f6BaFHGji22p4wEz1VkmUteLYJ7aRRYpGz
S6HX5ysCogLwkPlBc2NUg8ZkAjLXT8p9sIQqGFWl2OStOnzJB2ye7iRyKt8DbBNUeLJJ2PGzf68t
761Qb9bgiOglGmo1vbFWxLshbkyXgCRX4ov8PM9jeIG9eh+aoYJBFLjE6o99ibCrfn+LyBep/ooh
mxi70MPThdHKHHQj/Q1uJH0FOEsXC1sIrXUtE/ALDsNv1o+dqXbNEoEEU2SNFhyaYjf+nbUEyC7B
Wn14J0vK1yDPPxZPHdejjJ6WW8Qfv0ZvC4hatTx6kIaToJGQ5VGFVw2PZtnhF9S8r5tYi87Cz5+l
eAm+VBcA9js8HxVxUlPkaKUEbwgZuZpWHakXQVy95uKDwrY6CIvfqbGbHzPUQLo9UXmET4BLzO0X
8rIxXZkSvYUToDXLg4LJx+AWXFrwvI41Nh9eqX3jYI35EsXfj20fXu5pMleWj0JlkUg7LSffa/JE
SbMuLe7MyCfKIwDA4LUMDMKBIphzktwEuI7HzBIsQiItZkZHnVyQCOxfFwnc7XEHdPmTfT0JSoDC
5EpY+SardxoxUP5+gcEQVVt8ioP1NYj6GRjTb2DArw8UjZi+TxVJaoJyrhme0A5cSaVECcysjVT0
KjG4N/cD9UPXe518vP8WfGOhUsJDQoNXP/w+1s6s74lcFaeLroNwt68pFhelY+iew5nxUUh3tGuA
OGultNZryWi7G62kEu5OANNfzd1wGs8NS6z0prPMetSeMiE1zBhZ2TBUfwMLwH5pV7dyCKLK69c/
T8xPe7YooL3jMl450IRvic05eSdNUql2oVX04ZJppx5nPw6yo9xrls4bxJYC3e/D9N8HC85O6crf
NP+grS+9XiPtXpBZN4GnJ+WRP71Qzesw3j/KYfK/nBtGP8oJAa6uhLHodFHkqNNLIvNa82mOI5cb
T2Ff+2ZBU5giuu7GPBPXNnVnwH7sXaoKI34wxEXI9lTRWR51MKkuqmMHsW0rjb98cWaaapiLHy8L
6NtrXFEu7pVzkYwv4N3Td6oG0t6PaCEjzaLgoOqf2A4MSG4vy2idz3DmdnlZMZ373XpHPYIWuss4
8M5fv5P2+5I9kB2IG/8e/sDLKUvQWP82fvvC1zro5boZjNeV4A1KaF/mwwG9CRJWsj7qLvf2v9GN
UM9vekFvp4FJLYkVD964vsUX1gvyhabLKnQFsJLz0F3l5FIj71h28rXIKSSL/44Sw97NZ2ehfQE7
N/xEUBeZ7UthWo7wGgICavJ8+1Ma8aNkuuDEuit830qelv2ftHjUpLo+BOXPm5Ax8OtCEqpVK+dm
gSN3lsiOUWJItndAzr4zre72SfhzwZpUET7GMQ5GRL+ii+E8vVG49Dra0fLexjBNQiLXCdaCRqVP
lIIW35ukPti7HNaRZuEiraZwcAHR/Zc46rSG/T+rjh9VCxROlJQklgoogkm1zAITAnygVpeRjK0N
vhEULqTf33AP3QLJSLaG5wTvlvOPPVKcwtEPJudPijNPRZkC3Mtmg6h3gadPkwZhwT0/IOdfd5gc
VUjJrQ8PjECSNwBkUDcOqHdrSMx1AzM/AskSNuDZGcKqaQkGBTVElG5tn6g3OgIOYdngjx5uBw0x
P3zcUwNVECaAbeOVCxis1Nl1Wlv9+J2lN6AN0eZxQlta0oeu7w2zBUobw8xZuJXniW1zBFcGZP2Z
tFFHHU6QIcxKfKqpppCd5584vvRVmVw7X3FF77PPuDfTPxfqRW0q3YltvJQqls6GmufCTsr/hH/z
0pvQrV9EL3nrAYUFkXsFVKKhsPQx0NLJx+3XlaoKZzY5mGUUUgziyZ00FfTd58HVfj+nQ4bG3SFp
O7uMbFymlPlIvx4ix6ipu9P7oVlbzmAfK7Y6eUnlkzltBsyVMldZdyusfijMQeEFX/1jiRrk0d0r
yEEgv1ZHeE1sueMS9zRDHWCKzisv6kucUFzpmwvjk1dxeTybXXRnOz2cZv/DlekcOzaq19L2aBqb
LNtzXC0mBO3ZaI8dJ17KT08eBKw8XVn5e8k6TAcjsvVNICZvNnNa5+/SaHRMVi4yq0JhOPlUXEhm
eSlSe0dHhtdVu4w+KYIQOu97jRAuxJ7v3yw4K66I3s7ZKhwQOGG3TkAKbBxMSDrtkR+ypqI6jnf7
tXk9Pf0oVbqzFuCOWMdDx+/ICRJVtDpxMdHTIZWGTdE6pLGUFZYB4Jgg0y7zQxsgDLieqPMzgq4h
i0hD2SPue++dJc0XitdOjqFad/17ki6eWqpbtvmfrr3vSu6VZgzi6BQOyKqgqyf+x2whn+0hUCbN
wINIPaHO0/vzWfdK0TQgimPydm/QSK/nySOrzNYz0U5r9l2l/3rn10X5b2+lET+kJkRObuQGERHT
430Vas2TvwTBy14eQR+6Iji7v5SqHNH4ReoEVgsT4ZkKtspLeLBtqtWhyO4+vbigWwwkD+xsm9DG
NwXaJxxgllPtFzgj65/ngGHGkoNSOF9JK+uahdnqneXrn7kFtNioOD8DX0RcM1xUx2xtXVbL6wnG
d2ipKol+0EbGh0OLYibBGgT1trOeR792qFzP3nowiiS468LyzstZkqMQ1toBOi5QVZ0Hl+v7cm8M
fg3kMT20YSRKgO/ik63+wwkgrdxp1hmPMV0JzuBjzbGeEl0+IpzMPl6r05iEHoGHPKGe6zUQ/cUk
Dc3xjW9rHUuppY/ZoKXzg5PKhHdPtN9pH7ngl3wDmi6HiY3m140tSHd1YGzNnru+AXq/m2q898Gx
82Q6XzutNcQCDCdhRvGxJphUYlCwV+J/VN2KggHzC7tcwynxkKU2ZQMks5AERVLvsBxJaPltCzil
rLwjChlm3hGNFp/bpn8Xl3aFurdHGPWljjdbQLTywaP4wGbrClfCSOBEHL8/SjqSCXiTHjwQWw0U
6bh0iA4YdympJ2sz/bRSw9Wxn7RL/GrOc2eisk19krrC4nRcD5zzRazSF3x5apdorxuEeaLoxKTt
K2L2egW5+wQ58vSxNd+S3t/eaInsJHlyf8LzfD+9+fNcTg2qTIbgrWgI5Qweht9IzZ9KWVJR1Cxk
5lHeC1x4MFfHGNy4gQfdFEnAYOPnOnEBUFBjw8U78xMCgh0SUY+4P+yDgk46nYf9jj+e1rT4t8r7
OpRR3ERWzXAY3sU3ZqN4Sfo6c0n6+DfCCyX4idxcVE3k7+AJTBRjY5Eke0FmnmIPxyMXFF/0VN0i
C7aW6QcMvFYI3Aqc5TcbPLokSb60Vu4IH1y7FwI0vAvWWvYkwq23OKWdQzdwuNnYThsXQAhhiIhL
LacrpeOkSVYb/fFByfgGiMdJHobp6hvgNBbzVArnc8LWKYU0CkT3ym4halBfRqPDlFCfxIDwA9V+
4dBRLmfXMPbOdR7XRd74sN0Nf7ZcyW3XUFls/PaJOx7QNqmaP8pnhy9m59rHid7WC0u2aMfz3grz
hxq4b6H+AQ98td7YoEWs55bSILAXdu6ySt5tdqM21D7UZt6pgKVJQYirEUFDpWpON8FABaS1voHN
f4an6GH+N9ZQ+nVmQzMufWKbhzHET0CNAHajGxTO9p750ORDy3KekzF1gJ0j/mRWdJWv/RIheUBk
68PXl1j/ZcJn/W07CxyJc/rPGeG9m5b14na2hnikkjQHCEdSk+BcxVcJFUlkxa4MvVNre8G+0fZ2
8MYDnatxAePcqPNSPVnE0mUiCDU3hc4v/24Tb5HJ4ep2xnUeZmxUwY3Gc0D3YDeEPFfm/YlI8z6q
O2S1WV0cyihQG9lc59vPrzR1Me8fJ1/nJ4oA0CW5nLm2HRy5GgLLMVXLeKe6EXXmE9LsT10Au+kR
41ZJe2g53DCEtIxAFpem6c1bjRJ9rdIDoihVsHUHm2O+Q1kGDBSm4gDjcvDBWxtsDlmzjzcWfdFs
+p7RIairj9KrNy7/C/FHyuLDZjNb18YvC7XfUz/dJYTNTMPJ1at8MN92Y+PjSYGZmJw/7XcnfSmh
PGJHzxME/2RFdo6KPzLCcF+LEnPdKE+TpFpltyXuxPV8t/kWUhwkOaLOcoO5Prg1q7uTJG9HJQJG
D7wB7OzHZkiFJs1yl2HDIkTUfxRoDKAvwE9b47FoflcggThCD9sXaPIOPXh94550GR1ldWBtt0Fk
XJ/tJkCUIHVWGigh+SVIMdxQ4mJVfHqd+SDnGKY/+/OxrDqBvvTL8e7Ymla/ak559NsIKvhu99nB
tzr3OHpH6Zw1PUMkQdxMcR3DLpQ1Ayxr22aLoWsBaYyrdLVstiderlzfbtz1xvAeO4EVdYIdN4Ll
Jffy/htdiGc/RSQC3vzD2hKlKmnU1j6iWLagU6Ij7n97qtIm82yHFD7NLjZUTejX4p5z+lP46r9y
o3oPqyvVMWeNeXYXxTLxJ2dLr/SXkhk0PffB8j2FQVr6B4+tOGAh6H9I0nWU2hUuaiWNpDIj1/kf
hdMWvtY3YAtcLcAtPNk5nFsbzofgjNEPTVK5Deq4Qh/yq74JuGmNMFqSINC5nrx37aIehg3Sv2Lx
R66mbfgpwreiFeuCw608CdM1kYm9epMw0YhBBqz/et5nTTQljL7njXH12cD7ZknzHh8SAtelmQ+P
p7asjO84xdJjCcQ2D87oQRwrbyMBr6we3tFnEiIo5q1dY+WapCj+cU9ErJYcRKbuQbPyfpEC9rPu
JsA1erExryNgdzmyFARD5w0g/g8SAlSgiA1FPN4VJrdcM/JrgQD8z1rkZjzyL6G5XKMDQkLKWx5f
hfFZgfpXw0fhKl227a0CoGLLKFjVE44Uj66kfTRlKeYF7p6PpQ6QL4f8UGk/l6BbkeBPHOl6JaoL
6jYnz6pEq9FRmImoVbafYV5ZsiEVJUe/4LZkqPumIXHVvGzMefNNsmg4YMG9E0RbU4t8BS5HsnQ5
vpHctYpUkzWBLIrZ6bJG3TMDAHb2/Jx+JnspGKaEJMqCGmhCd6GLpIhnNiyWEO6yz7rmZOPjEobd
CoEerwdbNmNkji2SZOXez6hKN+rFqcaDbAFrZSj26rgtJuZ9vGMfky/7P9tzI8EsmbS9T7TyGn3O
fuotMZ6tAnfrt0Rz2ncd1QUKnJqM5FxNvOBLH00JWG9RNC1pqVLxC4JGZN8tn7CJZ9AoQTzIvIbL
oPdHGUPTVRNzsEifyX8xwcV4JmtZSx5jqGefY4quJo0BHEKPrOic8/OAxSj2A0RdaaTzDpBVyL2X
sEusoHctC1guqnvfQVWr0wLbNVnGbQrOOr7cm66JfFy3JxdoXiWufTnYKflc4UVw0IKMZfVBL+tm
FdbcDLBe55pR0+JlTIDzxLT9+5ZqdpVtp4x6u07bCDZpIJfctPyJ9k/uH3TSLiD6+SKuYNRYgIBI
ZzvxYRhPJ4vbAz3CoW4UemJgvZoyJgk351iOBv1ZSp9noDdRIaR0ksLNgbRxVyKdS1Kz2Xt91KXs
rydWK4vmnGRZ7mo2QunHeLl6g1zKLI9U6LDFCKAUfXQvi+0MkT4H8baYJBHeZAC2IqYhNjckOjmG
d9ytbas70pOUVJ8tdR49y0x2igveijbBxa4V4Ut8fLXKyj9VuIBSHauPjoIPAAfwsguewdWYSxAZ
wwFcDU3phw9i/bXKXzDpP6ojX/qnAi3IZInANlvxtfVUpfiRLAOq4b2CP3yXeow2CqE7XDHtQHM3
jxmNKzLVZQUm4cnQCIy9SYNusLqTAKrtfQVhZxVmAp+42bxkBsSUqLMXj30vNigc9b/UKwGECHj0
jJZUvvynOkhpj+6E0L+q2hggfmKNbLpiHGtbbyZaEVLdbI47RGO5KXtv8zvZhKBPTVrbe9kZRHQB
Hf0uuqjpE8kg0fLXeo03BKcDVZegaWakz08+Nr+rTb0yeZ5ocvpX9eTau3z9B9jDjU2DAIlXwdv8
qiRMsetvLmilpNNMU7UJ7yWgGLxIC50+hRNZEO8nGtsiau5LOrHwiRz7efGYlOkvm5B6a1KGCy4t
8+tefwCoRBuo8W50cuT0zu9IvO/i7y++0iOHnrbJ9FalJY8gnqO0RGy/z3X0N0Q0ZbJahUZbzvtW
O1vdeZ1bBgouqXpAaOXH/12FXzWCRrqkz4o9FVFUZCGnTwdzG+M61kv7RW6VSFoV0IUhzGOfzULZ
xmJr+NUm1IB06yD+KncMFkAStSFNSt7O6zJQzEKw1ktZ9xRN4PIpifGfBmNNPUQYP/JUng2Twkr5
oVXKy2uLnXgwLYZtTY+HE9/s+86AunkmRe/yTnwHLg6iFTQhDjdis0M6L2TGW4tocZ8j6KEC8KeV
Z0kx/uxFQyPyKsFKw3+kc71B943quoZ/wDa6gS2s8wd1EFZXQ19ipjG7G/+58fkVgSHinJ+UGqxQ
Do3g1nmcS1oQ+jg67SkeyCyWPUAg3CoFjal5DtlbRSjJwDEZqcMihZfApTQ+4O+InPHhAqQgznwm
AXwr9uZbufG2HI3OuhDj22fpL6qy83vCehuPsLh5gEzCym8iopl6pWkIwBusUP/S/xpG2W5R2zHE
xV9I6ddBuAuJn/ti0oVC07Xy6V+OIIM9p4Yx6MAeaFL/73o8XnXCX5rUsq/xBe4+y33zdw9nAh90
HB9fqCoKnNIUPP1lYMxifJvMkS+F157bAR63Z7WefnVV/Ls4cf6zcy+iu/lT2xz4dAHa7kFs7wn/
hyByIcAe47VJvoZ4Y0aR14NKvbl0RlrKhwAuOSQMfeYU2XHKyuGRx2Gi/XRQLHIUO9CfWqPAFVBY
VyD4p2RIO6rQkWF1T2JOELlqRrELarRGtAd0XppQ7L9WmAcX0+12NxtJfV4IInRvq3/Q5bDZN0cK
fX3AjwbPk/6jDEYuVT/A7xhnpL833CdnX0MrTmWIulnYg7ODlt6qPjmRQVeKnXGboe3zZLavnbL0
MacDfNmWf1GXpd8k/MmYUTyHnWn7RuJ7/aWV4VOnMxK6uiiLpTgWCxaPoNOEcZ5Gb8bqDgXrzOYL
J7m5HKK41wWUelyya+G4RhALT9wt/NK1YoZFvwCDoyHiaF6I5UhLelJss6jE5rIDkLryLE8wpQSj
Hr0KkCj2bRbfRU9BuZ2wtnogk54616G3K9frMZ8Bz6DR4j08y75O9kbuajrQlYKpdLj+Kbcsd1rV
Uja2kggsdIGAtC7qP/Q28FStwcdLV4jolJsHWK1ZFIZqUj8hKdlzRe6J80jv3RFfnPsVvR9xYKlY
RlWJRLc/79Ezzwk5R2Uwuo5Q4Kb5Zv2Snz2CD+oMPNiojDBuvEsT/7L0XK+UIYX72ssJ1JmjYWyv
rUNGGyc1Q3/JrJ//jIfXpcKWnj20QXPXFvUn2XvCkEQMDCGwfb4tcPAxnsrHWo6al1isCKvyHcbq
0VDFc3BjdkfDHw+kpuuQ9GzM9d4VQs+3PGBDsJ/vy5Kh148MfvbVwaieE2qKbRgfkx92RjpGcgXx
xJAe/l4vdkjV6hw3mWzR1avPQU7KEJmu6LwYONDkfmeUSwCmxybMcnM3dD1PmTX8vBW3QMrHKMSA
C/mKLGfxS6pRsvLhRA7oxB7Oxxl0OVF57dwLt0n2JEA7l4iQ0cwC7dM3eNJ9bTgZpS1/E+wpTqdy
0NEiS7S639GoNVhAglQ3hrWJPtvCszUNKPHPXCzjy1A50v2CkQGfcrAVySzbT3CrH6CQEtSwRfl5
v32EYc7SPQT3C66ZPhhmwmBLoThb/N8mpgLOgn5j++zUCcDWrcYgko+cWP4cUERyiWmZEwYYTnWH
6rzhY52SQJIn6tCCjMqdmYAnOxYtTPK+CScr3rgAZfEbRG22Ln2s8+WXv0s3oYnZY8sR1JaRzX1A
x+l3yt9uBk4WpdC2zEsOJf+wopmkupLEnpk9X9+jGGbYodFgMP3A9lU0NSFLMOZPkDnjB5aJdcdH
1XXfOe1gAx2QGKy0KBncropoalHb7VNhYKbqVJsxLRLQoEZYKCx3RKd/IwrWP9vOR209cLQYGyb4
U6sbZfu4XvOzseVizAr93xxAR5kUI480SZWqbAmoUjZOAhrX45/RIiw/JwiVI+i8siM0Y+l0xeXq
e7qM/zdlvJFM1AjFBE0Des+iJ1BVTpZD/rtQ1veHhSxDucZ730iVq7rYAzHxBVz/zh/ugB6oPyBL
HwsJGwn6E4UGDObMyeyt6n6Kfl+z9ga5hG39D6XowmlVb/9hh0BpMNhegNKWMBsKcsuwbZeYAr9Y
Kwa3+YuYzPeQdHN3XiEmwpZxPQCDk6JPtxt/eby2oFrfkD7EX8kwubano9q7S7gbOwDFAAU7UY6s
83UNId2B464FoqdKRtDJI0YCT7N6KWjFXOrZ18NEkkD/RMRem2t6ksirByPFeQDEx3kfG5uAfcnH
lfdfx4unX0S8nTQgB1WyjTaX0rlpVE4LWMMgC/fqzYEbmWq0uoYw1vTLND/AxvuOhYFHPRc42o9a
3eOc4SGkwSYyJi3R04+aRE2rvhDtgasUAaHTY3D7cMFARvOOTxJQF1vaLQtsXbNgB5Ke8/ve8qhk
rLjqWsNeMWr6+g+EnYWMelvVKhJXHLtDYj33W7GOkove1g1oE7+GZiWPMxWgsXkZW0UQgAWIF7AI
b0pNw3Z+wWyzTKT6patJm0hF2EESvcARWyU4VnLTbTxJq94y6Xt9TYeGed4cLShuGSb7yg5SskhV
ocAyTTCChtHabWudD4EwS6sMwnxHIHrDidYC/88lFVZzYQiP5KsLTJeWNp5sLw8rrRPaw8pbl6CK
udmdTBnmfzl1hBj5MW5yjvL/pgDNvYR+Durq9mBLLxYrX/GU5ieLomLoj+3pHYVoq/Z9R4cAAkDU
mLLv2FuV2zl5gisF3NKMBg+GPlxD9rn9+BnxrayWp9dSBQqncEbrjAUfL59gJApZrM7MD4UijYA7
dJd1GRm5TpihpCapcymx5XvcnfYlx2hjHpSqnHKpl/ka2WJ/MIcOpdSCoGOKHWJPkya7AvtqbXPj
ohta5AVMbiEq5B4Wso9Ubt7PBPr8raZ/4B+73FId/Tm47o1LYTgZdZrBqZTA2E8ctxA7x2037ltZ
Z8T17Mv7rFMfZ6t04HnyNq7WujRRE1e9XlPfD4SEmsBgVJTMI7PCoK5kGYmSr7aXJVVwbUd991QG
W2IncRdc5DXZVxY43qpBx54QEaYdQtNjrCygTIF7epNW+/7JkoVvY/wl4sjnAN5EpiESqtBgw5Za
earbOkqshZEjWue3rrhbrXip8WnBZo5hBsfdsY8BcjoxCF0D3KKluG+p9GLBOmiBjZJ3O4Hl9jer
k08vinOJhEohtC5FfJg53R8jjWrbSZEfuFiH1Bvy2BNg4dB6Twa0N7lj5pKpRjCx08d4wwMvmKPO
THHOlEQxKs3maWNnwGfcuHgqwpkk70Dy8DAT4EpI6P/apalyh/iOIYhWZJ9dlOmQ7SZ21Q+jCGG7
MQE3bb/yKORcCXJIA1uNdXEhOlPBIhFIZp9we4ffX19xvMDEHMlR+GebTgvT8EJQrBd7+JgOMsaI
HrU2/BoCI41fjA/qnEQM422CPAD8a3P95RjQ6XBppX6qDrsqPdExmfR3VNkDtUqYq00Y0Fe6hEh4
RssJ28N/3HzuyOFom6rBL6Mus224dbuqCjMfLixu8/sR2rPO9e38BRWZJCStPmnAel/RlgDx7VrH
sQM9omY8i+bkW2LB0PsJ+fb/g1wzNtAJq+RKdTBIe12fqSNH/F2RYZ3QuFFAm7+h3bC3Dkd09iQ9
OHtUyunAz9yZ0tW9G9wVwO3jStyslRfP9YvORB0fv/WC+i36qWb8wJY8pfolrre5vIZLBhe7rTMk
MuDSe9raOmxrQ+lNXwlj5sd3++7Z28DSheTq0Gc5Z8WdRM7djXRv/WyNJJaIxL6isbZUtLuJZHOM
Qjk5PU9zxaReNmNdBC8QBn7aZeoOpEkR1GOcX2SJrl4frvz5zlE0S0jvPjb7x07aCctaqPOKM2Cg
xOUMG21nXGYlmlfdeXUXdEbyuuk5SJHwRyB2EMM1XlqeD1who2dthAoCBojplmnUBNU0cRLLCZde
yPbQt4ckuh7JXdklCb5dx39h0BYUK6SE5vlJcxyYvTOJRr+QQ48Tcarrqs6T/nLFu5arJI0VgJfb
rP331VIuKf9/i4rTGJ77ujD60J4RhASHH0k1ZiVveKiKs6Flm2GQ+uyx7l1orXwyGpBiWiY2dB1l
PAFIjC29vMT0k+fi+tv/yZhgKCRxgq5T2sSE+gC2eMWVgCjZa641jO4LmCgJjmDZKa5ft52VD+QQ
ilhuJWt8EwHHQsVTOBqOhRr09bpfAQPV290OnzB0dw7qMuxpPcdkRdX0zy7L95KbLNQz1CWWbADa
aCyj2Ar4r2KdEkPhd0qYScsjceAZXHYJxcmBmh5DVH2AbLaiAJ9uFubk68I5BrMfYmhPZo6qImCI
UnjtcZy3rCWhD5G3HzaCmpmvYshIXjXP6+h8GKTupf8FbxZm3FnYzi2i3dBaSZP942T6STrm6FXx
sw9vcHSYiZt4bHTA5ccNIRhilTri0gXWSWrq+/8bhwDlqhWmz5Tz9h7Owzeo1mpFkRSDJzbo5sNH
ZwI2klWhpiI/GpMCQ5SN0zMLfyBLZhHtSAzeF8sURsOw+ZFffyZ2EWlVvxq3Aq/Cj6uxu+OiZOey
GZmZx5HTsRDS6LTCrBPiCjP5DzHgwBF1+V4UnqxPQDXqLA7xW/en6jT+FfQPIXqUxRP1vGnMZrUk
Bw534I66UPbEwBTscsZOnmtJUDIHASHkHJJ4O2NasecxUfjte/eUyL2/RtcC3kI/ZspcA/o1nwiY
xl1q/z5RR48N+GpBbxMQOnR2tsHZ76l4LRLD/3n0SfgYc1hBbGXZk8mfn0aCOLXHKY+9B7xBACb8
6B9LVBWTGgPfMwUX9ja0z1NZVEwfwPKxd6RIXyPPGaIxx2VMBZrQMJDCm4zdbQBqH0e4YrmRKe9N
T7JvHfLTUSd2yXlvUgqFiO7WTBVCR2CXfF4xMZ3kHrYCZ7TCabfX2+IZ6QZYjtEC+c9Eu0WzFddi
D1KBfsuxTGSXF9w0+99DDYIJpj1eZtQuNW4rNFntCmXCgrgoW5R6S4ysAg4sdVQZY4LAeS6nHzW5
eYDZdXsEQuTpVVZX1lhXHo3rj7eUf9VvmpCFr3t6Znx7x8Cts+VQQGq1Dy43gqfPm5QNn42X7vcE
2yPVfm+a12tDD+UEtBZ7xhQb2HWm0QkZBCvOU72zJ4HCjfIkOnvw3xLV8CKu2aAb5mDhSkmxpJ4A
fDbn0MwPHxGx6m+LbX8UX7LLJVus3h4LPmmaq+DRoyRhkCXeAHVF6/PD6QYo44qkSXWOGRp9ZlIK
ainfz5HIt/T7o/w6APkcEsmCcABiusi9BIKDjL5jQLj9aoixr6D5HtQWhy93lbJ8B+c1i6ejLbmE
VtcYCR+8PicqoojwmLSG219kO6Gd4HBVcfgdJy5FM4QibFX8TEyE3i+wdxAZyKxqJ2fao+NzwxOr
8cp2JCdN94Po6Jfe4ph2aUXINUdh1QFcIgVrBXuLa4Es9x3DOrelXjGIyNKdHpbGe5YbNPSOR0B2
yPZ58sPOoTJir35RnW9wkrggGWZSvuxAzMLf3M6HeAkRnazAOk6zSEGY1blh9e7nfbccpZ/DbwAt
rufW67Dk0vxc1zUC9y/GROFFpwMR2XHLXR1LxpYrFmzb4e4U8OajwygfZf10JN5JzOyLqTz/BRhU
ZaSZXWzv12+aUgoY+nrPsjeNNCBZYB8vEWGwl3CnRCXBYUwYk5U75Zocehe9opwYU6ALFmEurtOx
tRf1YsBUCOouWBp1Cg7n/nIEd9itaQIWtiEqnnhrHj8+Ok5wmy3ciuh4fbJa8A9jHnOiwaQdRoMn
CXvM2J4KleQ0ou6lotSpOw+o8wpcOVQrxCFM9zhCkni+dhUb3T98DFXYjgm9yu5oze4GHLP29Fx9
r79zb5nEF1Gx6gSnETKUmY8VEpTNe7mO5yQ/Vws2PKzaxKAdoGzqBrbuMyXY3bEo8dPaFW3uEoS9
pRwwOfYMyfNknRNaZrnPJ+mdFn4p65AB3QEhsBoKmL9LwASTcZ5yM5MX6vnC/Q/NDKJY6u5QtU5N
WjsVEj25SUy++RisCX9OXhhHAy41pH9XEujOSMUzQPgnRrhTvEeYoTkcsUnePMF45usMCmytmwHu
MQsnq5yfgqQDfpl2IHhIbpdKG3SI+wuizd4YyMePVivCBLZ9aCWCYByx3f2tg5zwF0pkvNCwxR48
PM58hBkicU7qY3g5qVJBiX37Bnw1KIKoGTkoKKUnN7HonmkaTQijh9rE+MypJagxv+hxGVombaUD
QTKK70eHuLp7Q5Wis1JTeaOnrX6cah2iIYjXNQqKFlNS7gwvkezdtqAGeAEZ7TIeeQ4Exe0ZbKSN
TT/V++q70t0EnaBrUCIBpwa1/WO7ztTZExfOqEOqz0AlDehqv3W988JlM9ph4SpcfCcsdzeXNCvo
Oh877JTHWOdPgh7Tq2myIh2NA3JRr52uhvZQ/YhzZ7fLsJa2WQz4YKyx44vA8Vc6x61f9d7qxB0R
AmSgDh5y8vNBNjizAe3LpIXTorYjFu1RYV/43qWyaniEBz1qV7KrZcsbByXwnkDLbKoGfr3eMRVY
DDgCuC2A9+hS53Jhrf3Mobxs/4S4/J4xykagPqJo/Osn3FATC4LzYYqUgzoRGJTW/g3bP91hADJt
4Kaugr5sA7MIdzcCMC9EQdzjGvDJebsE4rDV03ng4D6xgzLmLAspz1pyoxvhoNLbeHznRMsfwQXz
8gxLrctXTsRgWfBg8ZPagD7kccRYJpxvZJPYtq7JwFszjbZr/YFKl/aK5MwT2yNMxZ2NVCCZFYSY
42njaV23h6QMXCq8iRFy/FA5rJ+SX5ZRaX2glzgS8hzFOt6Xv7VXM99hFpMBcQpssUxg/8P8fHVd
i06XgdiqJVZgvFpv04Rgf1mR0MEkULQt0DBB/wcrmyDRkNKJCallhrCrMV7IZUQ0j2IJb/6WP3uY
xgoO3q/5YOt8pSSFAeyIFPgg0BmXvpDH/d0UfbVyd9PeR7c7rsew/n/7ebRBVx7TzG6Uaf1LlOv7
ganDIPx4LQLeE1wqqfE32Q1vlTt4WgsXIhw49JKQsLLLazFGhOQjBTfbySSFsrg8Fj+lEtAc6VGz
Sfs8ChoY34Av1fw3BCjphKw01xUvqSjhAqYRHeo5ARevye1s6OHpGtKXI/LsJEWXW4/HN/XXcPWE
D/nf45jZNOiKNMwPkAZxqAkH+CJADIeYhsnzgfTH4Ia7TiTERdPmZC04si5PjYPlM5/2Jq9o/MOj
uypRwnlM9gras0yRbmVxFaOwIj8mVaArthCWkcV6KDxrGNTNygdRBVTEyvQ8QJjG5++vfO24Ndjj
4APJnabr2XAvGzh092tN7pPGJfoy4nVIvw6B1YiVquGXyrreBTh2UOtJtYSVz+Ben73TH3Uuvio9
8jiwiS3QVAPdqSFZaNOY85AB0eJAbaA/FQBmt4ho1j/9uqQ/8iFcwtpDTIxCEbvQ3RtDco1JAPmh
h3QYYNsqC04ptlaOxfK2S6qFs6gSDP+u1dgiP5ixNKre7sMp2je01W+NUVHdfEtW2N4VurB4ge2+
ab9d3fgVwx7gL88vasl2b0qqw9rZh2LHQEyR8cf6yw8aYA/zJl/x5kAO9our8bIW4S6LhjQMDSky
SWL7l1gWpjW1SuKJ0fBuDxOvyYtO24ZljYM6nRIrrHXsxX4rPGeSupVK80N20WaUijf2KWcmwJ43
87CcTeRuQzgVj8lPOJrs8u2wIiZLx8A1bIUEuHiU8CxwkG5/RlN+miadzCZ5Wm/E6dWDyvPVwJkf
4UWn6mB37lfUzJS1L3a0xnvEKhqZRaX2OoZlU3LSCTtNEvoejawXv88qYyJcxkVvSyC+i+UOppTa
3qRqyprtqNCLJOFPFeAcm2KkpWLT+AGM1tGpOzprR/sggqThLDkyIhA6dPMJp2HHWDYTFDHaES2N
pnTzK4dub7kUa0n7FkWgA8Hu1ed6CYwnz/GX5lnQGr7iAP1gw71shr+pKJns2zwfEkyM/hUnmB5C
qSTSpK2fzYOc8/6hx0ej+mu23VwqlAVhqTbqmVxzdp/VZ7zeJPt7T422RxDFb8kfrIulUwA6d/jE
8WCqwgFMKAsovkmwenogEwoIdB83mPAbiIQoBZU6we3rZWXM8Pw2D8crkTwv1Xcmglu552gGcSok
8efccnegpoVt66H3HJ791wq0AnHkYmmJFWk9u1/UViRaNzyT4IJWh3XAN/g3TdsfrXHlSmHUYfSw
96fcP9s6iiQ/JAChxrxI3zJxYJs+/FYICtGhAEFtfZC2WpUjcEMP5vOVMB0FHtYEjVc1fQ4HUww8
HAoNO+gTsaHfNgaTvTgrQ0ePXtTPLXcWaHf+ae7DKJIrtmZpbC7kFiXpapNwGs2u6sGOZoqw5TWO
bgDU9G3NYvqwd1+MCxAS/hjAr13Hv/9e+3qqE9+GF4LDGMj6TpOXNmmUaKKF/UqHQw2nGMTUyWD4
tDP+ZJKybh5pVT7uaVsg3aLj8flhI8kEAhXl6iWPzy6ctoPOPcXcrY0aDN/JzAjmFCWMSIOraZjT
RTeBN9vQEeNrC9qkZKKGzkI/eL6U+WSKh+q7l4m9djxXjcPwe7hRIo2lvcg7kPctedNF1CFADfpY
TEl8AKftobfkmgjhpG4LtAp66MLL4XTdgmoAceYDqMkqjR8EIwWmENvJFX+GM2Vt73nxjy4doBrw
4fzX4NePSf5Sj5EX2SozNwPzx6+FZzl8quv8jYVZo5tC1c5Tni0O3fC3hjnlUWq5RnbFetqGOU7K
Ybhe/4DepXRzsf5+r3RhZU8DF92ukRS0/iGckPQ7A5ckGadAx1gBT07urSiiRtj55CI7pHQx6cwb
Tumb7aFMpBBLTnV+6kT84+97VLJ3WrgKOCXtDDVulvOre9lRA7dBZVwRclyVmG5XtMr/qLf9ILin
/J7H1hZH+FbcLufH2UdA3LHxaRL2a4nC53w1oO9xCM9YjF5LUj4HB8nU6bap3P3pQBqJAF0WXmfD
Z8Ky59/ecflhcLXd3nQA76flOY8a5YuLH4Dg6VeoLdNkhpwSNvj20yqwIOXLFFMOmw+SV64HU3qT
YVikcXx4mDXEkUg3XHFAtwtmg7ljUSOfUiF4DAFzRFjT4XzqpbBl0S1LAG5h/gvSJWjrynxmyKPw
OCTlXDgXsTN27PkpCoFf9pesgKZhBM9HJuGao15pbstz/UqwYFTfM8cmCw5oOOol6nD2WXWEdpeG
Bz+G96U/ucZI12F7aoBSx3ht115QH4UmXEGJSARSeJYaeIBc2sMSMn1cZssamfd2J/IDzAVI4dZS
wH5NzMeITQAzrxkUOYpn/KoQJ7PLKF1mGoL/oOy5sYNju1BYfujf0sGrhQoNEppTcul2LXb4Hd91
8wdtP9lPpbDkd0iKwMagaRqjOhrhYNkbYmE0rbusgY+JRUDGzvMq8JrjzsXqIU++I6DvnyL6xo0g
KTdr6J5Cle2ziCxSnldUG+R+EKOUl545PJEobevmoKvegtZi/MsxIqrp5S3Jz08Hpt42KILxJ+4y
NqL3tk0Pdxz9kzKg2xarjhsJga/WKQgAKI6ue30aV+y+v0ev9K3aihyYBFQH98XqCQlNxsi0yzry
vuSHbbdcGVx8XsNsnxM0En2XsTUd4KyvxwtA33TZg6vqENA8oyMezw7ZuL2u04Y1sOePtdkpqc67
xDVv/jF4OIoe6s/gboIaZd+EuS/Zb+Ig0oGpolz7OYl9e59PTtH9lZ/V6kWBjnm3rx+cGQdzJ3eV
43sLiLQzhiF3L2UCtvJsWqfQ3WSalgEnBBhziBFcsQmfU6fZha6Rz2VWQQrjCKvC2PjDZsIQCoU9
nymQlw9Ta5pRQa8osPJnR6hYZ5K6kozMZBvsv2jrzkASjeK/A+FwRx4MdEEVLi7YjiZoimvw+/58
nne22UVhHemuF80qmkx3EXFqWfyl8BixW/WW8tBbolet5EEAidRPuNA3FXUzUJ/6KuOPVbN/j8a6
QBnGJKd2Rio8BzsuHft3s1DPhn3Du7x9ZcwLk9nTDvXozflIaFWkTA+L9tbF4G8l+OIQNn1iDiBK
v11L3+c8p3M7FBAkIqMHg3GbKlXKgBfEkC8GpmF6sxVISvzMr5NmJzsa0it2MLw1c7RRGb4EduFS
ZMnUj33YKaymxTPNG9zNAeQGK7C00NiBZPC7mmhQH89/g29p1si8i7zMAUH2W25Xz2Wa8tF+hglH
merByRU2MqI59ijsxa36Wq4zNcR7IPadRAqfsMNt0eC5E1Z/wvbClWjml7vap6UqjNTIUq4lMF6E
R+fL+Suffl1hwT47FkIJPduwaZB9LJC7cpwK76mSzxTWSPci8dSe0EPEr3glAOupRvUxcTZLizL6
JbF2+pl0EIFaVYOkpbSioG8bnkqiPlSquZHYhAO+GWoivcUPZR4e5j2i//iveYPtVgyKZ717zWQa
MuxmcceECiIsJK68eDLtXTKBdm64ZeJSWCsnFF9y+OTO7miQLSZxvHHqQAR1GXZTOiTn1AShQGx+
mRyXpERIgZgkCFE0QIlYETbvJ64+c63gueW+sn/B3/CgGon/OXk7XCXsde8wiV9oqoZv7rW52Hlt
79axeb55GdWTplT8oQBjFK6qNFm/LPBofS9MZ8zTaKmF4ZsVeUy7HN4FlvZF4yOqpo+JgdSw6pVP
/EOQE9NwmgBtgeN7QUZcTn8xAiHL7mBSg/2oQnzs0fDMUvrisa9ViERTbHwTv13fAjDaYcUviWkM
+p4ibe+EPxsyU4R2/EbM2NHvLzoxDwUd91LKCNcChRAT1ePJB+dKs9QT14/ueG9V1KA90aILfscW
/jua+v8sT8qYz0LTjD5s60ELlVUs4gjz8BtvQD5gVVEzxhSfJo/oo0Xo/xAM4ka1b7SNBpnX4tZy
M9ryK3qT8JiW/fUKu9Ka6MvA5BtVT+kpS4gOP1EhBajCLSSEzhnKCicfT67k70yPSHFHK+FTr3MH
iGpabyyr2T4L9/judcZ+bLhyx7Ff9yvWz9IKAG3sPX7XDFi/1+gzuFRydIYfhOBVcLijR7K79oJq
in7BfgYPjlqlD4QZ06Pk7YMR7IxB4qsYf75IdnJfg/0rdyzhuWUgN5otc8Vgg2Y5qawPVJzLpHqF
G8YuUYD7a8Dp86Yc6L/lj82r/+pta62V+6i9DZGp8fIMMaAqlPSFJCR+S4jHzU1igT4s+rZlcfYh
PfDpkvhVXet9PV/4QQj6tAYJbojMLJjGCiWk0//3awQXU7GomIkBfWhiPbPnPr7ZV00gtJWKOybY
ztI88XscwvhHkckZazHOaQbHCEcR9Bon0miIfggarkN0nh4qfX3bZHew4Y4VybhQC2qPB2gVVcKI
wvWTUNnqbu3uDbDsPMk9s6RsL/Mqx7US5l6obCYbr2TcVQfWNU5+v/W9nJdGSHHTbUJ+muvY1Squ
HzjdGAsO/hMyevO/qU4qM/9a4BSJ9vgi1UFQurRbOtgAZNOHWmQqJBm9w4Y//cS0OkeeK68DpWym
1SW9uoUXx9BprUehnoDgcugajMVb2dmG9vkbS9pavmhafJx0k/fnuZRXgYOYduO3fXL6zy77P2tt
Lt801lLdvMjOFWkLvtPVVgp2eKrCSx9PJpXl+FVSLDu+35lqZRbggORvlii4nwU26A/PQkZB6nsp
lgnmB3n7ni6Hw7jvL+doZaCvFUYoamRjI22WKiDGWk+nBoy+cPiWmbTcwDnFttN2COXtJkIstv8X
gfJ3R15ANlHTLKPYUDYrNu7kyqNFxS1x7ZDRoDpuZ4MxeHYlpaGyJ11WaKB1eTPGVWzujtR6bkGY
jhg7PcRq90QyEHWfZbtIxLvg5RXOQFTi76vI2MrTCPIqXG2hAi6/XaqvTCwSnzEPXXy6sBDtmrjG
ZhFbVLul139TU3a+6fdD6Ez6mRCs8yF5zwbvZTPhv30TqtpOprxfUTVujDBc8q60Pio8DCQlCt+L
Wj0PXkuf9nzZ9JlLGFXxMp5QVbiy7R2YjmEZyjaKhedAvcFYviSuuWHZCs2tyUMQ4+Epmf3KbKu4
vR+GKSv7Uo/LdhXp+7xwksurYbWTGjrR7PlKP9XnQobs4cn0Ud/Dw+8GHXk6pjXMV8N6IMUfvlGb
aY0ku2Tb3XgoO8eWk1OeF5l1Jaq8alYpTDODAhgOLheUaYnM6bgfxSMc+JLHjVP3xeHvTNMbYKtK
xg3z4xMrCAjQGjGgmWrqOxXRCYKIWI6BrG+SfOO20Gt6PSBaElLHxLB2TiwUWyoHRodaPV9uerDZ
SQcDYh3kRSGp8a12V8hjGnjVyQoszSjwHoE4xbN5zWPl9mkvzcpKT0eb1fQk/tKDnMTywEqVylH+
1GX8cpdu6Ip9Vz8+2hNSNPYw68n4jyGQ2DqF649jRuBQY4MVrn9wXS8JPaFnFpQfXPfd8VKmceY4
D21NtA5/7b9Y4SbMapDnuBlJ2eJXc31CLIr9ERHJrP8mSLXcvXXs4bxR6Xyy9atsMXnScHjuqTME
n1YvbHH9v/6tRfgKfQtTYI2/cNABBqTHoqhXFMcbFGEiBYR9eMNCWH1SGgVbuTKGApvfMM+Jr4Ej
pfwjixyXC1JpsINxk2yr7dUGmiupUaHVQQbynG3kbUguYvFPxA8tUIqXipjbHyP8RjfDWqJv//nE
v+GvJaErrJkY+wHqD9GjKM+MZnUqXxKk1eeIha4jQk7+2+EoagIpJfyyZSslPQL+Io05QplyfyBl
J0HhNAp2sf8n5/cidRXzLtYcC9Gi3DTP/Pm85jYWjo08YZqIiG337ZV5B1uS7/DO/PfPPC8Orzx5
AbUjKspbETui/0K7tXnqiptq+YvLNEV/PsK0lI3hwAKrD1Xa8EuXDWaYezsUeuaQfJxERBYI6P71
zhflLCBEDDzH1R2VL2M27t3KJXtC7BPgrHLnkY7DcW/jLmIBVrcBe5C0m2uLhdeTDRvLJR0hlFfZ
6mFdINIUQFq52q6NAtcJ5xQnx5AW1xxm12ayLgjp3iklpYj1goCWAjPet6FazJS9Sq1Rqohc1sZx
JBW6ZzZnG/j/G5yhAqJLWX537rgRaz4d1H7rQQwCsfQf4igimuMSAiMTEpr67KdEKv62ixKMLQKe
tmgYZaeK+FG49Hq0fAWBhVAcCZ7qWec20lSFjtrytVoMOPNGkJrA2Ip9Je7F+/S2PU9KIiVqkLvI
0O99tVZw4f0YxRmibaYS/qpifRgRyXGvmVZMps2RMQeEiFCT6hB0setVXnpUptAuFI8jhcBAaoi+
9x1hNJI43gA/SOHdrwdvFC984T8ouOHUuDIMHvfLJUnAmdb39I+hDc2a2Q6ggAspS2Ts7mDpIXAI
qMt04WKfrm9jT36iZnXRofkpE6QRrZSM2R3wiOCFFvLpQhwH8bPMkYCotC+Qlcy1VsjxV5sfEBrl
bcuPcHgdL7BvHe3mhuveGfLCj/jnNG4QBdhMCTxrNge0D03+/tpgqStmqYJpPcNrXsIzzg7zWjlA
MAAsJg1LczO6W4nax3iq1O0+Nr/ruK7hC2/1Dmp1IZjYMbQye89JplmmEFfg52xRL7IDsSMB9zoS
5sv0nqjHIqxQCrW3MLajdm6byEXCQpCmy19jIKnCVvMyNYgO8l4KT4UI4aZEW/VqLZvMDMjPTj2S
lujVuAzJspQiyrSiAWLKb2qaOhoKC66tUv04CHyL8094iuyUWCk2tIhthsNN5xgT4MNXDCBf/9Yb
EgsV0CymFHAhZ5uZszDR2llwzr3vnVQt8gAsQc/VPwoe4wztqqAkjFOoEUQKFeY4PX9wEaDbAcYd
6PtKwclr+ax6LFvi4dLm8QD9S1fwbfKzu8Hqf+aHKmIl7dg1pZMK77Y729GwGc8CcFWN2V+lINMm
95bRlAkV2cjlhe6+kEqETAaOu8WMT0UjO8xxgByW0i8KW901+JPvRmGQxxQewu/tGPbFL08fpTzi
/c1RcdgdiaiYNauRXnbf712gsv9i3rENxxoNpqF6rF6Fm4mBB8/OVWBvVvuW43/cWpyoBvTY0YE+
8Nw9E6Nq7I9L31CSg4LHX6wf1rlkwJl04i1JzYKWdMayK1TBV5V+BGQCXNeBu9569H2NTHrWe0OT
goVAPghYE2iBN5ZEWPsOGg+d+j3/FbhhcXt+E79y5y/KscJr+6TMVVx4QnpGXmmkt4t3s89tVT75
wyZKlJD+2bQby2yNFp1ZibrDTLYBM9e7A1AX1uw1I7B5KQsvgWuOFgQ63UkVP2MaPZbdP0taKOsd
9DdVHEdYwxzGOzesm96/BBq/2pGTzx90DevUdkkaa9a33wJaR5CGlZvQ8LSBRLLlKjniZQgTR49B
46wCZ0nEtRmJUwR6iu9OGhRGx/sCCLPuwhSa5O7HZjqils6W1GKD6y9uw0PJM16Mpatemv9/+aI9
m2U34ZkVPdX7hP9G5aGWUptKClZbA5oi9KyPJ+2iY8hq/wwMmrhTRH5rW7giKINKjxx41EYWGz5F
+ckuWX5v6EfRdtOwx2Eh/X6x8+PRm0sAthSvpi1ec/DOH2iT2MlshY74snMD4Dofs34GGh5ElDDf
TT3qX5fO7h7SRELvU2CIgVUsTUiPh/jmVzkTz46BDwSF7cZgx/BHQK7HvjzG9DCYwbI9ebfdFPzK
EesLECnwKjy52b5z0C8ZZRtt4UlrtcHVNUWYMveLDlZuU2jUHdfGUqLOeJAuF3pHupOfcYlbuD1P
FcSKfwTFdasABuReX/LvInErajI2x/gRBYaIAqq2bkK0B59GBxvo6M3PB17TfG1unq1FDaG/akt4
7FPDCtwQ2jJRgSsUFTgXLzvkLt+K7/3JIS8f+eWbY48gDcoBwj4B91w23OPPPyg8uXIZSirQPA76
mfTMkTga7b1Xmj+fL9PBhnITf65YPoMZhuqZSarx9TS+bw1k9p+C9Y2AmZhrHsAuffnSeD8Ic0vN
9ZNiLEwAccoC1nlJUVtVxU9XvsaXZmijSU9pjR8r+zwiky5S3+PqRsvJIyjBHfs8Ywt55yhAq4gm
IgGkAi7cfHZ/uJ7RT3RwRACjk4Ru5Q+mElCxQKgUJtPyixBs0upaTSwtTSKHXVfUWeWcie1oO8q6
wothVvgu6arKbpuR03MtVeW86VGbGD1yASDm+tleSVw05wXX81akjGBT/HHK7RP15GmOEmj2TscT
z3NOI2pGj6W9WWM1nF/noXIzxl4XaI/ibrkUcNl10Ab73jyuwUqWK63iYfoCHQCefIkVvr3hI6NL
V+IGyuRuQm10t/y6GQfw81kWnitMZK0GBvcEWdQUnIwXbSWfixB81P98djNWJB5D+rfDEgJ5Qwid
hJPxHtkgvrGBorpuc+YGgRWMYKXW371G8IY1EWvUade9T2oan4CUdpYV14Iuyl+tY2ps6SZx+r+V
7GZ0rpBY+HdVg6X7BeY7xJzGDuvDexUTmXUF/TbCeDDUhalBtm21Imo/KDy7tkpcZ/fsa/M9rUYn
8S0virbHUwX187rJTDbL8eVW4r0cADEyzc2kHyiJgR/M49WVNgBdc4uPQZCJZko7QUf4AEyzpjUK
/e6qx+Axw+PLFBhJxhT8Em98TQ0SaSl3Gml6wSWrFhdFQYwYWXyrr+UQG/qZnXH/JQu9zct8Po/k
Or78rYM4FhYYlANt7wOpr8M+rklZnJwqrvOvbVxBOHFqE/dzFQM6f6/RExuA0TjKc7jRqF0ERd50
BRfF3L+hYBnbcJNgGfKZmC45x7DzQZfB6eQvr9GI/ah4uE9jxVs327mp3EWjZIUpO4fv7zqE4dQs
zD40RRvj3ivJyL65LMSWF9Lp5bM4VBggWU/cArZSwR6GOubcXD6/DdZ3/aiWs8y6QFMihLvl7zYd
VxLnJYXIe0aGKUrkgE0DLTLN5Srcd6OuBzD/iBdvIlDL7laQt+mh4MIqeb+a/Ha0haN2RTqIJzEl
E56DtnYJOeddjLiTmrXhr92GHZSlw7LNOELtSom92O3HbUPmyaOWebztOHJ7+5ng3fl9WX31yK4r
3TO7AJgWI+AvJb/yN1mxmJlRC+idfk1onU+iq5Igh+Z3cXrJVjfwNaE7qvFxl6QQXY1BqoOJAxGu
3hRMTT1f01DaHf5cFSBIl6HH7CKtkijKIjsSw27YLHRqCZTpzIcQqBIU0C9pva5iZDfkM9QPU8Dy
MD3UVtzGnKDi23ENza5suu3qSzxU5MoUoRGCl/avKcprA5td+WeKRZmy/COcsd7ilOThrjdbphM7
MWtRAmQurLCQmnTGt3whFlJIfi5tleu8268o2/Be4bkbexQq14uMkdoYdS/5Dkt7GNyCcVqVCUr6
Z35ZMUVNTfO/3tiCVvpoGYttMK/D6T7eiOyfNtt3JVUPLyf+mbbkVYQ7Ri+QyMufsdU2KTzsJ/6B
wsO+fVrWzYvFUuPnvYEEDz3w8KP9Z+nXu/n7UMApy90VIhMuj/35LQQyt07t57SzZ4fQ/ZKXYC73
YU4BZ+vUGfoBxLvTIL5cfrLitbkAEgOTRU1or5vdsttIo9mBqFlAVT5UcRcmkV16xcVWqaSY0cjA
Xx4eOTOinGoe4UHrOLnIbphqXep11qc1Q58S5PU4obLsu/lvVtUzz+lC37yAP60W1lqUS9Ey6KZo
WJ/IDzzp8zcwe8rJnj1OFzdxFDjV0NUb6yC28JAe8N1zRFzY87VEIa57M3QqPiD/sJII9JkrJiE6
Iu5dzvZOJZxGOy7HBURGnC9tfq4JAAe0g6Oolq0iOM8npwadB20azf1meXQiuoH60ocWzPp9qCCa
qpQlTZFfC2vjXAjFyhRboq3xAqFpkHdubTFMKy2zfVEQ1VgPZZBLFc5ZrwqFTTMmkugTp977Y+8g
WFJMWArHdmvYNObZqXu4xXp097UrIyJStJUxHmK/jlPmhx7cUj9KNx/TxkN9IbYuMUVOaoEtDQ4V
pfkhKfcdRI+thqrKD24PUnC3vl9WJBOT7i5iCpKdNGkKvxMV0KK8hkQ5KB5lFtynA1L4fGFTcbfW
VgaWt7anE8Rl7LewKZl8aMdU1F2OSETi1hFi0OYEfoQw+n+ruLzBByZHnOsV3Ct9V+/graUHvaWs
STG0uLAnkWUbTPYeVJoSQfwpTgYacYulwPjpkB6PJtqubB0iODvoWd4rFvHSyj56E37OUJWVJI7j
zj3Dp/V0agGx7ac35j2H4QUtpoXM3AKH9DPBEjXgfk+kZyd9LUypHK0hrRqD1BuCVQLsAqcakx3P
ZduaogG2Oklz26I1pbyii2qyVKrsyrvwHZcSPkFjSyIJeDCTX0DBAex6Z5mxTcucka3wD5hD10OG
3TpR6BnnWv2Vz/XsFoSJLqjCbMTeTOmttdWQXmQIq0yjeBH2d2cMJUmK3+0wfq5WUvJ/pqRlhrV+
1BzSZDwAVmC3620KYoZW7aMvK8QLYT741lmVjZHUcI+95xo2a10ZAaM6sEYxXah9uLwcs9sB/qZL
18BzLwmfSi3Xs7LMFfgC3kxKd0WSgg37JoNiq5EzN1MfZHKsojVhmuK37S1b9Ra/3qhJj67lteo/
H4pojblCYxor5hXsPGZg36aFwVGHAB+IAXAa9LwRjSqxhwuYY3pSiJpmoXdDc1qUnsSLlbzLFkgx
iHc6no6rijHtwv6gPIN5cKELb08jEfUqLa0yAwdUxl1HEYjwwweprqoxUvdUrXIbQAZgj0SIP6w+
VPqxg/YkJ7xbCKftlwptNr4+efuQMyHwuPXyerBYJAkGvJ3NIDWA0SZfUYqJKDyQack0l2Q8gJMG
ll/6nt3lQTCRkSAA1hPwcdfvAqC5q52pCgwh+Bk8lDytFOg1oZSKCR0NskfSsygzfO/WJHSFfPu1
4NhUP6eMYuNimhPOEfvIqmAeQ4Afym2GIa6OVqbqv7qxnJdn1/QWVZw1UC923NSh3NZ67SOkG0aN
l/lgsvAgFRsTx/d/+sq0iLaw7XNk+gGgvTFvWB21x8SWYqPGyllBmra7KRmkF31tYmMJh8b9qKU3
RtxUpkG2KabkK7MyJHrvz9udQrtYv5vqMp3ZxCcjOQ2G4XRkR/LFdbfDiqcBMEHURwONiTMZpx70
YsWwMvbey82eHqNugxRwT0B5nJWTBqWZgipwKVNgzbOwCVGKR9f9q5abc+oO1DXbI9fCKUh5LUlM
zxEB/gPZN7RZeCVAvbAj/oxV3ApmkG1YaVf1AF1Ob7BzaovTOqGmV426A2KOsg3H8BfXAa1AvfG9
7Dbj9mX8c9cblebiRk7ORZ5ydZws8nzS90j4zajl8u5OCawf3+wCPMHwuC1B7DA0TIAGoGntUREh
1XhqhSVC1lL09qjRDKyBQ20AbNoMz20gqsGQuGm9Lum/o1zOFpS1EYMAya7keu2vbkxy9dE1dzTr
+1pfnyvU9aD14Frey9b6YpqIcPKnJ+GrrB4b54j8anlEzXxSQa0ocOgH9GirGB6RydtJ6G4/Rd5o
f5+Ebq5Fon+7L64HX8U28zWyOrL1e7sxJ+aKLjmsoMqfoPP+AQUbz8n3m0ma6uMIFoDzdnvmRP/O
glPX68OL8ktM0XRKeijkPR2gdmKxPKUSAXSmnQCU+ad1XRGWbKT+cvp2j2Ui+Bb86YbIULsc57IL
GToeoCsysnRT6ROO249ZsK/s7lQ8DBawRXMLraZvLPToGzjkCkV7l+eI9RoRbx/jX3BDJ4xEbGOg
p0Eqnw2hM0Tw641uJSTVDzlmbSmoLG1A+hnyT95wGhhAyd4X6mgIfV7YrMsbREAPAPRVAYow3iFy
ond65125qg7cO4yTylCScseOk8iDvMURFwDP4oyNt7oaiSbEA0HhXvGmdMco10yYIAd0U/4ZGy3v
Fm1sZGC288nFGiKJEfjLrPGd7ybR3j/uHwBLyom/4ihfcQoTY6mecetiFAndeJi20fSihxT/AN0S
Zr+aQcvCpuNyih73jACRhU2i3KtYFRHnQXvyohNsI+nB0EvAG0H3zeVVAKff8Sg1XUF7IG6kaWmo
szI5TnHEjGAlb8V6Y5io+Z2TAKjiFAFotrruZgRBeDOUZRh2egTYGMIpgb4ubmunLdm6ORZvVWZQ
XIyeVNSpBT4LBvOUvUZ52HRz9eTMeKyRqHlat9j4U7I3dqqd0J5k2f07khoHu/rY0oSg0sMkN0NA
aUB+PkFvIOMqtgj8Q7JNDUipmErm6w//R+nzhlDDcn/4706KK6U8SKyf9WkbFNyUUgJAUPmVHFTD
vyaJ2rJYI+1qRVzAFnGb1WXFsCF+oW3Dc6HvOcwbUqUZ4xal19yrrB7N5etgvUq9rk3VnctTvfaU
MX1hBdjtfWOml1bY6tvUtANVKuqyuUss1vW3Ve4gb1Wv9UH/8hyTyjbgdRxAxFxLpBaFNyjQB+xK
qZKycDnkJc04EdBCy6wmX6++b4bFy6OP/ndMN3F/EvUDiIoyGjRiEYl2AS4j3tGvoilZEpd/yQWv
HPmL83e/foM0KVF+eG4OqBNv30r81pD5/HBeX4AMWDOgljT+HQ3+Kqol8/stRhNEy5ubw9kuA5S4
ADjWfnV008YwSuXygTbNY4hta+C+dY6fZfWsF6jQhDhNZnMfXsc/p8JAeqbULhs6og8pf1l+KZYQ
hfQXqQnueSbuqnnNjORsKSDDGqkGTtlLilW1w+3+r0ARKT82Gi+w+i9n1J39UtxuJARQQA8las9e
yA1SrkJ7ii0zIUI58zIqGPRHqtLDeQM181A8ggNCi55Aqt5d3Yix8YDvmY9BTe9lnza+OAv/dN68
Rv8VjGkNSAQTl8GgKo9k/G5DLm/moZ5iw3XV7OEl7SNMQ4QQj5CUDbIYy9K1gAN28y0wq4aE6SFh
+eTYtB+bq1pTX1I5mfX0LqBjOwzxVjZ/NTm1aMy9qQ+vHQ76CHBwy70J9EVZhyJAvi4HUmWcdPcK
edEWu94GCluhGHXjfAatRENDGsO0XStAZNQMZP20XAwXmM67erD8zaedj0SnwJ9VovjE61x1kK6M
aWBfrXqCpwcGzp7JbU5Ld2ZDAfaqxXANV2oK2RFu/EVrYjbHEUBuVQ9MxArp9a7VJ/RwU1656pNq
KeFKqLnY5GUXtdrFpuhbEKDRruaQsERyJOZGdK0IirXdPBvoKwPK6IIr8VT5kcnoqH87hJ3cOC1n
Ll6tzx+4nt5XpGOUMkVtPMvuiK0p9AXfPlUzV6ZIdOR1alxWRLpohtnm2Db/ZfmpnTdDLjJz9HDd
hk8BqxBE4V1DDGqLcybEsfaVOM4J2e8SjHelBJ/1RjmNhGkXQz3QLwCJrY/VBZ3HRYy/lC+kL2bj
eQy6RPvdiskC3uEYeziFF+ho8KcivhKQQBywFWimCGPGSS5JJM2ZSbwtbV7QwBdMTfydxVYe0+NW
ao9emntJADO7xg7CtjEvBlbPDCdj/KRUWD+QzqjebD3dz6yMRR7kvTsHoAlwgdCHT2HM5+wcSoSV
Q0tOe0u++VI1cZvMk3jTPJ9g6zQLjwrN+wgTeOuQ59DD8/ofyUguT5Lef9Vp/x0XPPjvVEcL8yfa
HS2oc6s5zOeFEe9IpjDiygd8cKxEEbBRd5VU13AHjyLlJE7WbHIBIqk+mYJH0kb1YPqwYB7CVDhT
h1msHBVF/veE2tMMAzyd481OgYd0iPgk8YRK6WU1sDAvgisDHdvQA3w7quWo1kS+W8PKRLkkI6h4
e3+isXWQmBBCl67VxxfzDQIsFpjYzHHtI8cvyuG9tedFk/aJdgO0Nt+sv9/8U1UDBOSn97mHv9qB
Rb1gPEiR8dlzHoXk3nP5IW6eleOzjgtEFd//ad2S4HOgg/oP0ujeBnkEj0dQkqvxxIH0tCskO9LU
jip/VtsimbBlOj0cogJci0S/W+Z3jkRWhTEbWx0T9gTHL0ZlMcpsqL7CcbKxp22phfHu1HeFaIj9
wUwGoJsFnJI+KKDtePwTycuYjvwiwm/T1r7IeAzcOcxUpCorT4kpUcfaYaHS2EB6m8pq7inukACF
vDRwLhMq28g7KyapHt17cM7fCfuFObdT4glXGvN0dh3N2I4TPp3IemzXSueXqb+5YP+hQ6zGHDXE
gllEr+nqGkpUsdnfxO6H5m54kMxH+5JCmdkvtLv6A28L28VaDt/5f5Xx+VjARpz1C0Y/AY8d7PHt
KBr84xzXT5nLS8aTyDDw3FzolUOq0cCtd3WsE1Vg1yQ/U8zmTBVEtMTQs9HcdR5cw00ZJweR0wyj
cJhJsfV3FFDagVccNqcBgQWCh4xLAalfl9zCM81jtmYAND56LNsl88J3UC1xrFJVysEQBFQNOwZN
FfKuz08jcOht16ugOxHYTMBqdpLLb7EVRXzYSN4wzbHfR3IEPvpFc2u6SDhlvTWvZutXR+hqve+R
wNY7za4jlvjyxF1LfK7gke0hF3IZfMjPyBP74abcNDRtUZk8uSPP12og+rs5Mtc0g2RhVxv2QPo8
Y0Y4EyqrT7dyFs/aOxxrFVcBlJ4qbrHIR8+rIxANehIDa4GjdwbpxNdn1MvisHeNEMXnib0hyi2H
TYHa8ltl0ZPFdLxOm+W9nHEorzhMHj3Rzcp53YcR0HoFLI8UTt8c5KcikeB2LaZxBtyP4PE+U8y2
YO//v2ElodrQKBg2C8xY/ed25GU4vkuTU3PxCEp3EvDyGlaK3dv+MMAdG1lZHmzaxEOQmtuJasRQ
fOdYH1NIVH+IHcx00W85WGWvUFqwS62jLawoyt/tiABo1//rO43dJ6X3Uiag/VPezT6e+Sf1MbVK
SohhoDuTJ5u1a0y6XGEvQR4EDe8LA2j3YIucjD/tKoaaZT5Oz2RasL1E6Phkna/TeOef4sOOAWhr
/FcThvVn+jpe+wHVubyaPbnntvUje1N+HRFQmJvL5FnrKfqBlWXb2iRcIJ3nFWyRufD/DNsSaYoJ
93rU2xA8Wph1m7WqbVvs8+/53r7B/1RI0JXE5Zjum/FcDSzf4mP8iZEyE/ZaQ5xFtfkuNi8qtb6c
fmH+lqvRHIufecMVHaFoFsouICSYufqXQvc75XS4RMP2v4PFo4dXxSeuaWZG1RAAu0a1ZB6qQjjd
bm8UFqxOCRfNdD3hrw8WbH8+hq82ajGH4SHbW0mAN4jXWSRLoNmLCiHVqnX5j/jv6xBQu9p6ts6M
JgBIqH0uQkdx/ndckiWoVeCm7OazSgGUr5GAb1LaEyiyB5T6gTs4/p+jaRZXiL7+2uwV4LAtKEj4
tZs1/VyAULWc0mExZgBpFUBprLPze9InbFxCAYVRUu3otfJxobtGpdJC36CdQvC0E4W+wS7U2qvi
G46P3OWAWez9xUEktL+IcAx1zdazMrPpZ+zofU6fvERuKAejdD+CGfLh/pI8/pdQ/It3VxBmua8r
xscP5tdo244deudAyd26/9drVFALWOFYJSCsSYd8fiKZyv7tLYRMOx1l1uKY2s3UWeP2tP1TsJLW
+aUVwAWH/avY9e0YrST4J9H7woFQRnCWjFyx9FVANnSUJ7tnE2iXtBsbJm7HP1pqXxCF6fD7IusC
zGviQTKPG1EUQbGPDU02YWyWdxOAdd2gk3LKA6Q1kr72uqlmJShDmp3j9Php8AmuiB+OSqVzIL5x
UkSna2LmKdQVFR/+/dPO3Fm0J1wSHTDcU6OI/Uy9GqigYQCU/HUqbESkyrw8mHS5UN/XqTQS/cKD
380gr1xEafWW4GNDK6JpGdgc+pTNCnRSESutWh+hetTHSsNYgEIRjwxAs5/lhmA2ObxFdp4R6S4v
VE/kVILo8teWkSF4uaJWeOdF58DGpspEX7tq6GbA5Nqi6BERMaE2/4qDbhv5XWuUvzq71KnVGaxc
4L8b8tGPtVmdzKkJl7e9w+dGvCvM+r/1fKiYsOhPBIBNPpa6U8abiyGYjnO4ni14xJLfJDhHi4Tt
pqrT2BMnuqUEWWu2TjHFis43LP0AtRHFI2KW/tLVq5TeiUA57H3fqPugFhkw/YYNSuwSg7x0SRYL
CBgNNoA86tYVrd+3hJbXNf+VIBkJUUX2XrP37AWaueHfNyRJcUuQb/yMgvA0qVkezE3tKmOSKHnw
ZBnqh+pMWoDu6fJhaxGM1XwMltZPAX9yep8u24umYVz0m3e8nilD6fndLAJ76R0cg/8q841VTTV8
IqZnBSN4uaoxZc0Kef6BTZnrj55Os4XHZkz1r3wYpfZaVoZOaslnyL6jKDBDVlvoMjgpRBXX6qGm
AWOVZRhILPJRDhTV1m4yGeWYgsdQJhJ9VOS8RarplYTPPUxvijAgJzAMuL9fjFwUhJMKgHpE8E+x
MgN3vkbr5qDSwWCsTqYeFFp7aXAtQgFKeixF6BUcEDW5h6LMKHVxst466VoE2PhmmlIi7rrdh3er
TCjZtwtQNVmOGpUNTMXur/Kne0CL/x6HOyCZr6zz9+AsVTfq+VuobfL/hLv6bhltVwt2NzjojRb3
TYUGGvhL5vxI5fytl6b7zcUROkTrACsObrfwd7wwuR92nRY2fTccScwhBz84UZTFkye5ziNaBRRD
9gLiFgUSss/ww1jz3H75KgEAe+5UQ80M78FLQEP4rpE5tyKjS/qKw8ywYPeY4tgpk97jKZhp5v73
KwEwfSDHDl31KfXPC5WUHaFVlXd081l7QfsXc3lideEUhvNvq2xwjzLHs62GTaMJYx5Cp4PgPFyR
gBuwcCRC90ayhlCPX4G3eGiduButEYiFPghRWqo0MH610DA189gzQ1xzd509O55eFS8QABH+864A
LWNq7b4U6Vc0YwSmOEOgwTU4+NKkDpD9xy4tBCegWKbb8Abp4OESs82Iv9l6IU6U1v91ifBy0Nnf
JZY3IYroIpEOsRKrm3aNy/bp2kTrNmQ+6OSD2TPJwCrPgEh8L0Y24T24/yc9eC9/pPXLn2I736HW
DwvuhMoqBkjVcM/bJ9C0bJ4+F+iEGklUnYBNIj+7xK1ZWi42tKEgfA+tqpbHWtyXAs+4i71iSMzz
bAVhkPZdz7QjGfn08j9A6ZWciDS3MP7drFKroYECBNAH8o7FUgiO34RTHn+fwRVNZUC3Ixrz+HeF
JTlIUJNzuLu1Fn8wHYh+Lo2WXvXPsHZBqvlvsfxgbuMYYpznYuRbdQQ224kKWbM1kVYGvB8vdUFU
v8VigL0VOSZYn/PGhhBlOykeODllDVkKePG7Gw9UIsl8kb0MS+jwaXnPdrap3VSfSTf2lHGS+yJ3
LbmzYjtlcFJFCrRCkcHLg64YCn7maoAdPHvWJqMQ5+Mh9T+DMUEh3UbtL6hYTuNQJePd5gHXDqA7
/DAYzyrjQQw0tQ8S96J9K1tul0UHzjR3iFuUlU5h44e+iDujtQmoULwH3CmOeuuvOuvFq0SjZ5Y2
+r2gYe3GLKqMy00AHZqDvV70w/6epSpxGZP4bR81TN6kkDsbM1gq6lpfgLE4mzem5YOCqlp2bbfr
qL0F35EcDdO4HCUSwGXL+Qs1jJKRF+ZdSYHy175avOw8f8LuCZgKMzwZ4oEA7r3t0khTbMD57tVj
ceu8gN6uN1PKT5iZxyl07OTpqwvcR4JixQFFCMGF62FE7K/ND3ghNPBauvqZC0aFVPsVQDxTiJJ+
CsJwBzNm3FhKj3TQ9sB+U4RyhbsiUimOy9j1U8kL5oD+9Ng2K8JzWuSUdzSRKaWpP/0/5W89I4rL
J73E1PfZ3HCiD3hpEGB4jcxhTaLP9BKNH/N3qxbQR0uSl7VF80o7TiDv8U23dfidcsBbV5QvRi8L
ZnQV8YXJshk/vPIRnc73wsXofBTx7IXFsrvwrYO0thBlOwdvTKNCwx0Qom4HUdpHwvE736++Hrnv
pHzA4fNe1G/sCOysFdjuxwthuMWsFHbGc9pl5AdpLYu0QX/UUsh0dfHhX+a4U6wWgF79aaPq3kON
aMPPl0341zmm6yeeXontIACXDU1hBnEGFeER2gImG9ki51u+N8+7zps1SpG/S2aX0Yqmt05MeBnh
3YF1hyT0hVpfag5T1WtBmsRThWNQjz7C9+VylLeO5f5c8H9DpN8KPI3rFoUCXpHExXVuXIyYI3BQ
9/y0bokubhKMev2gB0JrHMLi8okeuoakO3eJaHDAn9SpTblwWLTkTHLA+w5DWotG3aApH6iuF+b3
XOpGGhkKvXchEZXr3jqIYk+c8Su/qXmbsgly3PokQswgY5YQjzC9pa3I8JaNFpl5zETWTdEwvT7t
NQYtrXiaPGUVtm7oxa7yMCH7YXUhLabQCiQ8HNIPR5ZJyZut47P7F0S3uuuxuKxtcqWaCRcNOcGb
N2favQZMSI617EGvZB3HSn6/w9K6+UM5F8pZfSCZlu5j9fTlI9FJ9jE1B7WJu68PHEpHNckWNo6g
X3lF/Wvv4/5dAWcGsW+QKqnKwOS3g/QHNdZ+ZuhKqxAQWgVjW8W1VvDATg/EMV4HXjzqr4B306xH
frlmnt+wbe5d2ZUZoXbgBNlGKTf1AFU/2EdIEF2uQMmnvumDIbfdnwuXP+qQ2BqqW4hKQ9K0Zt/Y
A+nc74uKMj+qDIp45Kyoklk6dl00eXdtQAAxIzcyp9jjNWNUx0UsOmUHIMhoC7lLrhB21izr0A4D
o6DHzQCyejfbG9jBesvv6UPn7UeVZ9xzT3aIf+hWmVu5qU/Wyv2ADpP9niHihmDz2PO0Qm96Ab5a
q9Ayf0r1JmJM7W7QpiQiy9xmCGFuwmaMHrpPwhT9y2ybkgvAztTqs3+4WaJeChl9iGzdi/OvXhQn
BDAUwWV9iNaOxoKh/8C+3tQwKd3InJlwJiuuAltX4I9/fb70BKRFXEvh5F+8/sMHQQehxfJ41R6T
fi4ZrWfxEL46NjVLyg5bykcPJePSRWBowqujzLaW3iRkQtqvP4LcT2w5juwvR+fd4nn758hb0SYe
CMnzZu4Fu05ocruqys1Sos3VfvlygJMlB79uE4xqXWWHWzKHGm8s8xo0qrPB205OSEQeNUOAkZ32
9sAJ1ebJsFeB79ZokmUU2gynIhhRTlCMkqyL/b2Sa7ftvvCBcryBuOyAn9takUOqfbJsQUbws8m5
ZV38m+MiVaDGnL+MgQ/GB4KBFw3zUDgk9g2Nh/izqWDfoW1FUT/bxrvIcBga8ofsrsGSZDjb6eFR
Ga97gQNtEJBuox3F40E84gR55XTSQ/3W1EQFkSUCLAxd/SgRpM99rBvyBELtY+t1NbdONCZ4+BLO
KoF4P1/oUtFU8W8vRDuLqcTEQEm28Uk9LSVT0FNiqh0SS3z8BXnP1mMiiDijNZlfvxME0HqSfC67
2Dt2/CEFwlB2QCW3lJ57PO0GUXjgAN7UK8+jBSfysfo7vENcLJhI2zuTgzE1M3W6+zcP8BtN2DJw
JgHbSSEEc69lhNhDqL2R8vOXIL/l2EZ+nFvVcSb/haSn74l16p7exV3kkfeeolfw1sGofpOm+dR4
MU0egQGJBB7eizJa6JxLDKhqstIxYa85Dlx7TH+ej1w30S128KlB8c4679Jr8x1UD7O04yqLb5lA
aofdwePraDYz/FhADd0lSZyszDJ1Y+pYkP3mr0k25eSb2/NALlSP4lKT0ETgSz5EI6TExR2+X8pX
jqz2bkMn4994QD9q4acflcLn3b1shG3AiR8eohOeDAHA0bZ/E4zCKNBPT8xGD+iD+LKWYZYORXhd
jl32BZAI9kmlD6b13+eu204KttlxJTwdCYXvZH0BJyWrNeIQb2KE1jgA4UXc1DwrTDmVcEZVMZDD
mQ6DrB6vXMu2zJSSkKe88sdTaoa4CdJjEJsy2/mphYd+dqIF66aNTGpwxtu/fSMqZydym1Pp+d/x
nPvaZ9EjZXS4a0m0C691Sdzf2CYnFYVYkOwuFNUmBrvO/vi1qMhIiEjdnpP96Djgms4+P2OBT6OZ
zQ1hL28Ai6B5ViP7mltP27/LcI/iSH8mWegsP3FonxaiSwaFHZ2wfUEmzj9Ck9HCbWbB9vfJI3Ob
aMetNZEkHRjeeAywZne4iLGaI/CPgXAnUSMDwkc/2bOi2kq+FFyLlzKhoatNQREeoJLZDwbpTOUL
N+DoJK+IdWLBMSUdiwQUBnG4oac04DYaM4KMXEG+hDMDMglZhW70abNUqY2aONHKadWjtKlvxWIk
bM5EJsEx/G3xWLSenZNQEeOGkSkSKptutmUchP0g+rpnrWMKdnrFb+kjyz3qvVUDegtQ1d2ttHD9
IvnFty3PdP2vYwUWvIn8Ufp6jzN2Vd6UWhoqS7dRqEDHh/2rYsGhJ/yvkLy/9GBsdktCAtn7MKlU
HSN2lBJ7P5UNbTs/AzZoOSO2hXse9J03wSMzNdyZgacAslTyRz4X9Yj0mMQwoC6UyfDuBNjiCO+1
MhprMbPKfR+wz+tiMj6ENq2KoJTxDxGkGUIV5DcpzcDcGV0VeNVfNkjQE0WkOewfWa2fzIj+ilIX
BClfUMmfy8pwRMccrM/YyIHDtTWGVE0WGKuRuqB1W51ULnUbhkQE6+YEIRpHlIt7qcSIjO55aBJK
VqznZj7gc9SpDWoXaK2Ph7im3f5O4ekHhBw8wEbPm6koKfKCvfeX7LhFRLIYIhcswxJ6+FV+Q3DZ
xkVrLU7xOsEu5Baz8oqD0g2/xpd1+H234Z02HEgL9S+FLiQ8PrlhmrQ0McTONSaJcraDvY33tday
R9YU8Lvya2bYtNH6LZ47RLPoDmaAa6IoMqruMfms/APORskgfECq96dG3jLzFHu+i7lQhNQ0e47E
c0W94q8yW253VcNTgW8v5h7dqYeB9Qgv6zMVJvikEUmP2hz/d1dDpPgDiDOZ2w1L19gG2dm8SKn1
mVUQyTkuC1QkL6A3wLQWaH3CQCmrOhHwLETsbDJ8j9cq5XbtoSM6lhPu9DTz/5pBEfSzW/1ngN+J
WyaQawy90wEQ3SHKn1uM8riTeXkXzWRvAC3kDOJiqDrKI+WWG2PqLuN7jp3bAIqSFoI/6ytqBNK5
gnqc8LuVGVYSYYVKZKNhJX2XRucmEQIshsRnPdMa6RBm0F9dMA9MC5zVXoQcV6VkHbs9UmwnAOjB
xGnfUud5H9g5u8hbRrB9LFwis3j7FWnrQoCtsLeS6slN0nV8xajONA4pLPl1+E8LDf5MAyqNNAJ1
8w5rrGz5OnkJi3Bulj51ilzAHiiBlWjM79itkvdmEXagTazEBgA4EzbllKkcQ3G/X5s0yBzLjOKv
8BT115BNQndxXDUkySo12YNZyvDrTYLt4y5grhqQXhnF4NAwonCRscgUXAqe/WXHh+paLap4mu5p
ot4gNLNwI8zePfjqcNyDsXpCJ82nmsMcx/7yvYvMlh6uQdsy8tOqYTZcA0ZIITmYI1v/Dg586th8
uGaFGX2yzGT5RCiSQp++TciMQA0/gHmQzDDjuZD+b6d+IlqGSWMHgnm+FZMGaVQcPDfyfDxHIpNj
+y5WEs0v19FnLHMnGFJEDki5se7UL1boFmzNoEKClrN2r0xNrjlUevoCyNSNJPWUun81YQi6Up7z
oXAkVG8gk9TRu/VGVUrp2Y7Arobxiw9p/eIe6hVitxbQptduF5Wj9w1mGS6KYI3Ndaqzpl9amMkI
MJT+a3nYj/FeFBfSCtf9MCXbyqjUNbA25u2vuFMioXjVhIX+3ViGLxJLrqYE32IpV5GBFIC0NBF7
+Q7rGNd4XoAfkXkbolgBNkyfGbs4oLNmjuURP9JKe7GNkndapkbjX07HAu+lW2KG68fW31aEiUhh
z3STGcyd/p7XJOUSrbzUaUVlKIxaxxeI5lX0rLAWAODTm9UW1k1hHZMk1ojV7Jh+8L5ZVuiU/NKW
lDqJIluT00y8/cIA55DDxaC50cF4P5EzaAnL2oF/7kG6X13wVHlcsCpMOdcWjYx8q0Ibynvcyd43
OREhWEIuAFNnNem8Gqwq+cZBeGt0XPTEhtVP8dLezZxttnh9VbPWlJ9TIsmlM/cH2eq+7ToXJkBL
FGcOVWbnbg+vKLZvsZxjE0YwOGa6rVWbrddhyU3OYEf+H7Z3aJL9bP0CoPa+9ldcBRlpm7/nDMXs
1ExO1yfFYuvjZLKBHAeHls7fHNfWcyjSuok/roogI/zxMC8BLvb6bnJDvvUyqJjMueURFlc+Y/dd
lg1qS/Eq3BckpOfkdF9DlzetmAezMiS5F0AkB9sWmvRyM5lOQXHakRuKZpmDyGRcXNHlCAoo6FX7
PXOz6bdUnvm2rd8PGozNUn8WfmUVq88cGPE0NyszSu2iYP6Ttef6guaiBcKqwrrIxlS8/+U9hAQj
R27UVoowEPptwCMbYbOmXYTKEV3zqfpH1FQVdaE0EHclx/9jdG3ydS9Dn79aC10Wkk+eGg/ZIkQG
z7YyHxlLgzkPfRQtP16a6HZpiVw0Tw9G7LWlF1istp4lVmirGVR1T3DNfJYdl4woMpUVx7wcYoIt
ZUxp74sXu75yFuEBa7zkpsRum7+7NSV/U1kC8uhiB40ZFA02xxYx1HMLV2uKWeII80N1QKvqHNuo
4zRRXfWMkT5WESSftq84aoIRJnz5eepGucCAw/AxUQQb5pwawpIQ5nB8yzO/LMPbfCCiGg5WYSSw
kLLwRRtl1tX0YzuQsfv6yn4lZxwmoDTyJpqw/LbgeozYww0xJtqRlilJWQKLLteeEzo5Rknj6XCu
T+zwxCHSOu4qPnal1gyeE00X3sKCz0sTwHx2pvj1rDU+jkXn74ZST5ueRkCS8V3EYNYf/BiLcHYC
VPgUnbUxwfLdGQ1tH7QEJpAEvtROSQjOE+lz7CVfDDZraImdrYQg9J3W4DaLmbnTseSuEskmPHQ0
Neneq+MOMaYNajiNQ0vxSYJz9MoUiwrsChawgCP3aMKmgb7Jo9tmqqQTLLBy1QQ2bOGYAcNja9Q1
cRPE37NYLfVCIqeiP46XdlwlvgYodOb7J48NvADRjpfgvwuXpt18zndhr17yWlRk7THRpQTa9Ggg
yVWgyJbJ+qRIeUN/mfrzfE5Mo+NjmKQOCT02R6ecWy+XLUsTBGmeSsEuHqhPnbJCP5kl4IGr1Xpk
oiZwi/CJ/uOrrb96eSbQi4aAXV5Y4YpublNSuV4Eb33d8EECjOyAej6mscupDix5E/HSEvkPbrKs
KnOzUNVyWoYVU2c26+2cNje9+t30ksC8qBYTuOy2oO+2qfG1fqfdCOqYVPZAZlxlUC0mTPl9Qvnb
6GsVDFUtOzq1YDci2P50vHhhj0oIHPjPc3FMkdrGbpMAX8IAb2pHBbinsl74YhjDec8yGeiIov5u
5TsLLvgDCGqcvCRtjHZ7AS230d081f04Qe7Kds4fxhgfdJRirRvScPXUJzQ5GWZMuoAHEHM9MIui
7Or/7U4KMNi5ow5eVvV+nlQjGeO3ARB2oK/f8h+pa0nZkm41O1jyc18bvdkaoz6oULUNJphdL0EC
j+Zx+otLBCND1+fagqtCcksb9rf2uYdq0TzP4AXsL/FnKw+9Hmu4yWMR0U1Y+kLBSy0yDe91eBPA
jkHvq2jzVaij23o33dbb+X3I5fJRiSgVfIaUu7NJci3yrUMPzvr12j8MEJ4DjOkayAtjwZg9WMT1
IQXC9DAvvtta0foZWoQLfA2IaFR1IcB2kYup/94kgcrcRvXZLYDP8rUBVSoGRMxLVmjI6I/8/Es1
pY49wULZHN9Dw21CT0dnJFK7z6mqOGzoUGVwtNyZws93TGOB3X1NREkYwJpwNjfzNwHenkLKjnKG
Z2MVZYeF7S/ZQ7aoZnHkkasMBtRFJgyUl9jcvyERMGpM35s2Sa/hrQifFkis/STZ/j0J3hmQyn0g
pYMNi/g141/chCBn3qGl7RoTyuMBJGOyl7o9flmToKbHVy6fgE/284NKJStZokg/ZygfSn2wV6G6
G7+3BeCfBdpGlCEgzqBpO2P9rlhFmxO8a+dRB63Rbim4o8q8R0q/Yi2nzM7P7wQH8K1JeswrRcm1
pQOOW+8aeINQCuSTlAPPOghpA+C8L/96fvgeYSsxiFaa2+Haoz5JGLYuTOnsNe+6AWWvu9pgLKgP
6KNJFD7PxOzSQOGrJ9y24gEo79tSYBs9eniRd6rIz4Df7TSTmv0wJ+OOHqm0aRpmf7YfELhvAQwt
vCPwnM+KlD45kwu/6Du8x1bvg2pZQpFr+zN17ueDchhKSg7pC3sS7WbZDeHYGltl1HBZcbfRL1la
KomiWRtvLZpuVVywflxP1dQWcaISGbNI7MJ5jDXPqXZiM4RiImKxWidvqoqrqubulnboIAObxBjV
bLw9GfxcHSU+o6x3SaVRSENrGeTOV4+2vDH1o4lP3m2gSaNmANMw3PkDiZzmEvfSIv3g/6U2vqPD
ZK1rnWauDgy7TnM1NMe8KtsXEpkqTNmFNAPwNC3Z0ePpEdM9t+pIr1ZRV1lSEL2c53uYEj0k7Lur
j7rGlUGty/sEWNr9cDCQxdCX12ntlA28vDmCU99S0QYBoggpC4/imAsC20Khq/0sbIkPRO9S0AEl
Bz+XTPttw0z+g4UzMQiuHJyAWTlJ1mNbFyabmwuBt/JQTikT/gKwbBJWDnAIRsWM7rgOGzUjSfmm
dTKdzzwKT85qgQUZ+ST6lBFd0OaA3ctWKp1Ie9qoVLSGPHEAyeT0u1Fm5Aaa9Chmw0+vR8ZpdnR4
ycrREaLQItHoWQ1LudOBpN1pvueuvrR+KcTnGKTLBwK8QqWtt9VC8vaedI0ZVIQncDU+lfCpxR1T
YVzwCgAPMIg7ns5JdoXDed5Wx34HT3qFRtAeJuVewu1gnk9OJOmFdlmUWQitYS/W35YYHHhC9wMI
b+4VTcU+iF+TSRH/luqFf08j+ZH/E4hRqzCTYwBMJkkWVxHPghatzI8kDMzBde6/nkV8VXHa67/+
B7ICLg5JQIg3u06WWOnF5Ob9X+HLLy414Uai+kl53nailC5zGkUDU35RbE+Q+u0Q4kIlop8t7g+S
meNOpGA1QlDLCV1R7L1Ds0XDqCaHNzuvnsK1DRQVqmHPQXKSpVJCUDhZnfJivkxXVlKJXCsCz5bV
gI3g2tugebyxu5i1HRXQOX5PojjXI0+p0ij5hZS0TRM2CZusU0N4Nc4sGENsj8Sezoq8MNJb7eKf
O+STdjgbsNtKULQzeafGRNVatQelfyd3H/wNRWgr8rELJXR/FdCdq4+PZl39NYbmsw/Dc3JZye5p
F0bC0Rth2HNnQ8DrVA5SUgWUBHQAKa2f1DeWdfHLgKXeYGOHitkxHdcEuQOM5FmAjac5WUJwK8yY
oaZo2HEIl3kcD2iqhvr0/9iROBqSU6A99bEuPyE7beHq0ohJY+iXy9gOPe7HufkkQU5pBSuzEM12
HkudY3uQuw4KG0kXfbJhxiNK5GUshUfCKa4jAHDrseJHURMdlAknlIb2i0lI3bpYI8CzOMobvHjO
BkSvd+i+I3KEhPoch3393Tl7zfyjM0pTaWhlyrM5DPZKV0Eu2c/OO/64PeuddrEsslL1cMq8XvoG
hoDTnfx6U60G+UejnUac4qAIutyTvLTfhq7dJnBA5IHwVjLa1MZtiHvdZvafzobFaUQOa0qr/hPO
c1OhEG4cy0/2zoFGd6nxWkRjwIICQjGZUw1oADKMxmQ9ZjF5VPXM+5FiBV/2qZAnF7OJtLvN14MH
RB+eajamUpSCDvtyPq9Qx8G+FEGic5+f/DhH9bwa/lleXIX8xywJ499ea+bkVmSRIZgjrn/ptumB
22cT+qSn1lG22ze7dsuQ6U9fYMQCZ06Py5W8fZ2MZRGm7qrjSSm3LXWapfiXbKd3Y0T3NBKddeeE
LzvxEXcJfvXEFFLWDsn2w2ZnWEfhFzkQjsoP7Pg9GmSSjMZSyget7lRsv7W/v+ULCaiuAYMOWi5/
saqvQ780ubuKGBjw0vNWFBH9H4/4tdUIo1GlX1rECrK5s4qTeOL3ARB7yCPUh2Rj93lolrQXZUb2
F3Y+3RwmGkRIZEev1FXx60u6afRdxrr8DjimsrShsmTTAuCnAYWJveQiHES13jhFkHu2rdhiKg9Q
FZmye3Pt94627WwcDtpxxU7yIz25MDwo8mTPqm/jvsGbhaF2jrpWDosRHHdfgigJP+ampPFUX8Zo
797hukSNADO1DYRFbBqPuLkWL65GADo5TpjcCVllUNHRMRiJj+wQ51a4mx/1LKrhRSXs5DnjJ7D+
iKFcyGPncVTQDwcfE3ceo3ODOxhZdJfYFIBUuMaac56ODJEELiWTsFoPy6JBPaNQTU52VqE2tyvG
uaQdT2PZp3Kn81PlFBCREuSHKqbc5hjyf9QeCxf904ULCgv2EHMV+TpE9fPfCdhfD1S/cvGGk+l1
LoexCIU1df62YpNw+U56USSUUdIP56cW/WJHdahOglPQ9TsrKMYJjUVMq7Z/l3Y+fmPWw80EQulj
hRSW4firYKR9A7fCd/MDoZG/SNbGX4+/sPl43PMtypK2gvYEa3P467BLNtuhMgYhlRatkF493k5b
SafTb+xcfRqxwoRJcBFVcRjRPNKe/8SVvRBlwBX/SEOvajvunS6IuFpakrEYVZsFuMdNv8Z2uN9/
KMilcUxfLO03996sbL7mKHaf4nY3ink6m+2P1y0yZog34fE9CYEHLFXiRwJdasAi8mI+KMF/fDD1
PThufEMvNL5krWAXA1U8btPLGQZMUe29Eokefg94XBrpTKmNaaWAQIBCCFPtBjjuTeZ0PzorOsve
NLXjJVBNT9ryqwt8D8+pbnAmqQdUjZg+5a8dYMBvOLTEtODlDTllH6OWbSxPvt7xUqHiFrkpe3OI
gNYE2ieH8eid8EMA0oMpPFdwMf5iP5QiOpilYIAq2dcAhrpANFqOJjgkKyJagy88v6oWHJMJbFyg
P1ZM0Ymv6BJkICnndG3Xf1MXQcD/4Vu+4YX9XfRUKKGC4iVts6iXEC+u4Abjlk7FxcivMk0h0G4w
Qr92lboaa9fiPdNvu8h3kIedCMgKW1G2bR32GoDTRXRcJ8UneSGWgw+6m3w6YnT/XQOZSYkZuTU5
eDK+0TFKPSuzO09tbsu29BQzP3uwlHuaow8o4JNDpRojAB2QbigDVCoAram6rcAJTARZR6K6WyDR
3ZEp7lCXxz6idACpW1YN3kw3qlp5KC+zB81EBvZAhZgfcIWEIXfgdaQVWnvAL1gJvIFoR+g/gOOu
8PF1Elbp2jAPqwUiDbqj/XE2KsB3puA1vG5nr7PZb2iymyce7RoqXnvo87ZWCR6KFXDEgqUrXqPu
pMQwIs2ZxIcbmLdqL+gSN5wwL0Tc8OjCZEdFrtLbw3Kt00RYSWVE4+yZAJ1oRltjPWuBLnogVmOX
s1jyPGxvEFUP0Nt0kKWh95Vt1wriS/AGNA2SquuZaXKkLcOB337Juv3IKVFJLbiAloAwSi9fPB32
01Q/YHGYtmkd+Q7oGUlm7Yo6bqi5fH5JiGaR5AHqnPkSM/gRwvDkBUwRK9szywo7Rd/c5p4s1c9l
ZWy86wN3q6xZHf3dGdza02SFDVi3PrdoA90TpQqZfz9t2KnxYnsbbuR6sjjk8DwO9HhLDTrWoqOR
77VzcxTB7LmrYgGzYXDStKjfrftYqyUBE/xV15OMQDMGhD6MJO4FL7jEEJ9dKHDF4m+cuK+IbN0G
FrtQa+d2oEJwFJlKVVPSh9HaxGhYtPj766ZgiYTCA9XNLEMpRk+Pnqkwif1YdOAK3gInMqD9KXtY
r8v5cJ7NZPaqVREYLsYKOGE431ZVSZGV2pbTgbEenXKMdk2KLTYU4u3Hxe1REqqykeeFmB8OROp7
i8vG29A3XSg4SEsATvmG8OiIonluCeNEA0Rtf7XOY9Xk/ATTuZxUNEBpZfmqsrxEKU/34w4LmDuR
HzoA4ad8zPNxrLbx4aQ4Uc4JVpedcRlJnlYsNmsjtY9KZmj6ZP679LBJjSfx3dkBDfdu7b+iG+/P
fZhSiVNCmm62Ym07Wi4w6bI4S3IePyaepldXDXk4naz2TobtAVbhlSR8xFmAh2AY2HOXXDsysm4x
Ty2gb0Ll1TOxC/Ij89T5QIE3SCym17NuLYcp9KUkhIo/ExLgAutnk2Oc8V5L2LuFC99leBcxVlTW
lmthJYs2zwyd4lR3z/evib4R7Zv30CVwvhFtCQhCcKPXD683Tfy35WirsZ2hIZ2xjcgBUEehJAAa
mSe4gsoPs8LtkCrPCKFOssFzof/v/Fnbq8OKxqgDHpN8DDtcTVjWDgrPSKWtqRbYuV3GZdp3Ir+r
4wL7i/STQlDQOh+eLhn2HwrEV88s4jyuj2kogM9BVvNAl8sBXjtiE8kuxBzycKGHF6NUIQ9t0KMq
f355E2p1caQeqZtYgKZDZDncbba+bb4HpMGNa/c0Jlad6T9u4QmStCU7GF0AXVBYu1AfzS0/RDCc
qrTEuTMbD/8XtpTIQArUN2B+n6SUeMpxcsu1SkaJg8sZeSsAhNDvocQZ4ppDn99WGd4QStLryD38
i40rCb4Y/+WqNSF9KX+j7wCpUiIMB6Ba6dYWDlhKRi059r6Z8sIniIcmUtL9FVzJq4dj7He+4KfM
ryCyWHxqUdExy6+K6PvMh1fu4cMLlMU7IFlar4M6kN5CdUwSuZvYw5HK49Kc5ZRdp8/WGwoKBfji
TSBPMnAmHmAh9D4zgFedFbw3F+BKFxo7bcAx0/7XyRJcu0o0+aeMqxxOUKUjHPueEqSD0X8HDTKm
vRFZzg4oTDO10T1CYdXDRsIVMlY1NPez6HjvzziuNpMSmwKvkLf9a6BBettlN/OqTI6f9BMoSmiQ
+Q4x9Vn+YzDzrIeOZKCgsh3dCkin9QIZcbih9n9ZvHNARrontcZUbgm7dLoyN8+ZNge1a7tXRNhB
t9o6jYIEjhgSKnV9JpVacQuz0euMYtYx1u7ITpCdpuKRgPVPQWcsvSULR0bR9zhyC4stkWuQcC/h
ihTrFR8tpmRBPd8r6UmBjgKlRsC2P5FmVJdRB1lWSHua4F/Hk4IeDofgTAyxdE3Af5s9XbXNGXGM
Y06fE/FTzcYQ6camufg7JL57X2J6sthLgYsdrlpjnC0HHv9FL1DQptPSpUaL8oFsng48sB8SGAbx
998ptmcCfyXR9gXoyY0Q2fDTOmCddqv80pIEnDLh1K2J8Ke5VlTMqfKIjq+RUOmSqdUd/TQU0TbU
w9qLEXwA36skBk9K70ron3zyl4NMhFF9jWx715mbHMRTlUfFZYt/lW7Cye5Fl4lH78mZAVWhs9Aw
sLtDeaqAz4hDS5a2W+9RIEGNPX6/oql3a+N4LpHkxeqEunPv/faWARjyPoez3LtQQ8lK4dhzgfSq
ixifwQ9GWr0cwelnrMYIyk7sGolAJEIfiqpdhm1qDM9F+0sBVMQjAH5YcvZW63ya7cjLmfIScJ1y
LF54erwA2wiaCggzuIZ/E69oWRQJQzSZTsn7BG2+1vL28PfDcftDE3OnMJ57oN3/ZIY4i/NQmgQj
rU2riKtP3nWu/dZQtzP3CqxH70Z1NYfdwxF83ziEMAG+6X6nGD4A8zuwjVybAP7siGe8n9oSJwTq
aZ2xdR0eBPvS7z41EfKwwO9fX35oOkQIFz1gJaHBfqs3U4/oIAq5hyTblku8CPE8mNZzKZXU8yPM
9l8iWJPt6OKbBzZcGAYdymn9meDqe2lC9lMN91daNJBlNj5FQe+Du+u0I/xii++yLjzKJS6hyxhN
z7JuoXEDPM656mKQtbbz7azXuj3TJam4bcNw1FASwFGxsA6O1AqWJbbLiWhv4kIOOGsF8oLgEd0t
6F1ySTplUwzzngQ85rnKkgIeNxPDxSpSfmyNRvZXfYuJpIR99i3ctqSuqwiVMeqYldtIlFH73t0c
t8NY4w+BXBZCD81FQv8x/21pI0JivyskQulYLWO2hqPf86UrZCe+OGcXCjLjJObmPnjeAlPc0+c2
s8u96JkuU9Zzf/nAPRNrYwAIP9wUK/iySn9YIdMD+FKc7XKtbRujwUnNa9qewTRiSv+qZb7V6Y/O
B78hHnwL4N72rQStiZAzOgSnCshhK3szR2rWQP2Pen+RFkGENJTzkmB9fOX97q9BRhW7uxgpQQ0l
XlaqGHoJnnG6Tm3r29cWpGUXKDQCY8G+8+4hgJJJN0zYJQJ4XXgzeeKISZMuJB6DZr2YPwEznZaU
fjhXCQMjtkvU/g4kWitNMCoJgZDnoiFMykZq9nFvuSnxvi/yy/RLXFZEY2g1m0s/TEMP5SonIrk1
ByKOQD+yVfvS/WKsiA747FFPuqkxltGHVTpOtxFY6jZlALXT+MdAxu6ZlpsNiTlblr6SsmA4NFno
S2vYI6xqlATmm4VOHCAoFWInnNTRIcLWd66VcaSZduQkaYbkrjVK4Jl25dmEFpkdszh/Qss4eOsr
wLuKlMZZH2ylOoDlAC2BlHx17KAEEioMpmKBC0z76H1Ue7QgYLZrkRg4ZU5OUTEM8KqU7wtkXLRp
Zid2Qv65kH+OlTV38J7CJWMS6Y2SENxKaLolYXP62E0yMmitVVnLBRN0h0zeLDs80I9q2jHAiLyg
0zlVmDP4oYlkChbC+vcWWnbPEjXgEesCj6L/rYPtXik2kiQHPFv27uNG9lU3tN/yoybBQYF2YfgH
NBwDGFBi7qfPGalJYkgMLEI/FsDNhGjJ/9AP+kYZL55/apGInIiwBGsYE0VessVZYLK3Zxd92Lro
FtqtmjZ/MqXdYsaj7+xVS61+JWXsIzLfTQ/j5iu9RyLcwLsdR1yF62V98MPrQzpPClbJ/nGkURC3
K51TcHI3f9PGH46FuyF5ocgLpxBmySsQup7eV6fa1MLOXpbz3UkIcaS5Qp7Ryfm6zYf/ILFCLJ7w
HhFURVWH3WjRestHOjOQYiaNtGtaCmgfZDgW7HZBUTKgefKYAEPb4mkMPyedE+gaAlBiiaE+XkHS
nSELRQK2H+fIVWDq3iU0S8onpFmct2N4epB9eTVErAKN+ESqnmMAJIXe3mLMfRiS0QBAH6HpjNxO
l9Wy2qmh0UpBz3kcfBT86cOp60KaH/HoeOOk5EZs1Fd6DemHesdUltBZ4RSFGSglUSWMtW9Z0wu5
daq9m7FtCU1EfcfeKjG4NSjgBQVhNnshwYBvkJ8r9/c9ec45lRWU93ptDN0s2lusJCIHLCt4g51B
w2UhMgoqh9DJ6zYrDtyFVxF2rd7MvVTPiXcJC9J6yKeFf4/9GCkyuuo98WzH/XGXbU3/B4b+Xa6/
RZZ7kiL64ySjTPBFKSGjI/PQo4Ne5Et2NjngBcwj+sWPEwcfBJb9Pt7RlInXI2dgjav8DlVgXOwW
CkybruFPaayOl8tw02ZQ02ujS+pdYVjKm31pepwcOsPtFJP7bvPuh2SSMj1OgjwTacG7w0wLNn6S
0dVCdgBrHidocueKGhcrrDti6N196rzfg9AB4sW1AmsBnlR4sDXH+NMVRFga4j/kRASh2haOCygn
5EF5TtIsq11r+b485sN5t+dbISuvqbRSi6LJG8jhmspVxL8Caw9IvV2pTxSrYjz0Go3rJeAm2cR9
DaZiYIqWg5GkrhPJpQLLR1yyZcOfKIJoooKlCWuuCTEujUDQDqZZVpCHDiPg2H5mBZkidX58Kzjo
dAKugfypwqO3b97BBCm8ZzXrGGqxqjGFVlUxPeTJS+wO3IbqdSfkT62j0s7hqOTmLuz9UtcG+CUf
AKbtx9tuZhNHzLojrLNRxykz0Qu7dcVeJaEpv8h1wq9C1pSDyeCiXmhPdXYNT2fdulnryn/7e2tz
VvPZyPCeNb9vCrK79B7PP2xWkOajojxGp5XuLqPnt4c8zdUL0aB/IIM29/X8l+XqQs+LYM8Rsh69
01HxaynkZEpP/4cS23TfQxeKu4Vqdx+sPNbsiv9xqu/j9Jrnqt6Ir6nkDYORgAPfSJf/DIKff/TS
/upAevpAPm6STRSxAwuJol/ZjaCSHsw2BHA+bSeRe7/MRJjiayHCP8BNxUcfvwLZ6u6DB4JTWgpz
pOH87YPpyjHw+2QRxYiYfkkDP4XHOI8X24LhIYRWLz2O3Oyg3wkukmaBSkl75InPSSe04hh3/4nr
I8EH/oN+mBTC9BJ14Glv/M9pEkGkFj4rX9IuViLzYYzVzW8XLqxsoe9n3FeK+9/peR0uBKcSqi2U
f/2w9eAc1WWWMHOkqnp4J1qFpfONhNIb9/iMdlBl4LR8uEbalEOSlT6ROD0AU/TCGyKpmIyEWx9k
vj2BdQzp/TLxfDPybHmdoNhniig40knpCQzhziEJHU3cm2OIs5TSPXhSxDVgH1TpJS+pPN8XoYN2
cSNKot3MM5OQknGfkBBmdoyDRP4ThNxsJk5rZVdrn4bfQNcZ5eN8gcdJ3qbZ/fT5cz0TTuNh+bsZ
1jdN5LVNp6oKz8T2DgEp3b/9gNlT5rxpVKpbfuqIbeRP8Dw84kdfy86f0L7tGDTZfK85VlRl4vkA
Pgz/Awfvww7yqOze/LpjtFTHuud2kDgerIwJ7lYYJnKAm4q0oXvWw6Gn4CuEO348/Fi3Ab6sC8Yh
FRRXg3i9Pt8lSj1rn3Qdo4qaQO4FpblLoYlFOFr8UEtcHGauRioz7gv1uorEGu/uCk+HFub71qQf
OvQmrpcbYO4RIPrJizAdogjB2CNDG2dOrby+5Ixw6P2ldKKK219bN1ZbufFiM6Sa3q01vacvVeh1
w2X0AumB0njruPhKfYrWpIyXDIkcyyPSx5mSCA+G3UV4DgpBMmkiksFfZr//n9TpExqqIzclnqne
myhyh3cLDYP9iwNWZmejX4HTTqspwaX53fZcueuH8fFn+W9Q+bE9pTfvEvl7n/jrB5G+fhTUaao5
9shdKgC0MkxAvRpLNpfpsgfpeYGNYLq8Lc3G7J5m7JUWpGFdYBqo5WzhqIQj+nTjoBnCD1rr55T3
KK7RZtEwNrdBBOBivaj748+iOsOkKThyaeUpaOh/IfQH2KOk4QotnhnI16ZlfVyT/ZNKpUvAYmoU
eNgG8suBpdS6Vn7YC6eSJfRIbGdHykDcwFbOiuotOF8+2damwA79mTFs1wR+xJMlB+dAh/vMBGCR
KLVu8qc1cpLml7SvIplpOl02lbaT2hqXL8Ywu7LnmAmi7UC96iKmTOcZXBZeK8AdhdwRnRo+Ryuf
QceCG8Mh7CSUbspNTXObVH4LcM6qsO+8OrOTXGzNN2UQPQseC33WbutK/jgv3ogszCw5ohQTloO3
ZWB6pD2x4rP0Birrzlq91zhPj+ojwgSMPoqjtVADyK9UHj0i8F8dL1YNwdJdmvSr7PkyqHZpgAGG
V0ywMD3oaBoGs9eMEzefmPWhlF9NBIEZHVZC7ePcIhAVzVhBgNr6Hqs6+UGOzbUsc2oyjy1Fg6Uq
x4KnHAQKGj+UEnm0GgcBOifjClAmwQP5yTxE1t5WmKlrSsYhTDoL+CiKew5OmpW6NQa+aIl6gvfF
tPE4zEA1iMXM+ihnstUo0s8a4K8zRbIeAJOZaJdKjttgc/4H6bNN9BInDzFJfJZFv9jcuY5Yl4X2
CHMw52CVDZIng95j/StgJOZJt129QA/X3EySRE5Gukyv+dAvj61xtXRJARmMbbpj4d+xAQw2mu6L
Tum4SQeoiGPYNHOstSuMdp0F2HiUNRnXigku6/rtXRIAIkKddvbqwPI60Y6RtwkfSRKt9JJK1/Z8
BYjMbjp+uFvBKJqXopKQk1LC7mqSk0MenG6XrX8GcpjPV0X226ImUUwWrnGXheFEoYZmQafklX48
tOQhT2wqRm2gWnsczx/QIwnqQlf1wTI9XdNa8rin6IbrvGJEot11G7okePg+g1zG4iy6aBFFpdD6
wPkQVKT7prL9UjCu6Qf3Oci3JlfxMx6od2lko9Ee5ESxFJh1aOIYmV1mfrROgjFXeLsLmWn4duGq
e5qkqgaca/9y4AAepybt9V6JD8QaJzjZsbbS9l8NpOjSRGONAPu5+OYa5KAumoHNuCEE+WRdKHXC
yZxSzzuoHkcT5Y57wD1MiPMImfifQ0SN5QUjmSvCKnpYHaK4uGvYEpknTl99PZblinRESnB6+KTH
QteiHOnXMPRAnNqQZmOm8tpCTSNvAngDvqvrR7Lm7nu+AV5QbkshaRqjpcXBWSm8ge4ESekR4NVI
lnFDgCmnnF4S8X/FSfBweII4OG0nkGvoVOkZtDKp8mLNcctporbyYAzNq9Ndlgq7OyLsnfNqnmLl
EHpCrICZk1veNXGyg50dKxTn90wCkMjIvU93JJnoyezUOKtJkyTu5VCPL9oDTvRDa1RH52vWGPE5
0qhqsnspWVaazv/S9snzDqR21FK3E3+B0HhPXyFhwZf8kV0obbSoxwfCXN0Hw7nbm8ecqCglo5FY
Ld9ksu7LIl7o0qsrroGFch6s9CQs92iJfWb7DMuwQtzNEE3wDR7b2kkKD2CwVP2f5Pj6vAhJkWix
3MEdZT/D7m1vVZ11bb3Ii8lA5hPHRtTTyXdasSwm1F9VUNWNpHFPY/GGs08+pNGITtxUSDFSuEzm
fnB3o2ILX5rNEVKQGlvWHxNLWiPAKWzkV+ykFIHF3faC0lGEHdzG9Qj3R44xALLqRmjhqGbUKskl
sBQqw4Jr9Usevzgcjj4TNFBlpPkjTk779JUkp23N9KkxkEWvewVFKkt6MLrYAsO22rrELwFfhqj1
//L87+wAxbc8fm7DEG5NrFonExZkeoFw7q7cQWGNPh7VbWPuqMjHUnl46caanh3Kc1mJJ9ZxOuJJ
KqnYC623RpHlS67voXcm4pmEQiSz7WtO63uInaMynhQhMMUww7F7tm+RPqV0CIzUjIC3ygQnjjo+
UxLPTaAI34p6Zzmv6MbuJc4TK4hP2NH9KMLyTtTVHO7fMDZaBBE0DodwOKZ9G/roEBJ4uoEAkwEy
lJPP2Jfxtlj4AJrBL7uuAOaGZ3y63+vl37YSar5Goc/hp7dC9DH00Kx9AklPewLkgpi/DgGr9ca4
UmeY3nJac73sW8OPCV08b/4Rt+iRW9jQXPmG3tz8ipxWaX3TVa2s1KtrwjjN2rXwFbt5Fg6zcGrZ
DoN78KD1O3kcqw3XDhVA6NOVQY9Swrdmy5ak2AmM9YvgO6UPLtaFeZqNs3AFksJyHS2ypx/mOyA5
wJmi9LvRD14I6jJiXGnwkLEOio0I1KfuAq1RrOpLtkysKq8yer8O0eVGigVvpTRGUT1dGEaxNWGo
HmmtvrQSF1RgGCaPR4l0Inh9oPLiAm7YOg63Pw+5YOwzNhnrsgc8A3Q1yQoo7r/+ci72XYU/E/AQ
8CRkTd6CgarT/2JZzzURMXvBS/U6SVZLNnhPvUO0s98iHcEhM1Jy/VITLXfg6wCkhJEj1X5h9HiS
g9UkwdZTNCfgRtLrJUcnT0EjgkKCtxXN0lknUPr5CGMT5ImeApyRgRMQhbzeTYJtLjMzqd5GPTyi
FRQZ5Q1lv6QLjQMV4RAQxx+otBAEsGbK+SkU4BoaTTWfVZ0ncV9xU2K5XzxstOSx0+AgpRW5y1UB
DquNcJkNF1w5KOEPNd9ctf7d1j91YsLU1RvZApkU0BdAGG9roLjx8EVivqEBY54f62H9sJlI2/4Y
vfos+s+fNdJEOrilNDK2P2OLyOR3GX7FMaoMsOmKhu5BwL3aI5RJmsOV7VtQ60tapMYYXvHVxdCl
tlLoa3cP6jBjC0wqhUd2/1WDIfBDlMgOMEN/Kr5xa47tBoNC71ckvgiSCPWDGQSwQY7ssBa5TU0C
+deXuvK/vP/MXs3Pff5ppZB+1myH+xFPO41ARWdd7gR66EUDT84QS4fT0KU18HYoCQaDdUjBnfNo
dcpFwLa6VOBBcNXaKrbDAZquqx65pR9rvlqAd2QBXMF15myOMHYJ8FudEBbxcqMUy8UIBFlPmBDw
qtt7pGgF24b9rxzb4Q+RQSlnAaLtE4J6An8JUq6Q9+cq0diJ3VgGll6s+0uf/qhE0ffT3twn+fwU
r8BCL8HV5LvIeLZx17I1LovkxENSb2c+11YaiyJQFzg5oY77Ck6kn6KdJv5MNoHIV6xNbICkWyHB
FuRaIe57Zi8B9HW/oekS/ckQo+nZTJ/9vDJ9S3olEfevuKsH4t2+8yLNF1rA+md5PuPa8XpM/fCF
g1aTpkqZ8I7ARWM/mWzLjL8E/Egubnt21o8stjZQ1yLCG6d89yYiVCrqQ1QSkIbBV0qloZyI5dFr
f2GNdcezNarafNl0CP3aSB3m6YMz/zG7uysNLcMHsjUcXClVIXm1eIwsOrCsEX/229oKAUCUpqUi
VrKwu3iRvBoXOVJLSY1+ELBFrcaBS+Kx5FejJ6gw8bSfFWZsHOJ3/161rfJ+nv+ID6dx+pz9VQUs
hmt079EPUJMRyZBFv0bMpo8w2qw7Panpg0l2uO4Og5w4cKCMRwOYmF8WaJFvgF8gE1yIg+2oOhPD
1kL+vdcGS/w4IN59uDWqlj0OuIvdwbZpa28q/9juV883SFk5QPIU5X8RJi1F4TqNVk5xVUf09Xy+
mATz6QQQNh7l1jsefleBWUwVRs70WlDOq0Tn/5XfQegSQ6b7BebfaTMuJRS4Li2sjuvgsRSd4v8h
hvRYpl54PPso5A9bHw/W/7ObT7VK3xU/0+so/ewf6tiVkdLXjpOUISqfE7rpOZj4uATbaAFHWfg6
852rNstpp051CqOdOkJtatJVVMlErRY30IhICNJUyUAdI5842XzP7SCfnwQy/etwTOK2i2s25i/4
O5zJrroBh3irsM8/7sHDJOUPY+IJEbTG8JHB+JnR9OGG/xJ4tf7pDgrK5KZGqBuiLcvq4Q6QQ4ic
ox507eUO7Ql/uPDnuiTzBjEeppLZn1xqAQSq7mNL0POGQ+Z5tNXTVcbaDLH5ToD+sfprN6nlKLC1
nVrJZO7mrow8f5FGeLcUzthi+SkRib1JxHZRXipCGphshLy5+vhcb+OXNKeEHZVqpU4TGugLEOZQ
Zod53dUvduHheDxTQExxkbiU2zh7g1ufv9PxRspwW+SBQqLyHF0DRub9l/mgB1olWKIrkulsewMU
1AhfHFX7L0aH4E/TJyQu8bYlHzjpi8Gd95S/MoR3OywTrvzV47qNzwRqNuVpkJr5RDiQ2PfSQ+qd
vConyGU8j4v53Xmwwi4MMPqTij3Alfp3OvLAeEaBzMW0TPS+U3lOODnC0mYMnvp7SLtyURAdhX7e
o1ywX2vQJV/ksBiFJFErbcFKmdJ2YzNsv5Er8wzReoauw4uL3hDfCv/Zuoyr0tIQNUqRuDqlE72r
q0KRiwRdRDqSAToMtebYS6HqpPV7rZWwhcSDVQaP+kldjy+PBTTt+kSnlx230lo6I60gmt36J+2x
sKnR6Rk0Xj7c4IE0ZtT1iX3WN2jlcjGZCRI2ljzJkr8Nv8VU+/A9CroP42z68CacEDLOk9Sbax9F
rUxwzMTXJNmoFm9F/eDv+nUTRld0xipyfRmq3tq2E3fo8Md75wNFTc1gP2Bu4LkqfuGlCaNFcUIX
U2xQU/GdYJeCBzTqg4Uc+e/CUa1uNT6l+6YO2jVTWu4DBDTmNNaVQI1GvJ4XmtGdJDLfwFiBk9BH
9DVbn9u/opTGDDhL5bSQh9S6nVCObO6nNuqWxVcUTH3SKh76r6UukAAR6qFgp3LGzFQ5BqnGzhy3
odJPXINwVOHkMdRwHKDQL2fSeJMnoZedwCFifhxczKwLntivvxkqqU9fB9yIZSG/5AJNct7fCuvv
YZUabHhFBOJllnZWyja7B5w/2UGA1oQ5BofsMP4wFlOP/FixjfP/E5d4s95cyH/lZEojKqxsC2RB
iUX/t04Aa5YbzfFdjA7ZQQGNrj1+KYnRoUqGhutdom0SBlb3FZasgeW1r9BVy6azYbIpQwWzRlLe
dnI+TZGezhAKIwBKs9RCI5uz1PyZscqgH5AZYU3VpSKQaAIxaspTyNDZM38voS8Mawoe8HXEcoGl
V+Iho260K5ri6iW9vPMoBnf4tWri/ioF7nh0FMCUTptIpEKH3eS1XM5UUf1dtLBI6Ra2KD/JFZ6M
200OKFPnwDKOiZwDYtH6uXpt9/r/WBvQHetgmRcfKFBV4bHcHUPJY/DApK8gs8dsT9IwwjTy14wq
UYQ+A5wDeWX4V6QX3BWhxF6opfHQHMhW2pmeinQFvghM1Ujo7Ou/g+ettMiXDRTYI3XXCe4eRhyp
wnOCXHrxyGpr8SexLcciDvSUeINXUaEEIVYiYJtN9HwP9v+g1NYt8LJkVB44fudyc9BLKwluLexY
7dTkmit7fi9kIPlSQtADBjoO8XyzsasRmzOlBfv4wvEbDOz0iErNkPqGegPZkxboJtDupRgzhL+C
cVHZiLkLOzyWAoEUL8en7vat9klPxeO1AZ6BRfBZZwgUaVwzQea/64Es5oVImCLOkoTFd3k0lp6Z
/y/WTUJLOD1BnWE+nfUMw87mdkVs6Za2nNw0cIyUaNPhWLSZgPW9EyT6C/Td0nfJLqc1lUJ+WGKI
h+F089Fme7EkiwJigpJohrvZtF3Fv8EXbTjYOjD8phEUDX8yp6pf/tkXxkm3EjBRgeda2NeUNyc+
bQPNKH4qY+QIlfvqRluQH+gbw2dva+3ctu8PKcsUEJ0ccM5/kt8vAFevOfOXuhe/ojdtsrUK3LGM
5w07Fj5vef3/xp+4A3nsYvZxCu8S2Ijte+X7B54unl32AvtgmfUrJynbVXrYvgAA9ncaDtBjuzSY
lBx/BDSLaftcDjuYLGtN4AhcjAK5AFrkOCtD4dJJgYuiqNTJG84olafFhYIO4t1tVgefSe8THsP3
bMO1tqOXz2WKgGUHsxunCWKtN+G4Jfl5zjEGnGl098h/21ORZbTdzPpMZwUeh3ovl9KKO/DwTvxo
HzsMHQrSBIGrDZ2AmL9dUaYaKTQo61c4ZxEY1GYbGhz2DO3hqL6RSZOi9IxNnYfek/TFtlRfjh2X
qYxW04wVJhf+jQ+XkGDRKKRAG6AJbmfzyDY8fLn4fQP2tawumX3hxYruydeKHUNFCXpMijDd5P3t
VzyZ+l+duS4xSz0ziKKlKl8Cc/xieZKccSxPxEnzJXyItY4xhn0EQ8ouMAevTUyt02AHSbruOhZa
8KIqaOkHfqCLqP03L86mdQv+8mfhymiYePd6a9SnhQCaAhf07I4PcvEKE8PSOK29594gMS5c5ew3
VRKMh+A50O0WF+PSyJ4esdj4k9kvw0JI+9mRnP5AVBTIzCohRNQKXJQ1QQwHnxA86o1LqP5E4TRi
sSdbn/WLLT/tRx0QOLNEc0wwvVPtT6tWNWHhkCFjdrtAVPkk1cUN7dcj0q6LghXxBfl1n2Q0FKR9
2QnkWtomu8UKDkU502WxuIXxV1Lk6aeDxV+J9gPlpC7wBNGgb4Dx31yB0xbG0qP1Kcdbpw/p97CA
5BeUstdr/jye6S8Q0lGxRc6OWBrAZxI9/UtsOjev1FMbHpsEpogpBlu6RPhS4kb9A1BjHdFGY8WV
OU2mU5OTl46xBSgC82KjZDLOu8kzw3f8t1PrciA2r6PGaDjYUwW15KXYC/J8Ant/8I06AfLIogC4
OKMbHMesLJNgez3MqHTfT5g3R3d05EN9oShHSNE2aOM2ekRZfMeEfJGMz1A4XDZuZ1wXzeohTjyZ
O4fR6qCGN6Hy6jFMdJ0GdfQWovDO2rRl4OyQjiYr2TOMh/7v/pBzozXCTtDToEv49NI5dHLLBKgY
tZ160TXeP14BWqBx//AmcJU/RaWVOBiENYM5dEE4vxx6r7avEerRPsR+hrAvA2xZE6qHGEgIVXWw
RyAjtcLhE+oKKTzx8CVi7w67FOEyeLKBDQI0sWMp7om5E7d1lO7sdpGhtqovBGBVSZDlyzQ7QYxS
6agxTruGJVXFl247vMmJfHv3U81MVCCMi7d/k8/kUh9VttqQkZ5QbwV6MCRWRh9F/A0FCh8eKcGZ
doqrzlUhzh1E2iCZXjwqFWtPuo0rQpMj+1fXURjt7fRHmq34rXumyJ5hoEpjjSEo9oNcPSee3h/B
5i/FgWELFSccfKw0CZOtQ98J53RaC7XyaOlDkzG29RtRgD4z/fbufC843KOHR0VQao5rWPlSn1of
tnmxRAzXsKTAs6o28qQhxrMBDIzwVlTIAN8ta/DG20eCMf0sMNtpPBox4k0klMfyyrEeG6fvqOWP
MXyRZuL7zIIQdKuvk+ZS/4SWT17yErQ2gmXnzBcR6oh/zDgv70gO0xcbkJGwOn0HmfFXQtDN9Kfg
8boPaoNDbQGxn5J8Jcz6ZTxuFsLB/CqnWlt3HX0GewAzwfw1kuYfH5b5lEJ22+ANpq5G2Ymi1SKQ
KZpsdTto3ZWnCCE3rp1gegZ5fychDHK9tyUGgDN0G9mh61v+AjUIGkNl88beAIbMj34TKVgXZRPt
vu76IzZXUpT0B/4r8vEn16sWJR7WcUQA/8xsFBogl9qmRM/aeIypakiWkx2PU5vQ6N4fuiLwJHB9
PhP0RHeEv+K1ohBNUTx1zlVyiYRTvKK3NhsbOtB8NYfRFnKvWjHpF9LCQGTKvcseq6uvIfJQqOtc
obeUvwx19PPweE++p7rXvTd82Y7I4YBofT9E89on8jvNculCSh8Won7HwlbyHATYrbNTycTh3wXF
4mlRVdudlQ+ozF8qW4PNgpaktpwyARrs1M6VWp7TzoGeVe+w/eWWQu9B6/W6V99IDeg4iwMe3QSU
BvaloEToQM2M87qdDHB7v+JCMtjyUQk/62dainnys5Bv8376F7IW6UbOIbf4lQhKDUI7Z84OMbND
OsRk+Vt3m7GvUODqgYSURBQlEEOedwPqfQ5tK/lMmwyJkTo9hV9srY1Eql1GFW7TVItwKG3+z2q4
J1sESBaz/+dQoTJLxPrSvTeNhxKrf3R36H3cGOFgmC3qetdPgaopFs4mMvKtEKdW6fuHbp2dxDXf
RO+NsOg+4eRNsNtp2Ui+nFirZfivXZKMeJM8LADD1FJPp/fnBTpvE3R0cJoZvQ+y0lZDcut8EMZU
FskR4ohHhw6l5zFUrmZlQiSCDBXIqwcqDWsu+njJfbBcnVI+PLMPb2arfM4HgHRXpC7P2bEQjW1E
gLowCtOZ0f7SnrGE4kwqpoU8Z3B/ZYq3vCSDw6uSDh0vBJNPgde8K3jg1D1AbGTlSIXPJywjhrKv
9OHjjIcyOhG0ZF/yAaf7NRz+Bu7TI7QlG6efovHClncLKRYh8aEIgKEAX4SdHTfgqfok6L4y/1/K
4Q7OBDW23L23jPo4NzbZOaHeASVse3tvU7quusxisIdHkLwEu0wER6GXv7MJWla5nNknuaOs2fjW
uvtgYsyKfc/6f0h/StC4dYuyDEoZS2iBWymLWxVsLsdfmaFJYPCbeaEfqIme0sYMHWmPuBXeieUs
Ui0V1hiRW5lwnSB9+FJ/iUh7Vdupvt7dG4cO18vKVLJL7IGyWa41Zc2dwV2wYasRZjGMnzKoSc+o
6dBV8IPE0JYt9jIcc3xNONpGrYHej67mWaR0703bP53pp1g2heJyPt53w/bSX4JzUDWzzaqt7PHk
E8K4ASlqHXuqo6O4HwyrbdJJfSYaXct7yus2zZgjyBbF4U9zyOSweX5KurbtvVFkJEqwnoKW0mKE
/tvp1clHOAiICYxDkNNd2i7RD3uR1PzfKyJYDTPmzWkdIPHwGX/PqIj7HBY6ackli+EP/Xczj5J7
Lmx7FuJeurAKYWwRlP4BT52uPTf9karIWjypidXgbKPsYmVNfRUnR7F+2s0XkNdwn+x7JOveizi3
tkZTjB8qjfUvA7Y3Ruk4ZKkbKy1OQV4r+lKXQfNtuHbkH30+afvTHDP0/VFwoV6GWGSytEvtVihZ
8ae73/PoSLnuqA2u5YnPze7+HWlVyxtT9TIkysfrQvirdH0bzw11ANUOl88zOsujtUnzlXOueV25
7YRrurhVh9IbXF26MKw5tCM0x2c7y0JxZgFq8aTsHsBfGbsJgDWfhi+naVJodL3dqPf+ieBHVg05
RywDgjbdBExJuuzlxMEGrZPMisXT4ObZZYt1loGnRD8Sxhwb0xNyFmder8p9BQpmconDs/Od7Jjs
M7bo09nvF620/2U3ntZu1oUZtBPYIWgOWtQebQQLSPAKqGgRU+tRs6U5C8G5yQ9GyB/irVM9RJ3D
zoadeRnjNjAzKmy2bUAbZTBQ0cFy7k5lApyxWwzd5hqRDGT/MObOcbvx+M7OB4/S36DPHkSHV4Po
8iRBo8yx4jKW3T2taOIqDP/U2Kd/EhUkHGgnMM1mR0DRcNURsJiwBY3FOjo1cT+k4jd9VOznnrkh
bOkhKOFHIaHWqEkgIBXccIsnQQgwfIPtsYqPEURyM5Kjtyq8DqHUZwODsK5GHChKF3bcU5XZwbSG
pwyoXvAw7OQtg4d9UZV70C/s1XRysT8IqnaMJcYY6vptw4J8IUM+/kDKinCJ1PuFy0986tUimKU6
DWBypqgAIW19LlVYxyyWdknWDX0d/a/h14EuiHplyxC46JaxfPgk7g5xumCRTFWWJX+6cwKGeldn
q45pA6g5uCxMnts2/yATO94M0WH4qOl3QSyyvChN8idvnTXV7SSYWhRedJ3jxgw/f7B0tuvwmTuI
8qxW5qwmNxgVF29dn7Zq7a3k5ZeY0b5PBMjs0U8wO59UgonmwR0eGJLbsLtBf2ikTj3zWWkEaPNc
uJ1zhMOXdWJoDw+5RcvFJroarDQd/GfvzlDJpMXDvGR3GbZJq8mlSbVeTo+EIZgL4+UzQ3hRs62n
nfYfY51pRPOtmGTHM5woUBFM+emYB1qr4F/3CDlL/pexus0x8PZbob7K+uohYUzUoN+r2dQvhMrO
GEm2R4xFhPrQhoGFpxC0cE9aDO0IJ7PEl4OWb0iBU+fZFnA+S0OjySJ8f9ONOHWmR46ccq/zuUsK
BbWLihlpZPh1DXB+bBJ57BKcWlYzDkBlyn+dTJbzWhmlNgzoMyTdty3TXxZBRPSbi1epZzKQsLzN
QI6MnIvFvHs9+mMw4z4mgOPdUdbqrh9WCV+iKgdA6+w6IItwtXaxmorqe9/cKsjJCZfx8hR4BuVV
8ShmzPF1FPZUVgYjQg+DpcHowTda/3R2rw6+q2MkrOFzJTbv+qecKWfxVMIM0tzUwlPrHa159v0j
XRgyRVOwwDqE0QnE6h+EMu1W898UxmUKRlk7yEBNFrA77opvSqQvLZJrZibHlJPIz/tl45jyV45z
4OwUS2jUs3DEUnWmV4jm6LBDzWNwyVjTRfbg2xInbFwWULs9lkunrn+q8iPQdR8/Ei4bbZqp6twj
EQB6ZRxsX68RYXQqVdbzSRRWmD+AFPKs+T59hCizYtWd6gABOs558kXOL024YfHixoC14aJH+qsm
gr6JTOP0KZSVb4DgToMTHx1NF3prXMBoqi9Pmhh9vpPc8roahnOvHbUkGXm4AMx8q94RPIkaZi6f
UcP3svk6Z89J3olx9xDCyqqhxZnWxaWt2DNL1DFQLfx5S3X87NYHcpbC6p/QvjrxXPWsM8BSv7dm
b33V/daWO1ySDLocZiHuB6QtLiulo9MQDLYwvbsIQs3o+xiVSJihZ07UjeUmH7G67/brpws7HEuk
kqFUsNhD/VwKLbkcUD8umzHUlc6RuwbRaR1WtJAILfqkBzJyCj5yz3KK/S8Qx3s/tQVbhCTB3G1z
Xwyk8pFL4nYVt9mpLtxqo4FF4uk3iBKcOE0eOXDR3ntuiWNXFWfnKJhEX5edd8GrZnMJmwohvj5e
Km9tULTIZOBSf7YTxOvSPp12XsOhwoCso1OFMA4oqbxrD2F2kO60GUAC+CP6uR0/yqw1UoVOqiVf
yjqljccf4Chs1p3r4UzBMzkD1utYrM7T2W2sbytxGJwGplN3Vytw6OftMbFrcmstM3DiMWNHqhyx
GVEJAeJU4JEJ0okNkam5k2JPpAAotBTM9R69Dg1KpvU2kIVLkw5BjJ9dBiHJY5Uhehale9ZTHZ+/
pyPKxgGqqoU0ONbyIUhQiIxrErPIFNv9CBmH0IrjQj4ZjHJXMUrQ/E8wR7/TwQh1w/Jr62LCzhh1
4eVXXyqi6ln2Gi+xIDD8LBIbEmqtvM2Qnm5zP9Sj3IoTJjX0AorW1mgQeSICYOzGv6dUKFwSMlTC
mh8GIW/NG41Ml+EuD+dEdLKyc1LcbtqXZzLFSZnnbH6RJxlPo9Fo/LqDS0+MUdQD76OwAB7dZ8yV
GS/v+stX4JuDwF4a8Mq3FGGM3KNjZhZxHK+6M5ncbpPVJ9OrgzjRZJvM+fTbBUvGT30lMaWK8Rhj
HYzq6eaO9Xn4+mqsSLPJPkDFl1FkfN39fESRW89bYApoS4xKrz7b4ZmyFNPOjzEv003Nh1/DaM4K
FcyaYCgb5b1h0gU+PvckSrjXMP0b2hmO/ARcDcqKs9mL5e0ZX5w31Mn85/r3o29qyvrrsXNTEtzi
gUkSwAUWw+s/x9k5CFyloSGYVvGvkYxnsd6nsJxRgRcz4XSyKPYB02TaRiPF3FWmpzfskXsqcWp2
WDM97q+hMUdstcOlEBAkwj+3WQygw2YSquraXGC7b3tRqUxSBjRO2wuk7eRHD1UnOlNP3IswHq/Y
+wlOeHuggyM7jNaeRDAMIqxw9wMkCWPd6oRvsW/mlyEKi9bH1w/tlDeGtktQZ64Wd722KROo/6vU
ZEYNYgJjKRa5MWXjFvTimRfuEqm+1TQDyTTXyFlE/FaH+bDdsKzQHWIcRCwUtTmKbQC4mbTgt0/H
Ri2JbD0RPzlvdcCu2JFfkFxpa2HC2qX6rNPUJWAhpkSvsNzPRkXwyIQGSMQmP8MYiDJbg/Rys+Ic
53FO2j+ZxsSirA6osn9CzuudiaBQ1OM1sGaUCjshhgzbQnI/3wFXbAmDzC2NZJK9+Ti/LkAl46xE
5K7URL1BOVxDuyzEElDU9r1FJLDEqQD/f9NtWfK204S1/5ZG4d/YiFhNfQsvC6zEJIiGbr28cMcZ
Lpzh5XRlPUs1ZyfNEZlQwiSdDVfXBI7PVHpJ2L3BY9a+bCMtFUFppDAkxUqsiBO3uecar1mZ9ysG
NuV+4mrFesH0i2BYj58dEmO/LB2hqyCleJh7rHgS2tNxWqWHYK2vNtkGh+IYUdjvZoiVlVukZLWL
1vS1gptQD+J45v0eUlkvqFDvHQHTx+sSrR0cJBMco/+r7i8/vY8wt9gN50MLTvPzN9N8R3jJgW7P
ZoVyhFmWrpu+VyjGCP40ixni3QhGTDEjRLRmhPwF90dE+iCRyYk0q727JK73JOj9HLzZshDcfv2Y
qV3lmPRX2e0ZWK00ldjXbIf0fGSHtw5WMn/QDVMFjm7kU8ivdDgL2UkxqOM8s18yQ3XPiHr9VFYc
5KBiXMcVfyWdldDT1aRSUadNX5GEo6mJscm5iBZTPIC0oSjBfxxWn1vTfE/2O5Ti89TGtxcCE8M6
IJ0+iUzwddAHo6KR4KvKqsNuTBtvkxcCQJbxDtO4HJ9TVSebXSUVnkgG6Frt4prpNuxBU8H99EfA
sHvA2+eflTp7FenvIER0qN4GjYd1vI8jt406a2TRBUMSguPjcHAhGBB3QskLfFLlJNQ5w9P1v7hG
diMY9GgTH9QPUiad2sRx1FO9vmilfwjgSrClS2J5vgH8+Yumv+7zn1Q1QttESgCbd3eS2FpAq6YY
TE+Ti7H0h4BuGrPoIvk8sv5NooYnqXhIxSpRE0WTHS7bRAGO1j4Ez8BGxyAIKIHK4IWP9DmFKZmG
x/OotNJwtxhgCZpxrH16ErnK8bDPytXDTGCe/kH9jVXvIKH9PGYO4RtdlIKbp4F3CW+cSjQN7VQ1
fum4LBQ8IxJix6Bycto4oaWs0WSjf24vT0v+s0M2Wrz2SqZ07nMAKh8hKQ4arXNpwGpICbvtJaP0
aWkcKqNIGxx9cKSPU3RY8kvx6gzXpIa2sWDY6G9155JBlz2+s40ui73dJ8ra4awPDxrDlDpMU4sP
9iMS+6/OVXx8nr9oFMocMCEa2q0FNSpZM/f7bCYOYtlGS0KBom2DJB3CS7+mdzYIsTGSjZmzl72F
2gz2ucWcpjXwbLxZdaON2AHDA3jdC9d6iOIYCMqKL9qU+c2DB66VTRBU6DgS0Cn21gVCJ4Snldhp
7TftSvh4yQFHBlb7lD13Bh6zyw5UGSmLFv2FluTBkgR2Z3COH+qoAjc7uJ/PWQyKBgjJDFFLC028
g8STB/B86MAMMHcFBtc8bzC+y4CWC4vMOsEy/kYx2C3Jf5dOR+OvSNhdETMLaRxVVQlRNH3DIrew
lTqUMJvWMebdJdOhubHl/+GSsB5TxIFlw3OXg1m/ZIO568z5+utBzt1DS7AXzCdLPxTUT9rbVhPM
mZHaMkpqKSLLxSNtkl2pXu39W2q4OobdDk/FGfW9uhh8V7dsMyEybtvVhSv0wC2WWLHBaz9YdO2P
fXHq8gjZVmMv+cQsrqFrtWzgALoUthcxijsG8huyczzoFX+LucsWxB6a3f8GI3Nx0Svm0MDUkEXd
bCMiEOiewKCHK6UFvQS2+E5J45vWxGzt+pz+Wx3i4pNnKdzcbEvRyfWMpkJ3i38eKy8AybAvza62
o3yYT545IirsCM/a5pfsGjii0reoNDILgm29QYUJ2+rKQ+cRhzbAd3hb2Tv0SKwtMXN8vj+6J8LP
1itiEfC2o4dBft2pSjiN6s0nyNDNo2vFhAcm5nBVMxS/fcc0ev15a7fOrmTg8HVUij9KeLd7/R2b
WRJGaurYDhPA6796LyXn94qvFGL8qcNAWD1cB0FQMPtJdHVMs56ONMO0QQ15WJV3Gcs56YDOsYl/
ui7XQ2QLjFyNLYQaQJ5VKjejUPKS+B/ECI7ofjcRfjcBtq0jIEmptTe/FWod8X8/vmQQpFJalxYp
eOpfg21kSCmtDQOxvk6lc1THxWM+9b1+HnfhPIWJ/AkKp/ecsu+eaqT+nMARE3eCLZGVXBLh7Vvy
t01FTm9S1Rb8S8zKBgY9uIXn27z0WGgp/Y7iQdd96ZAwEMv9wSGVZTZvMKGyuSQBriNpvf+L3XZS
IVC5Kyusx/46r43SXVdX3xYewgHAz1yc2MlfZPtWk007Jx0pGx5DlYUlBWT+iZ7Ef1vzBihaTBdF
mVIXM91SDT54e9bRhfu5XNGgyai1TBuMPxKtVRRUwRbqoBaSYJRaWsF/4YMR9V8OQ8Al49UB1fLh
wnhH5aunnwD9EjbDt+I1+tDD3IKQsMBg6CF3UOmy223P+U7yMWgJEX46sKcTWg+K+PBeXDBWphfx
P2gjluCZPAPR7fb44XB//fQCtKGP7lh+Y9L994DfdkwiE+LzuMRhxxf8jtalT0rv5vv7tNRHpFQ3
o6tbjM6sBAA2X8j5/HkyXdOj8ANyUnVF4lPYOirFkFw68zTjJfMp7mcgDjItpHrAzZULBVIUkEbJ
j3vU9ollFdkTQEfxlYh4S4+VvWKH8/Fq6J5z8TwzUETyySRsYflIec0QwuP9s7SMRvoZR6hDm9KT
BpNF5e+3/HNvq3Zp88DzVlkWclorSqhMFabpLZ7t3pQtfYS1FoLpcUpmBdTC0eSN/cnxv+WG7BLD
6VqecKMLndf9rVzrrXrZC5Iqkr4zKnRIIIutPdVVTpa39kh8kriNVxdbxvKPB3q9kI0S+MtS4MS9
9y3sofK9m4jnvQuuKVMkuO1i1hXk7//9QaPdxUBCXBsmHD5Dw53/rzMyEPHONXXyArVbK4ZMJakH
vgLusn9figkaHSFNX3md56wRNEfZJoBO94NL2eVRmpcrEbbB7vg9zzFCQ21h/e+Ig43YYfaW8Ze0
im0M2eBz10f03SiqVK8KHmVacoWv4qlFmgEFn/vnqcYFRH4SkDQFCxtg+JH82uw0flasDbw58BMO
e+R8DorCrbb1TYXqzF4MsN+1PqNfBJ0w5MU03F5KljJKtsiPOeHx22MMpGXbPzv/zpUVijEJoa9O
w0I/jwGMiGu1VKdw9NAWUFrvfEFiOwJSOd2IiIyjwlRyQILa4qOy7cpuDSzrrU+YNnW05Jw4LtV0
Q4BeIPi75LvQ51YsZpGS8ETAvgzbsNu0eD+FXOz8PsoypkEbh0swrL/mdgJKtU0jBxJ41vDgvMgz
WXOalqBjYp7okxXvZO7dL19V27PmSDVBErk/7KPsoxlLg20fLcCd5mV9NEMNeNTcZU1ZGJla32WS
4lI5OY4mPYvsNjCIgvV6J7ZeNul70YYzy+Bb77+BmuBghUkaDGkUEO9JACn35ce45Cb6vVI6wg+u
LQGzN8V89LKYE1lpG3oCY5bX1p/ou5g036VRiNoJg+RNDB29nx7HjQAV8mc0D8rLP9iaOdgIdZmQ
1G9f35jvmeVjTx//JM3T8cnvIzX/4NeKxLZOTnqxKWpNX3APoUIiCUMdYwyZ7uXaDA9Y1G9bveLW
xAe92Aa/HAQHvSGpnjf7LSYXr/H48yDZrf8DhezUA7xIbdsFsZor7N8Wj1cbaRNSHrv+umYQosY2
JgBrWDYHkk7dpmwJkuMDG3gOhrRV8zWjV3bfYmyijJvtYFyCQh4AJCq44W28B/hODtcRryBDu+sR
587qlVL3XwMtZu0xiillZ6yURB8Q7mPxsEGMllLd9gCnf7MOpsr6UAscwPuywVRre3b172M7yUwa
2wG4xl4O4QgXhERMkbGlNX9BuUr26R2EVJANpTHx2VLyVjYD79dJShdqEeNHVBTErieCiX2qIbSI
JAFZKQY7FWIL9nG3SGrjusZNNOMKCn7OjdCs2l6rBENfvobeQCZUU1t/8H8FZtMspo7nMEEcfN3y
FQiltucTLKTaPRErhjaYa71AFC4+J6AR/bcVCBgVLJQrztb8T6zuUxH/TClEy3me2n9r0A0av8Mv
WqVj9+/Q6S1ejyN72ojhDCIZgO5YrtzZrDxXsdGMDCGdabg3wSgN6FTp7pSOPd6XczhIjBCTB2PA
3jVelr7ocd/sKGWCL0UQ3buKwUaG7SSeVo5WrHAQXrHL7GAuDyiGn2zsJOuyRUWSdE8HSGXSe2b9
HzmO/hTppsxvt8gBPr9ka05tR4ebpJVEzbt0CQD6VMQ2QVMcoo+adGCnNR52OtFf5nWb4ahSa+ft
k6FMD0Ize3KXVsvLeivEAcr5OkZS8FsSjc9FMD2xeo1NlFLg79ULE/90ew3Tuvrz9Dl/zuq5RW5z
cETzdm9dEXJfo75Jzo3esDIUUQTUDcGup4DBc4GPqF95rZTn45PRAWHuQ4v7T9Pro2MtnHuxdnom
PXRW7iiMSY5u8fyq83NHzuTdJfBeqmP/wf6N3bAYE7UoK2Ah4s+aXeTNvCgnGgf/8Cbm8XiuDUXT
F5wy1sEqU49gfq06dpGqsChBcS4jiPW2ZbtK/VCo/EAHarJdHsHlE1rpKGhADa96xh6iiVBSXNaZ
6U6GH+RPDYQUT+4oLXL9uwj4aupvNZ4FoP2p9uwMaUyTvFbA6rbPDigv5XaV3KTHQqnOSEUjUsoR
eoCi/QLZkx6eeuen3ay8bbE4L02X05v3ZxI46WVR5cohrL7f6XicBOMP0d7jFQ+wy4qbOD0H1k2e
BKMB/ec+ZUwoU8OShiiYON3+C8Aq+WXyIPWns7shvwb69hHojkyC6GKdoaUNcrwzc4yU2nHn0A4u
42XE+ThL39ox0A3l6Jla1M+2FxelIYtn6YESRYbCfn6hwFTBnUGunM7IObHw685Rh54Fb6Vf7THu
UICckkTaulFG7hZgnXn/xfoForaK4KkPtZ53rRoYaeFIXAxQUX157mZ+W7qwJU+oG7lqQy+sjklg
wjcPT/Aze7vV47C9yZfkcMY702H2e/Yd6RCYcfOzvrA/tx7QCyBqLXuvHtbg6p3pQSPNt2bARxc7
1cF24Ho7P7L6CV7mTDFeXblIkc7wFpzN7hXcK5M8MgzcCi8h8rTeTNwuyfXcbFKwO9536Y0QEZef
HesYey1X+SPzyMAFxfGyoAhjoe6p5dPOsXUQW8Qdntatk1LU7G4AviekCvrDjt6jTIWa28Xo9gPc
CmSxr9PEE70zQSst31pEo6AcQWNbCmgcDAmj8IaosNq2pJdzFYXhfh+goPklLD83zmVLxahRZMWG
TZyRsK5kuhXmv0ZSv8njAmuSCTnaOzhVgY+RKpPSi74tQmSPacDqss/mdX+G/kQPeAWUgy1JelnS
AktK5fVCVVbyb3qMf1w2mOOs0uZKx6BFWvfDnFKefu5iovWRvJMRst83mb2Jsur8XHPAi5/JTrnq
Ya683Q6iiGASRTJ4OUI+VKWCevY64IW683/QHRey+3eXfuEUq3LmbBh5XCUH5TKDxgQcn+DfXQMj
0LWIyjyEB/N/quX/qtWprfYGNyXPWKwzhHf1Uk7BoCmIAK4RlaMZ1AS9f9sFekEnULckf0SFS/Y3
rnwNe9t3e348YJ+umr8IthhCSJKCU0dyGeczz1hJsO4kx4Pt1l0U+kTNZRm3BUfjRChZa29IYk1Y
J0rCS6N8YTiNtfw8TKftDdM5o84pbkyVQtxcaM4SBfNi7pM3IcPmkfOit0WIZNQKoXMPZHKmvka8
q+3/xMhfWGxFSXmKLsUmzPXwWdlBYlYrh4h+NvnVnlddeobupEhPC1Ad9X5sUtHbvI/rqeP7GUCv
jpxrsCdNGo82qyXgDo6+yOX4bv3MjCMbhulwSJqWA7Ko/eSvtcSGtZA9GhR87EtrExquzBVFliIL
ee3+B/GUkJeVdOFMVhPyO09rH1VuEGPKAnfEzY2vzMEackvdJk4Ln9HN+pcSa7qBFj5VltQ3yfRz
zeUXtKJYLcj8aNPquRsovRLZ6+wZXrweu9m0Nf1HNBUOiZY/jG2g+8dehlDGDwD9PgjN5vyjZ876
TZtwgTanmsCZXNhJeGR7NuNP0hY75DPgWFUL4818gD82X6rSckmQVfBQmzGsiPw2Z3h5HR+TF89j
ofDb4EUYOGD0YzKDYApUIbtfpHyWuC73QJaiddVKNGBy0TrA8F8UKQnbCDbb4DjepZJJFRqkT4XP
4pv7UNqDnki9o+VFI+KpzBjxiaxgJd4W8qQ8Bp4MW0U5SPeYrrqO3H2C60Uw/lKmdze0tKtxDkQS
9HC+syVZc7tY4yxVRowW4APT4NCdavdyrRWbelv8gq5itJjSD1mPwj+q+2ScC2T/+gOoYPHlGAOt
02uWsienEdNzexjsKo8M6v/lRDjK/JJE1sAw9Vl1R3HcBmTHqXbVOvZq/qxxg0Cbul92rqNpQilh
L7b5VRnFVkOQTW9ERrfNStv3K7yr2BiBPqq99+lqr5P9BeegRM3Ia/JpQmjyDyjgwY/Q3rEW+E08
ouXDWE8jVVCthPcCA8td6BacCy4+IPnPnloDnwTRtioqz2y3YoRUJnZWzTy7BPlrrt9SHM+hurE3
H1BoXaMfJ1WkXusLRwgx3YaiHJkf8W5pmrhlpaLfr7NlbZHFh5wi5OERcpv6L8hMasvPdUZVsKgc
Rm1fO5dmlwnoFE0Ap/PsUoUBS4j3FWGFjG/bz8/Rh5uDKwKHDzTvZ37+bfjnphoELVLK6KfIxjA/
Vv6izES6Tko7B0HKAgrTFaGkRuGUd43cb1rkvrnxZ3QMvYiKM37nRGmmCKx1+fGUOTDpLJzdDsF+
+fkx0kclWpNLelKRbJPLoAAElgrTUrd9dXvLB8jmrc4sL/eu6JRKNgCF7xWAFL8DZKKDcGGaTfbC
p9E5QfiGYMWOdpPkyin79GylnbKSxjgYgzfVwQdbJBcNDxa/NWq1Mtb0tF/ALeNK/Z/KQchkiOlD
ezdwbV7VU4bASKORbq0gKPUGY2P5pP/BepC0eOrgl5zVgO87ACX0oAMALn3i/TlWnk1RYmfoH6XP
O5eUXg4LPl269PBwpd2+/hXWKPgE8lhYPQdmTBUtEvcD25Izsh6QAf6FeSXQzJfTq4N1vToUZ7Hu
d0zdoV24VU7iO3Pf7O/QBO2sr3vVLE+5ONXkseVQuH+W6HXmYDUb0ahlLGI0gLpIIytWMaizBALS
AzgaUEYaoM5yMi66SLSOiZRwYg1WAZM/e119wTgONbe/FQsuCPMZzKgpMaONG6TfP4jCIqTU2FD5
drkbJYAlAHfkvl0BUeTgHLOikuii4tfmsFJxyDMCF82h5aHYFlM9XYZGcZobMC7TaYV/rDzwnssZ
PwK9s7orXThgc2DuWbPZBX1sqbdiNYEqJz300NUMYic9mMaQsJkh5t+UzcNiVtLCdHG3FEd54shP
/nakGAtw4lvUdiUdoaj8duD/qoe0f25O7OcbpCZkk4GtjXmdy1dyDaQ7q7OZiAVTlX1BUNTaQQsL
CTYgs7lPxGPQP2WoGvgxJKNRca7PmIshSd9ddKhIkGpWwKsnZeXmatQp2zZjZTXdXqnYKlzKrayP
AJEufIlTLfKuEfbBQoB3iyvBI05xR0O2mdinVWFHjXhoDvbU9OpwxWhWAGKWaG2GUa2wEoEr0tBd
VvrRKN7EIQnzY7m1I2WgMGxt9K7G5tASUh7F5W3wbg5eLNMf3bU5Cx+teNPwKCf7gKCTkg1MTSws
028+t40mzu38AQ7ZqOggy3CmVlM6MBKVUU0m5PVV7cemWEzsRc4JImhpvAFocgFAo4YNVs74xpQ7
LeeMdNsY0lxUHmJJykg8pMYgOHXedxvlLBIUpNyt/AdPuiB28tTnu5COr9u47p3EdS30ozxkVSkq
YoD4qu4Yo3FNBXm5Vt3kdCkOviSmreQSucFCnUZR2NerMeIwhGKonMs1Q3MDNpsnEu3MVX0UkF4p
SE2UaQ/IQNeYsFJIjQ9e5aXjCMqBxevApP6cWohJdkv3cUdC34NUw97wyhTj/sR8nT3oczLt73+3
El8PTASbzyUXXsU5PjX0VF7NMoNGIGKPuetJeSJFDHqex6vqcXlMtSfNXlG6AE+t8ojRD/uLJj9V
dEDjlBhRwrDfppDCXcCl4WsCbSmBRyprJFqObyXxCNw9+Yb/3KG0bv4Ir5W3+wpO8oQX/SEubNKq
O24sShvmF3uBi/UlKpCNmBYytsF0BACKBYKxERSCnikm9o5ssLkSYlTzNu4FvsGltf5fTTBUQn0p
hSGUaXMd2m3GXv/YGK7cBqQS65lRRoZticmHtwiuugWXfmcXp2hbiIRRCWSW4xlLx5Jk5L3U3dPy
U+v0+34bUvtAXsE1uN5BOIQjfYnzM3HjPDFFzri4yvx8UOp50LucKyowLQrj0vKtupoaYTtYhubl
v5+0Np2fZ2OhgW/p3VvIKSjPFkJ3C8Jz+DsDTQxPL3ciM8cvtnUviLj4NzMphf6cCWeLuUsytTb1
ziLpBlG3zMAXqG4mnaqbgakLGtZmmfp2Ndfs+7ooplMH0MT7qbqYFkLeqhIXHsMaTv8uawsY6Acm
b1ZhkcXexlmwu6r45t9vWIeasx6BvFVaLzB/tOA5PglnxruYvm8Sl99odkMu61rKBLpLlW4VgAgi
f2oSv9KZvPyr6qB/toezq7pYV7bgUn3SqRy2g/DvZDpeVqLwcDZqybVaw785BHggqfxStdcazaWX
ENFbHFp2gC7Dp8dzthBqK9D6t3fLCsv+YAqCpPvaLq1U2DGxegOPRp5QEkdZhWY6IZrI+qSF4HQx
9jzNqkQhTP8gaMMBb1ybSeg4FExczE3g7izxtvxmRvqRq5GywZHOGeZPKFOjeSBhDSRUiK4fbE3U
qaYPKqKZjNwWG15vsK1KIRXCiHGE4cmBZVQLfZ2HsSmWtUjE/pxAS2rk1ngFjdrUJThvItGWg5pc
NP37Hs5mHooqUn1R/kh5e1B5nd182TnBPr5+G/3z328Jy9Sbspd3t8QQoaNOLyYLfSjhTtzkQm7T
O10beGKjT90WsLyQsxMnzRz8o9dU+2kyso47LNBJ4L8LZqNwj0tMkgt6x+aE1oWNiBxxSPAccvOw
Xhb3f02XFmkO/be7MA7E95ed5IghYs0yvQquLZjYi19pQhSBbSI07H7Au3ZijGYqVlCBQ5fbGrHS
KAURBf07eO5bMXeGBhHmmbRDm/C4WjmXw1+nscrMrSufwmzG6MV65sV/9Rio3ZOiDdS1l3ua4j8X
8gGTikoEX9sEApLUskcONg+UMXpKZUTb/STam/kaa1E0BHWjNcGAq2XC6Cqgn22GMJGsKD4HpMRW
aVxrWr1vySThHCYxG5dgzk6HZqcIZtTo3zm0Lez72C1CQXENxyLcfCIosOtwzf4YV4b6jsJnOB/c
xSSQIKgy/Eh01F3mUbDyq15lgyfU4Kn1dh5KcCxSNCnkhiOUiMip4IkWg22w3pn3/UQg9WRStU1m
nZkKIewcLltTuWiNEJjOLNmwYFtEA7e1QbvM9eyJlOtB/2+PGFZgY168gXKigk/RRQ9pbDeQguEB
FUz9w8DmoRB6Dt0mHVzZgxxFAE9RZ9gweQPEmZuQMXij0qUYLL9n7dWYdFjeIhyF69nQbbIxIdxi
NhguEU+qu7CVil5GORjYgdlhCOkZ+LF9h5mL0IApB8QelzHTaVP20UV60JqlhgdQJsyNco57l6Jn
zCySHeD/dw0zfLUOY4GZKIsytIDy2AvPgv/Wy9vzb2L/9Z/b46OOJFGgNjsazT0OIu1fKlMqQ82p
JEcEkoPgX0N31S7Osjd5dHfvefex3r9iRYILPxou9/EQ8VK0AUETzwQxUY2oHpT1jY1G2SVpomwn
w83tMk0Zfy27Os08sPu0Yvrq+a3wE4fPhF8dloRwLbyLJ7SesI82DnSqfR+h2UGrIERTPoO0grWr
3pEMekgsz7RCkOSTSgmUgsdkNNuuoEuf5jqzTuEliFAg4Trw4xEOYXl8K5Y2BrR6EBMykD6aljAF
rn3I4sT6aZnc/RCR/aDBD+SGX5t6pj4g71KJH7O52BvjO+FYroW8ELZYq5fmW4/TymZ3JGVqr5My
Kdz6NxOz7FIff2BXmTgGPCEIjVsbvaurvv3Kpbe9OMlXog6jiYVJV2lYT3FikQNQYfZoC5jJJVst
GbOW3b2gEpYjOjqnwpbAla5PQ3oeV3MeY4E1MqqplNF6rnBiRyeKHrUsWGCw/P67wfTtpIqY82TS
P0Qgjjmybmkxn8IA+CXc8oz1LEf545aSOqVzx6XrU81oRwQyhAaurvIvPhN5SuecbrilhSKtCe02
CNb1L/6BAsN5ovsIX937B+i/MfoPb4Y3CxiCM1y34tO1jml7QMseVN/cK1HCk5PeQIwc1aYaGNlD
MBxZwqQnotryLmFEczZLqRZPMwbaDs5sCAXfLMqR/GYL+squ3g5g/sEGuOJSCe5wzkl9T3FYYxZ9
/bzpucmjw69q/kzMIKPHkvvNk6pAYAczegDNSRukIjsYRxpz92i6rW4BLyf64LprjfTVBbcF0vPv
0c70SAcXe+CV7hnKV7ExPgKGbhcj1Y8/qfh35LmgidqET6lqFqgoY6mqykP7RBI3AO4NZdroACBS
8SiUG9EInL00vw8PaKbM38cvPmkPDFYVP87cZB7+soSmribJEpwMwRKuu8/EuNpKaX+EjGMAZrZl
pYcLRUME0e7zi43uvFD6Vzv+wsMTTKFRMwquyQvsaB8vhUm5QYFHsk7iq/a4bH5W7x6u/4p4Qu5y
ZL6+s3QKcbQ915P29Ts/XUVlW+/ncnAD20xMeO9XB525ZnX4xKRGnHKQHrB588BS1EN3sTu4Nsnj
glJsKT8rkF40suK1Hdv9E/ooHnVtVIBc8kdB1ovRCiM5Ryh7AXV95k3+75erFXgWNF2EVoGlz0zR
cWsfatGzX8kR/Z7vjotDE/O5wfrKrAfS7mkkM1DixpdNV4IEEDbP5FD9it0imTjGnd5aCstb8D//
Hdh8+nTT4Wm59/DI/yYiXxdVcoSwf9eVZ6O9zKxZ1GCBo7qOIXoOEWlBIE5qxFyI2y3MsDHcbNmr
1+4HimcediwZk53Ye8i37o6EHdcmpgQ5VX4cV2CX8Oee/WDRQG+DBeQM3iITdZr/I1mARIf96pGE
bHBeJnqarkmOiSXPTlPCRUlWXjWD1LQKUBJ6FL9or4uDpqEus12TPruvkH5Din4C8yIuSo3AyKGs
OrdXbf14G9YTesb9VQRb1Ftx8Zoq7kV8xlrj35ybgymbxvYdTcgR5jsSTPyYrTcsBrLGKfxCdQoK
tOp+GEprvwQ33wfBvSvli+P/VDhEq/Hdaj2D1W9eWWg5kF8xTOqmlaDCYCOXFyY971nFGUpRXjCe
NhlzgiWRSWzi79g2LXcK7qIaQn+yurSJRoz4atZVBb+tEyyFlqOyPAXYpM1SRAh/ijQnccewoIMq
XbBtMdYirY9T6C0sUd/EJgIallvs9RE4y/kPOdB+wSikqNedcfAUccCkTt3H8j73Y0FXwSNj9GVe
2O9wXdJ4xSEmv11XzdrdCcLyUKHyI1WiuZdXq2+dbV8hsxF8x9N3F1VjANMlS/XZdyPHI8WL9Ul9
sdh5bKe2AiY1NblSxXFe8tVIwyh/f2Cy7dOXTwyHA6+sHNNV3+KcIfXnXVIPfdLenwEMFKtLh+E2
dLCrwAe40ZrLLp325aFxp4xy4fS/UNm7HgeSixNqaKTH64jf+0LQ5lsftro4KiVCSF435WYfyiSa
684G7ArbgsBcvz59CIJuYAFc+Kfs7aCELXuysgLkauLg08zqP3ggmGvpI9vbVpmbtve0jO4nC9FT
30L80nEqc5CeSZJUS8FBk9BwPjuujayCig5ruAePjw0ay9FrWYJAnTXqP1hs0yRQSJRCHjPGcBzR
c0qKvz/sxkDl01CULyOwo2rnzljCy0J2BF1DNjOxd2eNh6KJu/JiNHwintYYgymI4Vtlath698GZ
nOWXaVC7JfSzySgKpFC7EJz7IG+jk8Bs92t6jZOXw8dafA5+phMzd4O0kWeW0HySj5M9uEmERaSn
MlvceC+JCJ3RoOtOHsBclGKppIyJ9GVAV0n6BGmi4ArGKt6njowiEABGNBL+kuRZGaCblC5vQcPA
OyA8r4sNZih7v2WVhbj0m9ziYEl/vIodoEqB6PZiKHk2LRumhoVoFE7zIbSTNNc2ZtTuRkbUy7Qw
Rk167ZqZY5jVRmlVAgUQUXX+igpw/T5Y+sp3wSywOl2U0VqySIvxteAVMkL0SxWdcyH2jfsaNlXR
dwnRuQS8tzcwb33mIF6TlC+lfUifM7gl+RLsrJPgO/laMBkV4aJ/ailuSZ/iyq2F9qbE/XS23unw
bDFtHnF/rEAD7UF6VdYiF1LQVc+KHnzE8yRQuolwUpTijanQqgYntoUqCQ17dS2S1kz7B3D+Z1tD
umeB8DZEqRjr2vRQm7TZgkFpyEbeT2DoHtWM27LSEh7qQUBKoaEd2x9j88ZwoISWbEz0vW0cDvXu
ObLtNvP9FYyFpDp7Evyll6TrJPIpDWm4p9IQhZU+apsFUoTt3pUkmfuImAjuM7P8WuKDSZmLrJMS
LYcpCcevJfUQClgA6JyisrlbFRPxmGlPeqCfrrio731oH/XQgzjXjnStTuIelYRnLKa3pd7fDE4q
792bL8siHexiir4/HrYpKgxRNA/xOgUbEesmUfNNtXVIPp7lwDIU1BM5SukqExJqrBkLomFx11Ln
WCDpYX/S3NkFi79kCrbIA9A9hiYdO0VPrTFmLC0nxmAJwz4vogBmErWpQlTQG9OJ42YOfe7/5mGr
mo7/bkwQqnYr47ZfswrGZY2I9mqKBLGDgWZAljRBzKyMnKCAOjQaEyx1+jKWBKCP3PIP0Mvyo1H1
CU/AkiTb4fuhFbeip18H+Hr/VNQ5GDebRKR1rueWkjEclZOT6/874WYQat2LMw9VRgJNyZR/9Cmt
woLZJ/lWaTFN1ypEz3+dGnjE6Q+zkb1+M/7iWSpwVQWmsFbw6HhrvRGmQTbCTV5uFvHJUT8g5XqV
hCKWeK/dfr72wIhXC6dtL4mDaPTX0L4i9X7zF8Ku68qQaaWJ8Lks2L9wX33b4GBbn8Jmet76mujM
wTW1EcDInd8Ndnnf0sLt6+RuStObPJhLhXS2Cgbu5qIJaQ7JfdpopFyrVirV8QPL2jxnIPH3luMt
HLm9tCggsaaPeKdiooRFU9iaDaV+grFe0joRkIIRFmnLnQJtmrIPOATHm3McloyKR2jJRDkSpQL8
AX+Oz0YlEc3UHxh0aevSpAY/QKSFGNp+btmxc7GKQK4whAQi1bGtTh4xhlCQcSeqeAxk/sKtxjgE
+c+IOcCsDYx9bxEviSjlHz0DDf6ik0LnR4RGwmjnofn+u5IkdL34XK6LqSJGMiL9myawMBks8BmJ
HKEWmPKUlNO34iBK03Ag1RClvuR2SxnjT6n7gh7aw0f61QCg2dMI+SSKpzSszEJJonCjm/J3UiFe
Io/muB+9HKwQy96LyvC4uJvszCUNaxtudb+wsuOjRQ2CBnFlgTCnNKTVZeVCiQzUHVA776rXDT4a
rxhCiRgYIanGAC8yw7u9iRAe971AQyQtF4EkEQWbIwStmm5oAuaCxt5gne6OwzavCoXxiPpKClnK
izMr/dIqd4p5WIWAzrQ3FGRaM98uUksPdnlroIhj1Y4zY6MEBRHpFOR/hXKV2l4VFuIZeOOLr+Mu
CEUcuxEnY5/dxF/mmBJP4ReFrnw+umg5o6qeD8Xyq1YWH/05/1fIID5mC28jnbzfTxG5WxbaFDcQ
7pwAQRJQFRNR2UJQKUBB3EUUzrnKtAKZm3pn9YV08Yq/PL1+0qk+Wb1ER53Y8PHBrn/U1NqhVP/Z
RstcV+CksV3UUfnYLkkvRoGeQ3B0rLfeC7nZ0YrMJD8VlFFjzO8D2pZL8iLyT1HxGDv/ch0wswZ5
96r4FFF0sHNd0Wk0BKvXpy8N9cTVo1P8e7jwsXZGVYUfn1/ZJ3aBOFJIEOXglBfWN2ETHmYLnc+z
H+m7jcKvJtW7f9P0WhFsnQlZ52gqc94kqDbh6slCnvS6STzfkIhPHjPrmtA1WoCpRtZSuYs8wt00
mzhYiRTcchBQooCD1GK8rybHPoBQRCjmQp6j65pdRZwwhndMc61CuA2ch/o0Ep73zQzJVctiEnj+
BRHInA0vTrGW4Xk4pSNmXNNm0P5/oEcltbXnGGWgD7d9KFeZNgkhN7wDrrXtpHa49Cm3+kw+Ig5f
YDc2EHFy/06jUibP5czPCZNJ9SqEad+SsTfXJ3zPCN0Uz0se/v/zocxO+v9W0vgiY2lkGuFBqXXu
Ip70uQBENt8OsXLzxZA8Y2hhbB8TB5rgvnmL6XiVjvBv2JvoAJ9Yv+u/xrVj111gx88TE0+OKRFI
9dAHG3B5SwvmxuKJ9sUDEKTqIILeCYrxZeWcblPeEvHVxTQcrKdJMoBkIKwO2inoiT50IBT6x0i9
XM53VEFWbZ3tQRJMz8NY+r3rJnTibz9ybbhcaX/hL8jo9d0/v2Qvb253FHriKbvYaeD0IA2QL0P5
iRN3o89DBopwkEiTyxUBzC7rAi+YnDxw94fTp/EhApC9rYy4lFY2nxOm5Pj+R6YTpPfsTSi8D+sC
2u1EQoZj3QOJvgJS9zEwbh7HeSMYdEF93zSeu1Ub2dHkLV9AkVstlD90Hxg1jLeWR2nCLX0ErB8t
XFm4mwbHUSNLx3/fS+YNr+b5tqTJJg1USrfL2DVArhTSig+pTv1nKMecjpFpocZV1NQsV1blkrDc
/HEhaJ/GHHZlVs48O+wihGch96Ad8xkVDlArSxB3YJpq6EoM3AlDz/xLu6tBocgzRyF3dZUIxL2x
b3pwxcX02IRMNPwtTPqeqtlkTGfjfFYD4/SJCtunQynqUmMy42oA5YEnYZOgzS63D4tMrd5UQ6Vt
MxWHPvbW6O+iH2vx72NJpbV13s/uTdjzfBw8PuS3NZsXph93GlDuPpNvdqxeSgr2G9OHdliV+MyL
UtC7YAv5yBOagLtT2vlhHm1xseyBlT9A5t/Rzq8ClWMS3JMAgiofwsr8L6qlxw7ecYXmFk5llpwS
2pS/K/8Mu+ASTHuOiebsohOc52QEfmhQfCl+3y2ILQsNcK6VSnB3oj6o/v4gBOPngaHzAaIHW/Db
Lz4TKZadLuWCO7qAx0zEH9TV037K+/DP+0g1U7Y202kdQg11s8x3WqIhz9jIumDJ1WhjW49m3aST
Y5A7ShaAPkshyVl22jtchlchOC3uIyOee7oDXHC5ET0IcAkRm2mDk6ozuep4HIXgn7jI/3Li0cF0
iyHR0IlIlyWnvdukylgsS0TdUuLXeKQUQBA37IWvjywq2FUeuxUUhrc084Bxday23ZqE539qVkSv
6WM6ZdzA+yCTkv1Ig2rH1NRNXy1E1HvGJTgAoAt8G1LnszxkmH4/SvbuTtNs6a6PCbVIElChlzWC
w7yLVtA0nNRnSyN1/6kmZRmz6HCYH2Ljo+lc7DfY0oTZFyeJYcyoDPGKfo3BrgUh+RyJq4USRa3o
AY7D/z5qAuF00q/FT4oygrqS6sNm8RXD0/hy07FmD2IXUp47Ldl7fakQT/mlAcslTlNXcPK84Z+t
f2GmXzjEwJB6GOf1VP+YrtK21F5sY2AaPJMGraOECIEdo2tixYH2bxywUubVn0xSL3gPPc5xt9BU
4HUnAjeu0UPa1lV49MJDbdwVKHQMLN60qvOWv/KhqYm3r90iNFWLb78y0sckUtV5NGT82KQNDtJy
2WF3dEAG/OJ3vFMDXUVk1Gw2WCDEW1A1r2nBoG9NdY29/7Z6vdPbELNOVU5dPOevaPDL7VEvRHCx
Ok+BpYe6xFW04EMnuC+IB+Wwx3ig19urOpiSVgjrhrEqiTkd8j1UWDnTZ/H2ki5mt8ynBVEaCFph
HTK1xpvQKmzan2/olUwB0oKNdztt/9wpgd9DB/wzmtG6x6F2lyDHmw4u+guuX5XXuskx4rEFMACm
QgtkoghXVYGpfYN440wuVzMXWkdJ6i4RWNeXDHxgRd+YF7+cpxPgmlAv9q4IR40e83YTRvUPyWIX
9LtIAlOGI1kOKEkMlY663rUEphbQp1eEmTlFIzW1j9+pQ5F/4xtbY6xVvT+eMO2zRYHZOkq4wqf6
Ytr4ANl1LNwB18IB/rQwOTQKEkR1vfur9tZJFNMXHf9FJwIVf30HpaIyXqeVvV7HIbBAEan8PBUs
iiDqZaS0iSGRQyZHLr78YtVE/+xcTokPWWrNl76MYtxgOYAmcVVF2Qsfsv/jZwGPrvE/hBL16ega
NwboT4RSoMEt1eKi/97ocAffQxoUq5HPXCXqLzQd61P2Os/uaekWK8ZpzTY/h3cL9vvpGmatAsNA
DnkljPCoXnj6+FhuvhOOflsU/gS8bJb4EIIEAtyNjZMLlzzE2oDE2CdkVkjtzd/STrZiU6MvSKHo
B5Lor4aeJNMYmc42ewCEPk4ad3xlb7kAaorvqyXUdi9uw7iNitdTh5pyJkfO4W5IWq6N/mWNjf/D
wYK1r/NUUF5ZemkWZpvDQPhL/jyMJHNenNoR+iRvsNoX5e6UAStgsVDwIm/fnvPq7uDV3/Wykqp6
nQa5thoTHh+7C7dxPGW4TLkxdZ0B2K9T5E62sCgF9t1fZNOWVAgFm0x/Z367NSS6lPFPWGW0DMpb
KIyVrE7QsM1DlyEiK9avNvawclNxohD/R6gcQYn56JG0sSFWm5BoXBAj0jvD+XdqC2bTwOkdz8GF
NKizYceotSrg1xHU/hYnx/N8/o4OARvzj/AXgALWqf6ERnmi8/iQCay8DO8RGA9H98kcWmPA2Edq
Ip8f+2lhul69eXuF6OKerc6P+qkgKOFMVumM9wjuh7zd7pLt8K+QpF+oCEeErbCCkTEPsq2PoWdm
bkKBzyUuNHSHGsbiW10ljJZyPfLZauRPs56vUB0ki510lB4KpEntrlgUZBs662BKAw5K1oONCXkO
BVt7e9mw1WVMezFUVvVvbheNkAWMYY0Rn2JBssZJwoD9xVxCBhMR8wMaj4tMfgEzkw90/MmZOqpR
AWx5bJf5ID/mBTE8F1gU+SuSRv0pe08ffGWLGw31j7/No0RFS1Yn5PhfT6FclwTNXxgT+ro7CE3i
FWiiJhUrCIdRwusf7VYLACXXkVy2AgOIoQePuS2Kvr+sigL/upl6rrZoODTxopp3mpvkak7NXTab
PH1A738o5Wj/rpPtFOp3URxmXST1QB5hk0L2bR8tw5XzKh0S75fAxhGrWDs0wEuHnLdBaxvX1C6u
Kb6SU00acM5dS8kbqpUGZpvx7yZ8g+keiqcSLQmkcBvlGTKtX1PGwvc9pzm6FtF0HG9qR9zwDfDv
T3h5BLHEXV7BS6NXtMrnZmctLxhBIHxukyn1UkR0RP0bF7Z7FSVsF3NEDMtwf923OSuj03I0GzdX
F1ucqe3fDEdJ3ss0r9lIt6+zNQrC3AWESmSFDL04m2S82PXt7Llk3mlNl16sVa9XUWZYgCFbgRkt
3G3AfW3YHE+JrecpzFyLvXWvWEZ0KW8NRZf9OErTroqCew9v0RZF0JXSKXAc92n3FFspxXAk204f
kcLM9aqaXUkhefIVtEucnEkAzbAPF0/Cvwld3YwMPVIEtCo18tnD+w9tHNsvEDEkLjZ1viDORKVe
SR625gITnH3SGLOFQowyyDkyByPhvLwNmAXPpooPu5jbWxYx/L/6dLcJU6B5ZBDvI4HKSE+p/UUl
VAHGGvEU4HQI/OPpR6ewVYrUJKvSwBVG+Se2fn8BO6sPY/nT6iLgonAoUt2zeu9JCJ9zO1JcrfTk
4H/1PyzN+4TC1nZaqeOlA7GPC6mEE0WZkbH1lmuyoibpRVNrlZLeImK/6DGKdOTD5lXu3I9aTjSt
GFnEiUgUpe56juq3PcmW9G4x7CYcOoAZqwLwMc5ft7m1xtxNw8G/FXLKKYWtka5yt3kI6WzdqZnc
a1K8p0j+No85uzBjiQucm0FgFSBl42kRh/95upggezJK/sr50yLNTDk5YTzloWs5iRMruZPzg5lV
BuYwsDx505jQG4ZtpvKYwSW/wUpRkRK79d5Fz+XFbz7r46XjQ7XuUMpzFQOEUrtvouSZccI+DnXe
obtazPx1kXwmP5fJf2PqKDhFkPZmXrSNJH26t2pWDO8dZQH5Ut34I8WjmfRV8tfw0uMiL7ceUN1m
2f8nynu2qF/O+Bee/3xmolyVU496LOI/L36qFmJzTq39GZ77j+VUdnjUyDBxododIQqV151+Ifwj
jVngrqm0ihtgjWlEXwT/c+c2PXc2M9rqR8TMSKGQDQtwFX1S6vquxAWDLPkvAFQzzrfeu8bFIv3X
Sdmo/7T6FTawiDSS9ZvTxPl09U/7zmSa8jE8oUo/ruX+Tsk7lfzE4tHXCWQtCVxkMFiltYQMHeRd
RJw+LrEBBO+HiKFxr1a8tCfGxiQ98TcmJUCFkT9HAhEN40x+ka8nUC3YjDd1eAnRKo1XM5sHbR6G
re++OkTXy48w8AvnvqM/pdItjSEDnrLCriAQbOm1Yhvmdld66NUDbGD5zJAbZGhKS9MsFeXIRSJc
tiWy/DyWM0gfU07tFuGLNAOVn9pRBlc8cfBV1OwRsud7cqYyhQ9pcBeGIOKV9LPW1fPNYD43b9TJ
qwnIXcobO44vZX/IhcaC4fia7DmnYgriaFzVFG09ca6OxTdxVsABVExgkpKWbzc2qdHl8edooJOh
gjNVEVjcCVnzy5xdwWLvq42zJpQg8bGkfS47AxW/16JjfuXZ4Awkg+OtWXMB93ACDK6ExNrxPJ9u
S4ZF17yx46FXRUEGU5QV6QNYewP4Di/2kc/YFOH+SNUsIDwmkxIfBOWrfsaf/JFkNn5+SuW1KyWD
aHlRkKZSQxVdyjWxuKPP6WhMKYOEL5U9B6qdjyaJ2nRt57muWRfoOgPGoncIuCHuRuqJjaMZ/JKx
JSImyUItLD87oFgO7yWDqs1UVtugd/HRnp5Z7NhHTHEv5ygTkebLQxROqdkwa7YlrfAx/fmVoCYP
3b1zf+sygJUpBgc/mPpmX0M3AxKOPhZN8B0dPdpsVSFu7vgAYcjl6nuVwpoVrihjjL3ZrjgSmtGX
wy7Lxnv/olYa44IxqJiqljL/LvPihfMCLaHPnvH3+1N81ddHfRwiFsi1vF+Q3IjCkd9x825ENGX3
WFeGQ+WXCB7405bj6rbbxjzxxAY1Ap5lt5OGbtzHxrSoS9R9fQiqwHSoN5mDyxVaXw9nB27lJZzC
Kn/uKGt3b/AXtIgIgWp6cNNwz4O/y9yIu5kmADHVZnkp2YXIAERyhDN1qh2ra2j0JuyL0xa5w9Kd
BvvNKqDs9XMc4PXPmCjyDiLChoVSsGFfsfqIihk+NgwIYVM6iiE7PVQtMHc+NCtrDO+Y2E1Cyg4w
turZcKEs1gcHY3PtWddi471tspLJ8M81REFN8GpThifn36olHmiGtyEmsEAHiO2A5vlfP/EJlnv7
B1dzgZ7f8UQHTdaIzXNn4JahXkkN03H3A4aKpbLsHYJ81I4qVNBtlbxbcgqA38OZM46a6KxV3A8A
4NjV3k4RMzHyum3MNl8NO1tQ8PyY13Iy1ohRbIrXTwfXRNpo6iMO4S1CRxKqniUupEEgdLfs+VAi
EZke753ymPPmdWdSG78HCId343mH/81C8WYn9lNOrnUKnoij8laVxBA3YfHcHDycUvbAx/cfz48A
oRB7hP16T88H39mLj3kYaKVWBAJp9TNcRYcnAX11BoFI+Otd6aiLU2qfSgFVaf/62khFLBIe4ngc
47W/Y0KjMtw59C2FWkt2Row/ziiQ9V4y6IVuuKwokqOXCmLVI24obw2F/yhN5sfJB/vOyEmEvBCD
iS6OzAcgxBJv6X8YYdL63V/M1ErnxJtj3LvwdnLnBv0ltwh3FevaJhgY5MEiAiCiEVzmrapiCc62
CGsVEFeYtInWMlL1Q8Tn/FqieA6i3ULkAAwUvUcTyb0hdahLtdOKjJ59K8SlPvO7ojjLwd0UzABg
aQG3Yw9ngw+/b0iwk/Xo64UhgHSva/S2grs942pZE+ubNq3C+p8A9Uqgv7QSkNj8D+d4J9Ru1MIv
qnm39MHVH7qeLMXQsS8ruE/rmd8RZj345xy3ZApb0zwGdiOu8sV22zPzUc1HtHwwqvIQtyoTC80F
2oLHOOIwtL9iuMMovhi013P5uIoqc+hsLnLdeyojhuNH9ziyASLm9Di0zAlz+aYvW3+YPa/HkrSm
U7yandUKuexfhRYnfBsHXOH4kFJ/fQlsti0wY6I2zkZPAKgFN4AeTOm11WMBrUKz5ynIG3e6Wo+J
AV6IakBxcKbC2cfdmphSzXkxZeQGW55nfseYoInZa94pQli9wmjjTg39DpFZxWG9GeEe+S9KIC2c
Sey5GPqvYZ5WhaGkiku+EXkdS8ypv1cX0nlI5JT9U0vdvXJQcdBntfY8JJlRAN+Y/JnRaGlCEwJ8
vTreG4ZHbAi3+UBSTnkE+Ta8yGnRRth2YApSSQpF3Cf+vOg7R8Hl0LZbNB33tgCEUuK5JuvahmG4
qu3FrYLylWEc0b/KBfTG7MMXYQopaZKjtGOW09eqikcNr7v4/BenV9tjvmSujZh+NBVcS7tIqP8s
pJwcBP32OBkMFRUqVDALnJb8ogoD83A/WcVq/rSyA/FLUDM/LfX1R8OynX0y1UJ3jtQptZ/kBYNH
uuy87zYjk1/8OquqErqkww6THG0EYMxVyHBDJbUXFi4OKwof1jnSikolYK2fE4EFa2HYbC6IWj9K
S/mcAoKVTM51b20+EGK4N7priB84PIdWnC74JuD8cRmLKph1EeHBq7gagKXcN8azIxpB8+yka+kO
5nV7Ul/AYwUwFKc+JnHf8e7EyV+LclGN3Xe1BsTeso4r8Nr0MeKZII7bN1xOMioB5Knl+hdAqC1j
d3PvZF8HEB9+EZ7AfnSTiZXFRYEQY247BsMvCbpLxpkp/oA58LpGxmgWhEB9LH0NuUX8rlPmWPJ1
owwg6INiKCns8LsD7qko3FvO32NDXs6YVmDjxctQul10pNXJD2KSSnPU+GiUNU7BgByU3qnuB6Me
lp0sF7NLm/YlmEF15DrAOJ+j9FMJilWnGaP10KcjWgBXW5ZwUacAVY73cJAknQPfdwl0nAyb1cWH
mAjcalGNS3fYvfW25B9/JKQyYsPX6RUC7NN2Lbq6HIBjmiocMAYKKZyQOOxFMB4KLZiowfLhxPRl
nQz/N2hsmx53TUNNa3Q8kG+VGOgwDdd65+nt0T6vrFqCNonRFI79Z49vqhLXFdntTsqWjqzc60IU
zU1Ney09Rc8tOTUEK9axtwtcc/7yT+EUrVLorZIcvTCrqQI5CmhI9k5ROxLseSLaeMB8iZ+dAMLr
eEfZC3ct4dfwShitEUgj3MYLoZC3dcpOCTvaaZECtRdByz81DqFCxXsbySBhn+/EMIsM6gAHojOe
64AfJqr5rNHEF2rcKBTMk1+qSZHJIXDCmCLGKOB/uLA09uX6zFB3LZrM0lVH4K8r2avl9P9nlzxb
Nzlw983Y2P8bTxmV/kD8tW6h9PqafvDxNvZAEPnlpR0LgRMhUjwbiK1/W63QOBWYVGxlcMTmyt6n
fDHh/Gp7dxaC3e0k9s8X6XfYr9/JY+Ersj4CYgfvz4zp0N5+f5gm7pNTtjZPUq6LT/zss28jofZt
0u29qrMx6Us0gl6tnL1/7YfqT0+kIFZrHoHLKWaLoEvll52mt+Yw0Lu6U9Lm9xPBvwlJ8Ay+ET4z
9bn1ouU+vLYC/+M7ChXs77/Q4bj2E6iV6v08VmPWTVBYUAAEM4SR4Av2Hqvu0DCIKwF90930da43
rWzgnXJDLC9v1EnUjq5AW2+9JP2+5dZAaTYBA9WW0zle67Rgj4I6va1Y6pViKb6QHNtlcutLzfUK
FNMuYoulrH4RS1iIkpKCwHFlehGGieRZzVF8O7Aa2l9WomEgX5ZyiTZuEwGacX0qnngPVoD7xyKf
IAxEK82Nb7d7Py0VLdi+uaEPlgesHT+T0Mc9mXPzZXYUkwpEMCr01z2E618UmgNGdesKU3Pp9ypg
muK2CsQ9AKOl3afZVCW2lBFQPBgnfQkNloT4PL0JJZXmeeBA0+lkRX6rtI2mdIgSc1TcKQYJrajq
05R5UMZzpHjvABDk8JUt/AoNDkvOOTmWTuAPR7FDrMflWSDz2Eh6nFSNBwKo5GtBBhSOBRURknb2
4LyBbM0WGP98llrIlN0K+ngoFC4EBFRnKIebq+ToYNWqnBlsxdRBx2086RbUiU8Oh1a8J1msi3FY
iohjghm+W35hQBlBG3ZtymTGcPl7mBIucU5rhvi1/1jjX4u24lau9IOxft7MhuwXr2aD1JjSDudB
d2oHLXPCPGSf498dai8aA9W6xieipedJczGOD5MZ+sd9Os+BKaJCFxsxtFY58xhw2FdDEicdUiP7
3ooBSH0qpcZvrK26M001VBEc4xq1V2BFMOdJMFmE9icp5Ssd043SRTI+xXDgAAJsk8Xi0RiIdpDK
4cLP9cd2n3Z+EoFt/yQ19PPb4VWjAD7bEKy4g4+MT8YCqzv/yR4LB9YqmNeYWYWlI0BJ7nYjiV9B
IQvnHXk4rzKHQNbodFNuanYPyeN6gzcb8HEQWMXgV96J8Dra2lEQU6RfxOGEtKrcbyVoYfV+0Yft
m52MTGOxVP/IvN3tAEMgAQFr2x+UrzOGL6uzbSyAwfTLY+61rm+zGYOs5gwY/bg+NV4MDOVObeeA
dwTelf70q+XY8D8ZR6j2te28qK9j2IV4r0fjB8txWJTXjtI9liI1Gst5mjj1mJ5oCW3hCSsPPx7w
z0CvaTrzFtx/DiPJmPkEQrraOm+UzChAKp7Js8PwVK6B1at3rNMLC/UKnoLHqZiY5+NglbSFiohl
e3/CUezd+CB+h78ZosPKgj4ZJ3hO9fNqqxuEuCPu3MDvEWIP53wF6iENmcXTSBMdDa7T+a9rCAfM
9drqz1fRnNc/TBeqNWtHwVTqVlL5DAmf3prOBVazvYihXJ8lF2BTb/1kowq7WM0QxlyyQAML8seH
k33G/Qz1enLFkoYOBfEVGgUFfpUi0bJ3N+yuNFgy0t4/c6EkogIF0TYOcbKbq4fhPgYNZxmdOiOi
s7FJeLt0vYLTxcW9hCTqUBFsLJPr3jxXmgmAOdBuiRLs30kpTi9vO0xP8nFTBay6bqBmPwYyDLIf
mCRegfsImhA+eK8M4b63mq7L62r0BSv0WX9/AmSbTIJ2SrvoNp7BzvmS70QulkQLHPoojR9hqVH6
O22XrP7GNWeFZ3V4HEI9E3NJZfc7gn0nPolHrR6fnsU1P0gBVCteCawRlmAZypPCJOJccRl/goT9
czuXeU/XsUKG2kv7s3zH2vSJuqPAIu8iEvrlRf4N4Dl92l7cWEsUFt7fJX/MRb+McqmfizmdAEh2
9trjjmHJLXUrRGD59Eb3qwQ4ydpVJn/5cOsDCOjz+jGWoyHnBHh13/J54WTrveW24rycXW9lTm26
ZLCa59nV7cYQx++GkV5Q34gcQWwV7gCCAib5dvgUDFZ2rjvYjMlrFeY662MMjvlxBUrerkOU+4S+
D/OWP17O9YCfrGOvnrF6RHE2gNHWmPLxUJCQbVE2Uju2SSVrTatndoWI+UzHu9ITjta4VExBVEQx
wLiZGtG5vFNZ1AENQFGxMRSafFGSR7rXR8M24pQLMHFRWGSLhfPV1S01mDLlCbNokMjJRQlrEBOV
54TRJETJIoGWlBTmZY2P91Bavw633IMs0qm/5hjClh3pde3uefzrtHr2BhYbXZKBD3AZfVQA1M00
S79zM2GVRokUBIQMXX+FCNkafJiVgqdf9plapXVMmWwPW8mR3Fc0ZHu/gjlWCQ/GusliRZrwNPJW
lIWYbJE0TRqPm3Bo5pBGd9NWg8eoxcjI5c3SeBwrY6C+f0Zvw9XeNe9BboLJP9C2imvzOlK1aWA0
H76b2nPknvgw0L1RFmCZftgYBjREaKyB3kM1N1jWod8WVtwaPlg0qk6v1Bijv29zaTVOFn5FrRWX
1yLn4jR7Oqut7OcgzZKBYixSsEWZxFDx8njxieXAtnDrzpUytSxKVtODhGKRZtKT7iT1eDCeaSnZ
qFOGvqwmASLUjb2FZIDxAeGblfQ/V+lvPbvfSOxzVpZmet0IYgRuVMJYSKS8Wa/DFbVdxWBRH8b9
AHnh6T67toU+oki3Bmwcjv0lt3pPys06jdvxz/+r0GTQR/+RtqQCcaa2FWZr/feQbPnNgA38tZE9
TVt/H3VmpbAixlTtUeyIMjgpcqGxy3WOT9nxPlXJL4KCDx5b8qWsQ19Q5ZUCdmfNCAHtuZSrfJAL
YNuiV4qnwod0v+QmDt2JwVcC0KlfExkolSBIySf5rXo61lD4Cliil3dKYcoy91saZF6dwH74lUQ1
6+SiIOhZZieYbcv4PHPWXUvkjRNk/mbmls+tRRjbCcImrqdPNdkxb128P4dND/hZmWqNSVUa1DKB
x9W9ysY9+a+Ben27DUCvprEQdd69aUYcb5n5U5iovq+9a5SRtj2+GZWxm++CqxBfEL2wYMwReamq
A9LlZeX0Oss2kl6UGl2/o33h5YBDmUrQR+pjWIoDSMHEKL6nkGRpttPrAzvoDKEARw5hQZaco4UK
hDN9Bcrh63jZKK4lQ/AHRmIgkex4WTK//XOTK2kJrEaDnGg+/ggITlW+aQnJIchYLVReFOY1pCVt
La6ewWQ/Qx6pOBqTIA4ikLvm4GvOJg+Ct91hVshzAkurpIRMnNGedpTRyey6LZSlh/7zEdhzFez6
qTxGhXSFFJ4wJFeZYLelqGF138lmj1SnIguBl4FTy+LWSQFwsmPp5A7RU9nl+m7MbrmNKBQ2Oz8H
vySbsExtmSCuAWkS3xcWbT8Utg0y5pVxVRFHMREek5Cb6IvUuTPK44jwlHjmToJO4RmcNoIbDxC5
CW1JShwLKWmzTw3Ha2mFTseqDcDGvHAZlR7y6v6VU65kN3gycsCmyNu2xI5FYxnyiGZmErbOfAN4
/RGoMi5hrHZAVuJA4AIlpJyqVoeGlI+THSB1I0Oz8o0mf/4an2hoDlQogc4x+wGITUo4uaW3xuN/
eOe27Vo/kOkwqotIXQ85Zf7KEckX+mwzeenCGLKBdg8QjkwIXtmuX5K9FlCOXIXq7BzCQRt9rs2t
Ew5z4VYDO7q3YC1LjR7800khijotI5TD7xzY2sUxB4RNrQOWQBFx7tw4bpS7PwNCtpNYgI3hofPw
HVHtrfFALl3rfZ2pL5ZOGBMLWTINw67IyOO5HgeccYGsRe/1lR8bKuA/VfUI/8hYPqbGBHbVr40H
ILW4ZAQswgjM9+DEJtZpJWsTdKSC152fSQPqiTzEOMifbhzkAMmK3Uuu+9QXrp62DDOh9QSFViuk
CZppI5vDP/NmeHSiRd6LZbJJHhZIz+KyDBTqz3Ejodpz30sYh8EltMxNTAr8UJzeMscWhg5DJWCi
AP22s4k9ELEUmOWjPg3btFQLINJ5gFHyy+ifeYiYvP7MHz1Cxz4epqMMhcDiG71cet8VBkGv88oP
gc5FvGlu8MsewKBP4aVEN84BgjcFPxXcEoH9bdz8c3YUKZta6eGQY0uQdYC+ruQV4AlSL9z2pbt1
21aZfo5NMHE4Oq8KjBM8Ta5vZdVnArd96wB4dRNG1Z1rmWUS5Y88JBZ5Enrpqm5SmhtSgX6mEfGu
xFxyeBVn3rSOdykPaiWzipyHSezoy0fGNXIa4vqeOBYscK2eIl7IORfRCPpw2YwaUh0v+16rjOQ6
yLSKm4IXZN3qNQpOjyoTY8upKELJpPIRSyQB0d7ZyH5PvTX4GMxv9FO2r4Qcip6vr0x83htJ89vk
J6l/5KM+Sm3LMWSEHSsKTDTViFoDqIt51ADNvIqSIpnlMDoC7IYeXnF1a4ptNI4W+emDtokXJsnO
WiSEdIRbV8kuJBX6CoJqrq+5CSthBKk14ItXQCz8GQJY3Kr8/NfwvarljjBJbHeqR8CA1My6aTDi
32fa+agmMKhnB/MYOUIOT9IAmoufdAORdGoWdBVYliPSigP2xFJiWuZ+S4ef40KEL/9Rseb1YXJs
+IergGMn0Zv/IDH+bmpMrWXH9fusJv2p+jcYF9gn2Ts62CvJpfsiu0EOKbwRrxk8YQ2vdgIxRzXI
6H2WJ8nV8DkCarQ204yyi6KERQXAI3zAzeMgzz6cHHHvb+3mRsgu3T8LN7F4gyrpaLY9tuAN50Br
3xeBVkmUrQs0EYdUYAQOLion6zQXdv3BXvgmt9J3PppUOCYssnm3WMS/5jpaRzF+6ycJNXF/AeJb
wfzx1AiIpMc1BQ7+Y3DqJNPWe5ImVGq74L2PcFDPsC9n61eneIkQnEdzlMtuTbeX6bBqWKrX0Xa0
Ihm40lvzqzyzZUGxmyR5Zxur+eNgBdDZ++jCroa1ZVem1v9nfMZyFu9MIHt268cpKje8KkqbAsni
Klik/cekzHmd553pge+bVqhra+tVR1qWtYGsv+OtEbvpswiYyUYhWEsWWlzGviqs5A2YDbp4hH5g
yn5SOd1nkSB/N2htRUim1K374I0MjcwbzTuqN81MoJZQXXLlbOKXPPyr4gDESS9L+zNO9yd1AjUI
P8qA4ATlKDu+qMpJk4kYLaOg0mOcTgOoRUr1PwOL/kEFDbKMfDL+rnSvkb2vm38zcz7VO7DcgtxE
dLxWx1HmHRZKE6P4SvVBM7brseLkCg83AoWBZpVwIsK3EhR5Ro0f3dggrm1yXF15frbcy4CdQ1Rw
kIywwym9ox93+yjQXB5Etotzxo6u7OIaibyXASSV/VQPR7c/KNso9lO17AJ397ImJZ3h95yYfP9s
Pecfi1zAR/+RYf1VTfAZKaCzGJHSHYrB7/rMaxzNI11l9wo+OYQl0GCyItY3y2mSRDIQpAjweoJj
h0fyYofr2g66U9nsBC9h+hhnpHEW0A2vu1hH1h7KIChcKOlVQxCjTI18/Ti+1V76eQQRbimysYtO
Es3Na6XVDKpUllEG9cnRr41h812z7H9Zvuxwx3/g0pqIY7fXbC8REZLiwysnUVuityfWnpiVhKle
WCflw8wuXJL1cZiaUGOh2dzAweqh5j13TcOHbRzya6J5Q6YZSWdt8zW3l3hkj8AvsYQp5d5ZqGVX
YKHXPRhNgdrp14JmtjvIe+E+fnXNzoa0LwhzYIdO5DnWWbBiBhdKheQWS7KXbK6Jy5eN4uIFevP+
eflDRFNbTCPolmt/+MImPRxySgtN6a0jaY8nnABi78GJflRpY3T1S75Gy2c5fiNioNi2VQHTNY/Z
aXcm2D/14SJDqEFM2T3lhnCoWwjBWOyZUx/b2DpZFPFdkIAvGppKfBq6gUq1awW0u7S25Yv6RkY0
gcBIRsjCdhfmcF/Z16ddagdAcsr3lErmK2wkmMhl0eO0nj8X7rZJcoPnCLB9eqz2PXSIcvIAL/Do
VHw+j1ykCzwmecxjOJon5ndseY7etVectj+1g1SYVCYiyCh9q2eiauoLht6iibyVox0D9lgwb+yt
3OpblPD3kAVOlFU6LVUH/vGmSwiDUJ7SDiSrhRSMmsgOl8SMbrqGGO6/FI7x37dF/QKqF3Co3ml+
43a6d11SfZioDwvGLi0G5O+tAEMBs3xyjvPsKWycZ8JFK8t5XW+MNArzk5CLuEqIBmB/1yVT10xc
QWajwB+mCC3DKIwDniq/WDOulHjNIeSXXkDoWBwQZCcBTpucFzj46/s1VFMjzE9XOQnHW371qvyJ
Inx3k18zlnP/N+a6zqcvaXogwkVUzYnmLgkzKBrFJA8wMTHDuwg8XQr2cZqoqzwUevwvr7/9Co2X
4CVubUUWrS3MseueUMCuFtF3ip2sx3M4zXQnsbrR6pzXeK75BlKCxN6EiHsb67o/cI6ciIL2dQsx
gQV+Za6LtMKvnZOvQepqX7e7dKeZSaP3RWd6zaVdFK9LseFqStiZVsHYvGFe+EaECas/QmBNZnLq
cmo4Gkxim7WJGqrksF/yZE4JdX/BcfHg+h5Pi1VnkuOoPIYBmqf2waChtovRomd0kb/TFIjljk6V
r/ld+yHV4AprzDY5NWKcN+Yr+51SdgYNjpErvZYhWnzIcgrEHMHy2CRiOuSbtER+ZajWW/f6o75j
1q9HywduXlk3KgrkoSfJe+IAvnaCT0+Fx7m/Lx9Cs77XGDZpOvZdNnqhx2rfACY8DwQlInBAYtD9
ZUkkEZSs44tKoIX/11X27dR9NPed1zJfaXfBwqtb2Ii3JMasOgOkb/dSEFlmqHz43rvIK8ZOH9vK
wXHbPFvgR7tJ4Exq62HQyoCe+/1DRomp7/urWvy+AX5EMhfkg30UrD7+kzxNgArJLs22krmHVpvh
oDPN2OVWgcxztmyirEnqDp7OSuYVyFE1oSDii1KfEezbnBpZjoHm/P9KzEyfhKpxd/R6Tlj4WXGl
/0xljxJT6zPWHke9oVymQSkKnOe/ELbBjaGjkL9g9xT6w0dtkNz6KE/4w1yPuTeXxAELPq6x4u5U
/PnisTn42Un1KnYq0XrJDjB6PSa2ZD1B2xq3960twHAiKa+MM2LwLD/5WXR5KHx03Lbm84RHhDoe
O+PJPzg8VcYy/+/p4X2r+vDAYtBlbHJScQEWMpGcPIhxIDn4H/FLShgzk4MkkIrAAEoMyqJ8ocQ0
jRKKKjT7Y8RIf0zBSRQjdG5wuRc6twI4rJBrR7JWrrgLDke3Cb2gpnEVPiaQF/i1SXriVvtLDAis
Io6aajOfaWyvW0wq4MKPMcM3VIWHUDZrM4ye5laPTnrMO4+T5439sqaFEekzQooodATf5FlP8zHp
50et9ySYhOVNrtJee8jRdT7Y5bp48ITneb/6NUjCdZT/xoCETBaC4lFKTNSe3naHjkpRejevT4nq
0il95SMAS8gjM4Bpiy5NCcbLtK/8QOVFyCKzzRXQdpI/Iwe8tjbV4jHVszpfvausFbwcFFqjzo4S
BikTgbov6Q5hFkQgEOpDzfiCKzf4J48bs+b/40MmyLjFnGsf0loA52l4t4JIYs+3UmADZaH+jzGk
fBH/cacxq1R64Q5Ai9cXNNblucKCE8zXVtp2vTvUPY2diigcgAfC0OJuNUAqdPvD4xC4V2zhhDpx
SPx2KQM6aofqO9ZnEegtnyFohnc1x19SSsTD2RZjxsnj4XArmSg88YkDxUXkLq3PdtcPGL+bXHPK
UCyu6gKROlueRM/8RF03hLrHv2D1JbyCGMyeTPpm7EgnFgoIGRC1DaLeFLQWbIkalGtBtRtyJYwW
cigJQmLd6YKpA4Qs5hzs6+UwDrXLE6BxD3lVqbXbO22/Sj5eRvgGKNZlJIOxGm7RI/AoacIYOAhs
GMOmZtFF/ekhw37HDiR9xEdl5rWcn1Q0Yc/GbL+CVUE8x4gBim805m18N9Zyp8JJJSWry+XvpYTa
ZhjQPjlZmHLNJRTiA/U5BqGlqIaB0APPXbwV8E9PYdw+EieEJX8AHEvpCs0pfbDvSBFKsAR0H2m9
aWxF0W7A+SkkG29iAWGh4P2TDAaE2EDhsBz9j5VgOkRYcPa02Uord/mBMrPnrshQZ6Jh8cqDNA6G
k3j4CwJ55OaTkExw2l5VXzqpPxzqmPH4Mn44gV1uEZ2DX87y43Axeoqdo63Hmb5hBJGEXSRN1yu/
Wh+djb7BFIwt5RNOzoWkU0SfjV4yivDbyaMUu48Rdm7nPr5uvSl1J+5pXBvLyQXf/aSz5gRG/b9P
dx3+3Q+IZAmtPo+/4cUth05Gk+1QVF7yOrJOjYXJps/HtjUG8sLeq2/0C4v+IYX+YP+hE/bKuMNz
UIGMiagRV/cORj/LzBGwpudncqjZKlA/1N4Ms31PCy63np/PI/3hOWXo2Vc5rsuoe9b1VVLi30Vp
ujRSHbViqr79ZoEUKZGyH+F6ah+1uIC5plaL9ER+Oi3eNbI3di2hwxdshqoz/4o8WJPd1pYRt7SR
XpBYWwHrGi/K6VVkg3gc1kNxDgxkOxDh+ADOr11AjwfjqX/9PaQ/kI4V+h9yzy6GeNionY2k1tYK
Tl6XtmC7ahX35oj0TsLXTDuvdIR4/5/RxZYFPpDqIOYa5CnXhZRjDXsLaOwKSRZS7WnKs2YZP2sT
k12YS+TL9yEzDSnseIt4TqiRdL8iwz8n491vLFgLWFQrQU6ZsZxfwhI83E9kfuQ4UaednvesPAhN
CEpeSwMtQ1ULlk/UOb5u+wqFd8sL2kOojnjGcJzfIAKSjmOU5eGSW7GV8PkNnJAQI7vaUlw+f4Pq
Zl0auphwlg14ZLWiOPwMWfs3jCU/mTalnXRrRq+DqnyIPkzZI7u8LYLA9nX7etkrpQu+q6/75J/u
27PDGYTn6f1ZgEZfeAPTPwOAMoYYi4/MouFN2HTN5aPeCq+QG+nY+vOLoFJ1tMzjw6Pn3M9zhI8a
6ojcIcLegD+P1ueK17T5SeQdVEtungrO5FhLZgmA0vty2zMJ998OR+zlFRPgZI4Qt/ME5ijSbXRG
ly3u1BysD3gPx+w2bbJOVzH/2KMMKcNpLlfY+7+HO3jX5IGNqDPWGNyVey5chJ3iguTWzg0HEfy5
27wkhWMkmCZIEgG/LFYjN7O19B44Vi35OcKDu3zSrBsFeCgtXw7le6lsUdBf70fgAHgWHXjohM23
gibHrT+27d1WRWoKAqJzxgVuaC8MGV0IDAtNiJHK2bKV3LyUSRTrRZ9qOv1GQTeAhLAIAOROoWGS
8caU4pOVVTD2MQKLqYBOyXgFG03RIB1Rf741BXn4K2VG4izQtp5VZQWJHRLYRyni9Nm+VeGlbWVP
DR/VPkaUdnTF+AUIHR8lE/qhAHsqoInvIfuhjBI9ER8D4SopzNTr6KCd2y8KTy5GFoV0AwOTkgBX
NANpVRTQkCMfmNRIBsOKhTJxbNbDvzD4ODbk9FLwYpH6tmUK017hBAcFE6SMhWazKV1zs0/HMJT6
9dGaAP1B28/kGmvaTA10za9EdJUAfq2WzDuw0/cf9FMzo+9QNwP2lswV+EXYrD09rxbC68MJy5p+
qPZMj1cKXfgegJS8tpLcB3Av9cTVPQ2JLjKT9ppmRA5Y+gKnDFg5q62dqsnqZsVpccOO3sWTUH5D
SZpi21ACV1ieYqJq1HHXVJjaywKs0sNrHgiZb9DSqZ1Ad9FvNuNRVRJf0fisyjRQEPBYrLrnKr/7
HnnviOgtFNFhPWNV5+dbM9bTXZVl1uedhbQxMnXe/et/+w9vcVTd0P0XdnKK2uBOTOzvpUpB7y90
y7sXoC4Od/LvfKw1VaoKMal4MvSeSwrMMJ1ZHjaJ+6RPBeEVrtdKulUfGcyBrqd+InexT3E/4Qma
KOVkcI3vorYrQdMYMBfWap1Xv/gXKPyaY5w0sTZvLWNNXV9IIBxQPfPditFqbsmHZAvzleU8AQZq
ffcXwAPAEHtwINAZ4Aq/0goQOLRtrtzeA3j4KP+kpA2CjeY9wa29cf3yAM3DIlrK870LwEVtLM2r
WI69QIZNrYoZlDUt8y6eCsu9FuOOB8oDLi9hmCM83K4oqRjYgEJZVNCCj4u4jI0/fGjfpqCdFgud
XgUBh3BP5tl7dYiq4oLiqv9HlbYzuO79kpx1IgbSZ1wJpTQQnt+eVn0UbqEE8ATqGPTgGOiCC+UH
W3vcehbChdyfZes+K+Ka1DMTvQVriqds1+9P9ycWpm5TX/GvaHaNqoafND/PtLdDcHI8zjlxEaTl
VRlWISZdkUp0AuWoCXHkDXQOr1dfavBjiAEWWRp4FbaUmHb0AR4UQM2IXI3ryWmLp1nYilbnqQsA
Tg6bOMXK5A+3U+aRoiknNdbFQbLsk1PK2Uz2uhUSqr223IlDCYmEu7l3KoKEH1vIzzfNWaK6GpG5
61ppFmYwcd8kYpocAJxbM2znBZy6Ttc4ZYvZ1S+8CZcPQsHCYcEa7AqOy4JnOot08hH32KBKgqqc
gO+PrjRxxpKaLnO73vnXfXpYsvo9P0mCBrlku8kZarb81DOE21J3paFU8BaxPOwCknMLFGQSksbN
F12WtdtiumhT9Io3BKsoZGMIsr22Cjf4jUMjJsd+IhgXqFraCRt9yopN4O3ekMTrabMfrsWJfuZF
I7DNmd5GWbjMKi7rC6E+bFCs+4usT2EY9w7nVtMz8Ozq/PbGcs+6Erj0ejQROhHG5WNDA7bKhZJu
wMRy5LeadH62qm67AeNMIFg2jHvub5aYXqJbcCkjWKXt6EfQlTDygrJjyH6dVWztVjfibJjORsgg
p0Davlu8li8g/AdUsBSBdXmNB1XyolSVwdM0dqYiE8g1p5SdZ5DaEhPm5V5LG2Txm2Y1UDGgNEEH
kkaU3fBrgwI9ZZdXEnp5NGBtA4aAMZovc2VcL8xX8QssAnxK05mHDz6WvkoYEKrmkdgW7Uwjsq5r
LlHVNBKx9rAK90dM3eR6pDN4AJcrfF09yqQyoxRdybWXhI8plEVxt1F+qMdPWkw4LCZb42CleQCG
HzqVW253UCC6aZqNV9LYWjDEbjhdIph/D8dsMZnrU6dIwT2InoG5G6Z0Ol/Hf63IusDyE2aAFSUy
dx5DAnvDn+cjXGYTuuLqv7hYpnrw8FHqFqd2a7/mESnHujgMvL70NE8rMj0Av6E76ToOkJuMxf/J
pm+/LZ0aQnJHO+HyRDd1Hfk7oMmOIdoDHYv5f78w0BbeRXfG5600jFHnBfYXygcDAxgVjpmn1QEv
iMl2Rd9tYGy+gmDp2kG/bGvsiLKjNmUaWHO6tdbqhKhZ71aCYKN6yBJ+NKii5XsqVSg8surZbnIc
paVpB7fMxjBAU1aK8HKKo2fkmsJUVmJ5FRhzevlPus5kgBaAJWUJyzwGAvP73cXlMLhqvEEfB7xX
w+OKCt0flFApl2Q64CJHTgtafVwsBMzfxDQYYUl1vyvOPHbnwZlekaAqJGqkiFvhuHM1dNk1qCdv
seGGDWALATAQP8DfUgYBzOsZBbyjj/YunWpGtbv7D4TP/9qtcxwUz+h4/aJHwR1PbNY5/T+rksvL
VJ7GJyNdyrDQHp9I+5T/A7YFuU5Yshs3MnxIaAt72S57Z/uDWgf1+9p0vgaAc1I1NqPbPjdyRQ1f
dFo1uKuhuh4WbiSrSZIst/5klGRZ37hvaVfcO34aMihrJDDJcx42ATwVOgfK9vTf3UyFWw3I2A3g
/TR4bIU2hBDccAyrqqnnQB1oJ1JJwFLpWywGDzbmo6AbcYO8A6bnUq7bEfTVnhC4WdDfW4f2oNRf
nbGl0dDjH0opuP5MzA4ihtLfAOMmqgYJgm1KXUgExtECZ31UnOTcMOLlHA45U0ypYu0B7O3qaCQQ
edNMdExpLeJorM9uq62g6uWgjM04AbBI//SVRFV4Q017UqTS0y5QPW+Kkie3nRBmHnNxBZM01sZc
zNtVaU3N2F13iYY4oCJfanqXVWm5rtGssYKESHoMo0VCMkgLPeiHtZwGAnNMhE0BNsEEGjah4AiH
jaqhcdPZh8aIoHaxrpKcUI+VqEyZKOx17cZFDV+Vcz6otNb+ggzfaCM0KzNb75xcNGbC13KMcw3W
Z9RwGxYxQ3PqJKv4Z3mXLTAMBxy9vtD5hXipHdMx56VY4cFXsfOd+5xNOo6LxODx52cpQH+LQHiz
/DP7JxX5pkPQBbAT0cc4WbanJBpH7FOTdSg/z9Dsby50Xp9L0s+Kg9DpUEP6ucAr7Jgmnmmtx46o
oAnulsrNBznTa+Lfqo3KovtHXEAhwv4kyh0QDOZLLihcJwJ9r+btly+0jHSX4rsdlnAoBG4pCI0k
kPMCKgbKN5FwH/FWWhC2ZHKrMRdNCTWqo1noudmVaq8x45tVYoTWu2ak2MCyIi3ug3uKmpjas9wn
JuXDklemZE2hzUHgcO/khbC9UYO83LEJehSrRJrBfCmkB60ttrC1Amlvb7DiFKTIDI4R6B069KhB
Rl3foOryXQoOIMlBqhzx8ZnQ2ZaFkRFQ+I+dYtiIQTQo1Bxp4gbVlIjz8d4fWEeaTgvDxYCH5TjI
iS4ARdPYlH9IUB9ayavrqXfBp7Qu5q6m0JObNQdwNqxQX7S9GhszZl5XT5A7fI04gWoHBc5RdX8F
ewk1zMg8RMneG2E5lvyslkzh5V+23helj49DEavlrokseHeuroQ51FoFpy4bhVcBkPfTM9odCMFM
ObrjW9sXoj3Nx/4fYIEAojhP2bkQLZdbsMU66537GntgSwbyy/fM8zZjhva3bPxj5sakKpbNS/kp
2wenRHnxkNdw/5KGrFPq9+T0z8NALN3WhJiYwwXWBqEv5L6GGKmrtgtZmSpYN1xBxe+fwj6OroKQ
/D+tid5fhBuhMpldtjr7+dMMhk3sll3/tOXGO4bx7thSDXK9dhtOItrY1NR9qlXqFd4/iaG/yBUv
GioPogMKwmhfMNDvd54S5iTkNBtsZJrCsUr+t9udHMeWNX4TYz+9NshlsF0yKCwPLL4Bu8Y/ZPp9
W2Rxuro7KylLZWz3Js6gkLrhEIR4m5jtrnqAIZBwdp3tAHJmnCcT3NoCoRFNuulWYCuAY5EZ96av
MEOg/X7fl/TpM0KXdmWGqJ7AkSveLNxGv9V+Z7kVluCfQaduvqD8oF1Fc7LoDGBqYzZrDKtTIAiW
BIG4qQ/MsEKxqiil7k+ff7y/OXKidY74PDBjLa0dHPC1TkJ0helyjJohztR5R13Y9OdALVrlvG+3
VUK72WImZLkO7nagsomDeR5xwtfaLnKncrxoKMm19jSkB3AlvxyoXgPxL9ZsFwZOghu21fic/q7p
MRo1csTqF5vhrk+eKk/L1C5ae+zzaGnx25eWpMpeY5klnvue/0APrBMu7SVKqOeT5fAbmgXiMWHr
Dg4eWmU6ix48MO1+ZBpRLhjOjKlJIbYcpmOW7ECDY/9FnZ9HNIxvl6ApVNUfCqbYEHDl/U+ac8d8
BhkFy8nLt2fbBeswOI7HO7FU6vxD5has/wj49gAs/8b2LPjRsXKPMqbptYSrjZLiVyo+J1TgDn/Y
wv5mbC2DeonCSK9gH1BYXTChO5MnrgingJhHeEjEKc4VCTXqb3B7Ex4DYe3c4uPqTcqvook683RX
lbsNJRoafGwPbRjOsw2BjvrQD0NMwr4YZkGCY6bgaZD0/KOgwU1GAVU1caU14/2+Z1Tmq9i3PKr+
FYiP380oqqOSm54ZPScAO3d6YKdQs1gFTsOHmBzjiT/EBybbMYao6vAw91cI39BR+bfnOMcl5s/4
8zprfDkQ6E2VgJU0g6ro9hwbPVkhaNzkNVat1IBMtUELjcEtlECJBZxRKFc5hzSdje8KLJzQTogY
/j4nWv0PKkU+lUTN/0rpyf6aDEJwvFtuYVYUehJ+NM6zysh8PL318UkQ9VweUntz+wYLHFPeK3FW
LBEAOX2Lc1EyvtEZwuyDkjmf+CPA4y2Lypqst5hgMb6GjsoRSCzfJR5TBG4ZXjsqTO0n+ArJBktl
dyZwA54fz469MUJBunJ1zi59KJOXQ0BfA/+C8Bg1rDGbwv04RC4NXL78lhjGfR3Ho8EdpxuY4KaC
LcrYjoF7fn0ENB+jwe5BmmFk61v3BcR5s6stzGf8hjQdwEybXxAY6k79MMHsrFzkrlCMUoFOs+oV
e2wTvMyzWhIJjPmh4MVYX9KpMFLBB67bSKrNJauTX9NmMMAzbPh8ghVz3ulkpCrQGEWUA/W2kP2V
FBQnfCzP6bg91dMaUe6eMFzK4aMsF6X6TzB8HUXGliNUvy8Cq//X5Su2rB1BnGckvpukObAeYE8Z
uFZct1txSaXeKtkEj1u8UpyeWkxyeUP4KjNxPAHyfR5Oa2k3ERpiFInMO++0B0mNOPZTmMhACTDi
Qovq8QkQrxsqbbssxvwaBi+EMII3lHUfb9Hs6trEvD6514n5B9Xd0hMTZNUFoBDnNX+pQfihSVUu
DyquNJfem5MOFWguI9j2uZcWA9gKkuH6Qn/7diEf9ybhxonzoTXuF/z5u9vIhHrrFhSn1ZeKBiV9
HYc9NpF/df9OyuyG+4KipM7yssKuV2+8u/953eFqPxLfrv5BfMepcWh8OUwAi5Ve/gvmCVSUQHzx
/iuuuJxy+wkKi8EDxGLvFhBZ/liwTrbDOxeTLDtqlq4Cus/w165j05hjeZ7Kds9lMqosSNw2G/K/
mm718moNEh+k4aVTJ4Tu5LIWonog8aAPbG6Cur+23deQR725p1cYLjAZTa2Ifpz6PPv3wYzsB/XU
bn4kfMK7UBs+1S/c8DSL3BIHUHZyGsk3pzMmGxcWZmzOmRcXCVzUkx1rfNTzWmGWySUNQbr1EQOn
dGBu9Tk91s4w5OSMsH7QgC0qnzm4ltC0Hge6RcN41wIlzD4TQH8LfjbEWxbtpBipPXvq9y24P95/
hEPpKG7nD9qcHzUH9kg7pn9AOTrLqNWiM5Bw+Wjk9TF2xGsLAzgvoGmH3eQmLo1fCBllEM53VPqV
AA3muKiMusRE6un6ntc8KLEIz1v31ZKvyEWOVmaNWnAKeiuIAhidSd21nDHam3zqLTXeG/HLnzaZ
qI/x/dEkqo3FLyiDsq/KfyvSDB/1cjuk3zAHxopz9i9Ev1AtVa6qg+Ar0vM43OsHvfwx1PujIO0x
brFTDHl73oUlm0FrNWDaBtxLEtUNSeUdccxbkhZKCAXe/2T9aBVdR1rYQmPTDiT1VaDTGzcw7L3Y
VcTyVNdRTifPulac0vG+DRmkFuX/43jzUPDsQRmsO5m8ADSLLRn8Oq8o4w0jFZstIStpoop7t/ax
7RMgAdydEfPRLz9mLoDC+0SnB+geYiwVuqa4EzvwHCwAy5r1Lu78TB/g5DlPQiPH1l2a0jLDWpoQ
3qmjSW9x5M0I7SVC1U40Aa1etdpkfyELne0BUtI3TqXXtxy1t2lK2NFfQUdQXV6j/7vYV15sa0sS
Az5DlnkrdP66NUxCry5fdhPZ7Kptbs9DdFFkxtXxgp4ngAm7EWfwSY+bzgVx6nj9wUiYgB1H81uB
evV1YmKVFhzfwHYW7CpVmpKALniDaH4gWrgOjrD6iY7cTvfAPI4+S3NeMZRIY/TzIctQArYRHLeq
BuXnUm3wNurHRLyg3z7iObSs+JL/Zx1/KydmTNUktwFikdsoOqcM8JRi7nlzOvkh3wuuAmwjQnrY
Db2PFW6V3xIGcVX0RR8oBo6+Cl7s4OySKKehHTSYgkkO01aKjWWG7QNQEu/Gd/TB4Cun9rK5ub+p
rZEpVq3LY6LdenXyvgOlkUIbya8rwC9Ca90VSE5rU9f2PoZ/wCol7zpzZX/n2nlko+jSDZdYhf5S
BQNhtA16vABl+4aLDXq8L9nCIRBd3AM/qljNpstD/ETD3g8A4yUGj+k3hvjinh3AI+z5+rhs3+rC
r6jVg1qMVK8yXWGaa8VlTkcl62OwFa7h9IDL1UnjY1ae7WiBot5mq0c6tju/Tr4dSruo2pQIduA6
adVoiW2OcLPph9NJ7FjRV2+7yl3T2OlcazyGC1zpH5fsGRjLV67yF+4RC7mymaHESieVjQPrFaqK
UDMwsy2u4tqe5pLNSF1hv807wj6rIhc3/30ZbO/CloOPAPbwrB2wrsWp6/aUG7iVgwxKiv7CJpy2
xbLBFcYT73vHjiwN5hBEpp2eu4MpH+EooOBxhR5S595uCEQxpCUDwTufrFRkaLd7YyeGu8//vMP7
E+jtM4rq5zSC0/DhBdEHnvRLpc41bE/0g8EeVStP3EFxvaNQ+I2cPXPkpHGUN3aKrq5EK1qfrEXx
bhjONuOGC+uTz+AUkksl4oTi1utUcOcbTKN7GxWftKFk6eeGBOm2AhQCjxQVSqtbaIf+YqbpP1PZ
8vkux6W4Bduk1zGgcTTdS20s846xxovdf2yPahOnRS+4q7J+53KzHSepAd/R94+A7NGiGfWwHNZH
zEBQ3Q1mzswybuGkxco4glJS0ImrOPwp5eheOwa/X8D2obRdB8l1OlGpZMj2HhrQFlkDXJM1MlAq
DX1kf3h991cA52f+hkCfMzAALNtXK44JbDI4oBlxZiUC+dMvcRSxgNBzsx75SPh4t0sASzj5ju+r
vLi58K5tQ6meTr9KSiAL9S99Eyw2Mj1boO4sjfQ4xLOY7yllex4DvbztmoTtu6Cg9M8vwyEJqNW2
T8MqW2KTFYTVYNDajXdwirAsR7OHe9ROcAoN84pvPZQnvVNNrTAN76WBSX6tG7SzOFEvFGiR8yLg
NIcYhxsPpCXllJ3BBx4yXyYg0KDYZYht0JJ5vzjOAidK2nLO6/+/sYvjWo8B3SF+I+tifreFmO5E
IcluemRtHJzWhFZcZKRtHdSZFxeqD17zQYlUgVJZt5x1suI4aURVAuIgcWloGHSitLm79wTRyysk
dmVmint5B0hv8h4RyqUnlDlsn95mw8yXRzb1zUYn6nWisG27LdoyLm/EW4oUCtgTid8R24SEhC7K
7QW94gSx4zeqoML8HoSnsP8xTlXhXHiOCsSHtM8HvAMAY1To2N5fgmGNnzcVYYjgqFa+t8cvFJUE
LAfBoQ2mWBPcxRfMdWDKsgRhK5N3UIbsOuIJN+LihmlZcZmiELp/D72gvQDqgnkXnxTH/1AwUrWq
tV00mULg3h2n+gZnNkQMDeKS7fsNxUCUn+E6e7ND05iv/kX2Gq87ot7lb8l6k2DEptbzl1ScJATj
v9WkWjUPYj9jLIyhvCKZz0uK0CRm5BoO21WDgQFSiBNhicOPXp7K72cwwFyBnkturCalaQGzZHUA
qS56eozwxp0TVg7EOGtsrJ/6KeasZzydVMntI8gA2OooNhDIuJ+R1tHiijbGo4IPGBsdR75YKqDm
jLSvTmykndHAWiiFpZxa6E67BpFOXc9c3EKhF3jYJfNrV4Hv4M2sLRfFarff1De4tanMpMlAd9tM
SMmhLU85sMB4Guao6FOtUhtTMua4wAOXttWJb55kiUq2RybJwC54tK5HF0sQRqTPInfY5IwFUIVH
I+Sl683KsL1/hYxW5BB8UakHYzXi2DteMFzaZeT0yR+YYvbj7YS5L7/WeAJDhb7gFx4qxyLwVl6c
E1KH7stTEeV9nt0MLISiIJLWxIAxWBFjIauNN2p1ogxiluBpOgXaSpme/1fbmuSw5vUmQswjbnuJ
LttK//0kMM/fPrEJxXs1vN8Yk5Ky/XclrE/QnqYjcy3XiIWyKNKWZAYtWpK+/6ISsL77gq62ZUfb
h9ED+n8yVIjLXJZY59G2cKaqjmyPoLpq4qMabFTVY20mC1jF7RDnA+fuZaGml1SXK9IILHF1+g01
LZz3ipyqW3eK+fww/prVeTgKfWf1jDlvNS53lcbyCxl6B9P0eUs4UYZHznCQkass8ys+/wjTEbeY
N8RpHc+N8xvnU7kkc3LAsYGHVGdPWfbxMk9XOstoD55eNiXzwLWySTKN5cUELUo7MnYFBvZfvvAe
WVVQarL1GZrs4x9hqJisH0HNg+5OGHqgMuCLXxiQdaOH8lsw4Kqh1mIUV/x84Nk14pfvGray9UmF
EAKCjfUkCr046/NMsPvlIWtaxLMnr/jb6DI9Ov+QC3S4CX3TdHMQ6I0AQtYv7G5Elrs5bm7kCB4B
zGw++/Q1MjcJIkZBJ0sXqI5FrVaUYh4GwVu4ADLNQ/Agz4kGTypOKBnBCJ0KzbqhfUESfMFTIxOk
eYNIs3apybq0kKPnmAeSvZgdcp5O5tdjKK9NehJZ5PgQvXhMeCDsmOVGLXsnce84K/5ikd9Z0nBG
bzYUdb5r2HMb5KM2+bqTNQhF6cUSDXXKb+W8KbcHC8S/5Sy9z7PVXW0dzQJcKwF/ZNJAj4yxjUFi
lV7RRes5804AJjfRGr9eCV1DEAz/JqiL5wbe9mdrzUJJ3SmGpGrbA6JB/GpMCAvKpg37aFN6Uyuc
GjoBwwEXogymZYtHYTAZPcC8fevcfri+LlTHpAoOAlaqrYC49N3pgcVsvswRJ7c14XTNwT9V3m/4
MY3uvyepJ3gkAcw3IoouKex8FfAVeI5Na3pbctxQ040L9zVHgKjRZ3IBR+6YoEriqBqU+OyNSmj0
CBji1CNz+XhoukY8qE9lFuv0qIfP3uaANfAxwyPsvt73NvM5FsfcwBspP1ZMyhHWQxhEkqO7jO1V
hjFg6rySXRjRziStvQTNdfz5M1uGWL4EZKWatcNb1n8p5hgTxlBjyuqUn+G0rGC/FnpQsCYS4neS
+6KodDuqiQxaf/6UpRIwKpsUiW+4T9GC/gp5gkwpDvGmJM0onlIazuSuvh6pz2z0YY7Amu4vvHO2
qMbRuNPiGu/hE2RdPgn8EvzxGsHhO/HPkJUG9gn7TsGonDUuLDcg2ATfhAJg8XD4DrhYzrdEg5BF
eooduNwzcE7xdoo2lvGuXGCt3tXMRaSQSDzgY4IBJwnApjNP5wmuroPpG4yCHpBgf2IySEfdivxX
cgy/AIhEYUrjygl6NDLnYqGDoALLoDZFEnpLd5s/rho0lTvjjTakINHB5sv4xNS8PgLz5Yb0zy+e
6B3XV0mtOzuJa5+hry4+VRcAeTUFSZNYuAIAHvzvaDU9DNiDBI5KPwGOYoJvhJCr23M7DkQ/Rx8S
kFLKfmDdb7aP7U7vfkorGFbCbchhODkXnCBprrlhWoAOyde7vv8gkxcCTd2rwvyqyrVHE5+7F0/T
R0YoKkduu7WJF9PaTllz47ovAH7uJFZfKc71tcCsXgv1uobLVjktGIK8mSHckFN0nyYr7UhccUt9
Ka4BxYny9yecPlJ+x714DVm026Xaj66RDy5xS98mdLHGm3SKIwQbxRuJpQix5Ai0LAUsHkxGyzGe
31/Fyt28ZXJM5dbgrH0eH5qbKlzf5WeR8Hel1IInhR2cfXEWsBZYthrhIhynHRofzDnZAAdsIvF6
+SVbyagrXajoEEzXSE+MIJgXiijEi+li/8sFtNPUug4CMQ+mW9E7gx2wASXu8ipOWKsnmkKf3IFt
GFlb4znB90sXsUxgQ1BHGPP0KxzT4wglAyRX6tWj8pTNSicdPm5hOv8zGVv42YUJ/Wggo5h39uyy
EeLrQrdrzWSVGZeH9/nMwPARAyHg+PB2I8Xmi28OQecMttSddUTqIT/OIeGx5XOfTKysdLZlVHjS
Fqbr0QYJVrTp0dXo6qvxLEOfpSEe93RGR/p2KpPQRCUa+sA0WsxXDHa39OXFKx2cQo+vTi/U5CUI
kpNeXhGIOrDo/g1MUNhwmWIasX1s3X9mzHLtFVUhmBzcetNAUU4WQO/0Vxn8HoUeAzAZJZKhyWMy
81kNOEGiB3aUFcnG1LmwR7fKTeZjqyFCR5JgndSiXoEKnQRPDrQe0eY2NzYIjjKZ/y/Q1/9twqn/
dPEVo4HrsFG8a0cJUSdp3tMe3yduAAak2+muhrE7XGmNGpXihRPVW5hjyCQBxxia+kI8yjwTHCf4
eq2Vmpw1A1sLuth6DBipbTX7TpmerSeT8Rjx0CJrMei4Kn4eisCJxPKUzNM0YJAi+JGCKA643WFR
ncBpPQ8UsbucwIfUlP/y4JDy7AxXA1s3sCBBMCs6adFOfGpzUkElngJw3eYPR+EhH7BO3PG39C/9
sMBIWao/V7o3jIB1N4pHQdJlGVTSxs6Ywf6/4X0WlkLW7wwwavWX0hy85m1JGZd8MsW0sRTYcPYR
6Q0tR6864Y17AsGJoNGynRv3AFSZxVQOF3R6fOWl50Xg226dqcpRwSJgHwBEgsKt4F2iCq06fHxV
GihkaymsoJ7SopB+sKgk7myYzhwoLYiqW6JU2SQoHrz8mKswcxpcbe6jhzG2665Dx1N8DYBY10b+
rn/PMIXxoKMZe2yz+GT9Cv56oPVjXD9gFAb3Z5xg5Du7fEf8em55HZimwmROwHBrHR5nH5K3Occ/
OmUb/aFN1+DUWN1W3QNED7uUGnHWgyAL2DFsmxzYpneGStzcZh5OKeiXH5Nn3gdfTukgiUKCbFPZ
YSpZGxJF/7HijhV3j/YohhW68xNe/ChVPxg+GXiFVLgOQZaOwFqn+ibVtUVBd+73jsB72RhMFuA/
Lpz/+k0wp8vLoo3E544PM/ZmLmCuXpSzVa+K4JgQyjpZbXu4fJumCTgbMxb1oRD/IvKfNpvyIddK
NDq3jHT+9BOmJM+Y998i8yMyBF5ZEUNlzmjxLthqydXk75GUqDkG2bamlg8fYw6GHZ0/cBcasyQD
NbBIYWU9kkuSBd5DV08i7KukH+VbDToqbdVgt/QccPts/8R/d0N0WtPgZF+Dzt1EUOy78Ag+XqgC
hXYThKEm+DAy/DrvVqgTz++elaKoA1qdw932eXPI7hjG2qIaK3Hlf5gmazcmHqsNpwwOEDdTY48r
IU1YD3FkIOGidOGnwNjslo0JXdxj+sjJ1dGC8JUAm9DpJNMxCyw1OOM8ev+/YXSM32Opo/lH8SuL
kKv/Dh7K0TA7aQ4SFj9AruESSF5kxnPJO2q2XIWVuWRb0v/p+1kU1483YVg0AevIxekHM5GEjc7n
Q1fFL9IjxW+IOL5Ql3uR9VDfILCcD2ndoluMDAGi5DT3+VV8iBI5nEMv2CWddtEYuYr+XdaWHkfw
3TbLuH+NLF0iQ35Xt+nHpTHMkkgloPAmxXoa29ZMCZdFUqgqVwvQVpaoh1ikSmWmOcqLgalqKl8l
1BW0sl9sSyZxHPSYexsmgdburyzpVK3s32FA7y2J3tcNJD+it0sfKXPkka0An7FiW1Dor9lsn60z
NTN+OHFigCIA+QbVeVdK+iQlGIaysT1Q6G3mw7jnxQFPPFoH5PnyKL7NbD2p9aafglsskchLBE4n
uJcXhBInd+NG4TVriXGK5kcXltaEqLDqsZNtBLYoM0C2ONQoxJfuK45P7NXqq9MFZVD/zF4A+Opn
haVslfLIzCvRyLecemtAzj+R8R10vAQIpaztNa/eRwngB0QaH/LchJQkQWOqRXoEVr3y5B4gzbkX
DCb0zGFNW0PLaItjL2lrlwOo+IEgHKSh2yQY8lF4Nd/PxpnhtrGaUUiS56fZpxFlw9uMRZE6xDJI
ru8JX9xuLHm2Ub1PexRORlcPNJwkibKVS2cHQUkNRxm5XO56FiFaMLpuiqES7lBV1fAfuJAIwxnv
DP9N1jDZlFw0ZImLh40I42vCtyZDzAVDZOb1ufQn/2cKRqpmFRhjmgx2fnBK084pKAqAlWiG+Un1
HCsq7srlg/D9CWtM+oJV+Dcyx+unmA52zqwtWsBQyfyqOraUEaMdrDWV0nOie+YVGFvWSgyEeMzA
zXFBlPgwNj8obyPwoODtyKgbVzntkwFs6SsTuQG9QFnIMc/dY3q+ltE8AXT0FYNsdacxGsoCffFV
fdvdVk6d2ee78ew9PLQXHNIzsPOUgQyB/15w1c3AAcNiQnFVo6JfsJ0TvCxK57xoDW8uEmPJqQEl
4AVYfySetO+3xDFaKxcvm+d/07F/1YiBSwRjO9yWmM8zYGo82swZQUakFpXksPLXydzPgKbJD/2L
hTjQXRJ0PxXmC+OD3jDQxNqsfPoYTU2ZhBwt6iF2ZQgTpIjuY9rHsNiNEhTF8c4pKPHjwG+zWPie
ax0PGo1PxjtpnjOstGC5dCj1N5VWRlqy7q8KmtiRmVb8nFEDm9w+kTXzDpVvJ5n8Xa4ouOCGR/gG
DhCZ6yABtEWq2+4Iux3oy7tmTck5IQWU9qq2ATWjHkW3BgswdM9jtIjoloEroct4/KG4aMM/js6S
z2irHyq+uR5Tb/XNdq+fZglkYaL9CTnxca7MFyi9i6V1UAiTEQw2iLcQkNYq19ZkVo9INyV2N4Lp
HurMqbKtJuCkdmSUpOYsmevRnUAu9X0vrJMu50LDHWKzQx3JbUg84RVi44jrXwnWJb2ZMzyRU6VQ
4XdFvkNZNwDi2+0M82PvQkMVL743D+k3+l6Hc4xvW9f7mx43l6Fd7PjAJlS/9mi1eF+k3rK97mGR
8rYm3QLJtSd6YV9Yl3VNS3lnmYLuBkQn4voC6wjfMuy0azgqD2K01IYkEmcVGpspFc2GEyicUEpy
Ru6tykKPC9LBsul8nFYDItoCAccm3WHxKHei/+Sm/yrX0K3b119XC4ksdoAUKkPHxuwDeufRvyUf
ieibomaVVYqQENH67fKnXK5Ks/nVCvZZtYjcouYszmD8j8qs0ti0EiUwWqKYgONUUCg0x+3wAzuw
hMUDhr6bU0K3/gliEGLWaGTFSD3I03+4MroB5Itx9WyyWDQoQgTsxkOfFwbOMULuoWKZ8M2nSJNf
+IhkivJ2COm0WiZ7/LMXJbl27jVC7USwQwMglbvyvakoPYSzSYED1xfXUEdC+uywXBvK5DPK8zjp
Wcm1I+zWnvjtfl5dndKdAcT319YLbWuApC94y6r7jdkHwzQri5CMmre5maapS56gftxfdaZ9qTpK
6uRcVXdzm39JGmKu/zD/6VzSkELjXdn4ocCIoGxC/vowPdZvWm+9MN7QEfEjXNr2L2SlKKAzTdpC
419rafG1vESWbO/Dq84YWfk+wyyeUoKy+fLxqOM6jzbcmzPAFMqWlVK6F6gimih3A5+H1zcSDb8X
2lls/OqLrVz2YlZEOBtE2I7Q50AoTEea7lYb2J9l0h3l1FcT3+O4vzE5Aa7/HE0A3N3iY/IGqkXA
Z8Q+p/0woVvFQLUvcvqkGLY3dUpFRXOyXBBTPLXIKmhYd/XvplParZukc1MgNAjtDodQpJIIdvV1
kAWxbylYGu+mZwRzQWCeVjsBLmA/lMJYukNaI0fTNngwnKsEGW6F9EH9yZFth6E7qoBheHgHNHDl
D7jMe0zSTXjpRcsAP8SYhxtEV/sXorTms6FesbRLrOz6et4dEzDj2OuCJ3T/nW+I4/q4Bhr0Snre
khFgSCB74R74VrPsoDfs6GUP/hh26+81hPKzJ7wTvRzmnmPH6wkIlNBehz/sHpiUMXLhTkSDmtXf
S8WupnOgZdDfvJ8DSLr6eYc1g8ABoO26fQIzFuDyg221ZgjcXNVLsXD3ZOaylZZtF9eaXme89Txs
A51sG+//MnRy5WsFYUpnWsR5Q0iFFb520n3xSb2yLLRvBkOBi3PeehUjVbtbdAfO4Z+mfNk0+u+N
WVXnoTwsQUUlrMBz8jqhZkp0kr4hKpNmXT8kBJ+CyeA2t0+Q8Ng8OjRfd0n7b/lUxGjuulIRNZfQ
mrLESN1DmL3xRCXGTFvvdd5x1jLXsQ2/WxFgGGbjBZAl2wEz1Zo8btcyggD9HxbxfdsPtoANTV3d
vRzMC6W4Ks5zKGXLRXdz7b9EE9e/2E5oauyYzID9z3W9Eh+W54GxM6DGSFjqqsivVQ6DINWspEW3
lUMBryBo6sohmJSmpmoJkMA4D6hw+csMRqKBs1ZjVqZmrufwtNqNvDRPXvVHY92DuDnKTiCJGJnU
gUTMsyR/wlXhMzFFaNlC6P51Drf8IJrBpMpWlfhZ2evlfYuRsu/SyvCfOLilENyyPZTBmJGLUBZF
gv3jDuZ0gcMqdmffB93HI7oKU+T3rVA3mHLmUadFV5uOZ3IRAHIAPr6ocn8t13477j/xzen34Cdv
L8JDtaC7MfNMyddc0eKSgWxm2472wH7VPjo60qvuIEU5NKLDAfOgU3e4Gz6b5KavAq70dcWkeRSw
6XeZn6H30EBNW5MEXwwY4aSdBgQHLDBsrsGbWOgsVnOFCO2FvJfmfoMNjmXzCU1coo+Ub8mbVR0/
AjkvOUy2ZZPH0mp+Ty8xBLnu9IZrc7q0qcuuahZXik7rMusQGS/LdtZ9VimvWfoG41m20tyyyU3y
n05lENCZ8h+ZcM5nLALubcFb4RvhziR+9ikfonNfp5E2nnIR2Pbh0l1C1zV/sRm7cx03oUI0RnZ3
qQiy9jT3p4CUJyrkt3ZlI/vsjjs+FPirxybBwuUm3FjkJ6GdW1KCAV6v1JZLHeE5bcGOAs31Bks1
vQ7UCu9aKDS+sNenBAMfns/C/ifZnTIRZUCDrwzYZmnk8yTqOWHKjHJJhT8JH9daDeW/RzfEOsLE
CKo2v2K4wfugkI43CfLdIc9ybza/X7sxfazTrY5MHW2aD995/KOhxrzgeoqU80It8ZVnW+nHd5kl
9npbWt0i2R8EOK6EQkFDQxk3ohvM8WE7yTAh/NlNUz0luQ1dV5DgzKiBGJqbtV3+IJVUNsQmevvx
XLPdCWFk9Zej/MEjeahH/LuEjTzYtDuMnfHEkkLMuH/rx+kl6V8xgQX8Y1RKojsZ6/rC6PFyTH9h
EKnE50nUjn/wY0r1WUVzU1vdkYFiMYIVW02HtDcwU3IMKNjTy2VUI5IKQjeCJ58QJqwZ0Hc1xw+T
s1sQSDs44cliSRQuxJShXJJoTR0IIJWym/U1lKdePwRfeszhqwy4LbcZ16Uh2kQzT1UZ+Y5u/dA+
ZARcro0VA+8asFY8FAvqOTLIuKFmJrgu0qrZ9FtQ+/LsSOIjcAoJjZF4PlRXP/lsNc6KF+PS7g19
to+8xv/lEOZLJwPX+yiHXe8/cWDpaiutZ3moqMLOy1Bo00kPbuQ12udahkep51RYABjzX6mCtpm9
xwkQYC+KhBttl5gRXzGltYK4MpzDb2JRmcqPFWZVkJam5p3PehGOdYUTpZevYezWQHRWDaQUxUMu
SXXIYxIpgb+QpgorPcHPtst76AbdSEMZ95ks6GbOaKKdNhtlWmxWE3bSc2xLr5nlnggsLv+QXH70
CDb/gZXJF/3qiAFUEb/KL5cN0iU4DaKTbPcyGaAoAyM6dIEgGjA4fZUB1MwOjxD68JtFjnU2r/gn
H9U7AnnDWhTy3Q1A0aMw4uvhSeuxhViWlyMJJVIH9AKm6Su8VemyNSC+JY36TnpE7DkPaotao+Kv
Ip/KdPH7+YXHh4pPfGvGpclGedeB8tnVLe7Dh10RZCEC+QvnPCaxYwbaKS7FP0trWhNg7jdV/ya7
s33D+dXDHRwca5VQ2drKdp7U8oHSlvUwoKVEEeXuQq1gmuf+IDAsVrOC7xvqzmAaLoA59uHRiY+Q
jERZJYq6ZqIfkYWua9swhzs/jnrYtcrn0dFI0ALTRMuDeFraIr1tZdEzacAbvJ2/4HL7kERaaZIa
cCjUFowwLnGADbfdK0ICJgoxV+VAwXeieq5VJ4lYEBbh3Wi1Hcf2PvYXCYc0IRlM4du0DiOyWkGL
roucKkMLpf9YgBkE/qq40n76gmh+w4o7uB8CHwSWsWfsqSNXSiAuUW5ArIBqks/8RjJwfPiYRNhy
mWA5TG611nTCOTKAGx02h/Kl93DEzVrT0qMqCsgi2P5sbMvPHnfhTlDtLDOOXyHzMPwdfZMY+MPc
dHW7S9MizkWPPMRAJAiQPPL+UCDU30elajh3M9TgRaeAM4r8ZCMSYWbwgnqXzQ4Ddao4vHj7le8B
IWEkLi6AKq4a5cYOZAwFFiLDCV2XxkYioPh4cJ9oINd3hw83iixtz57WQYR3mu/2rwRbrHSFQhgf
k3GimKCzfR1LdzAR1M/fNiI7hemz7GnGvNPDZS1FJiHTkREO0nuiZxzdzxvz20d5XI7cBIVkF6/i
FBDYD/jNxgaGZDxP9BDQ0i6xCJ8xYIwFUSw/ERjg+g4DXRvyzSa5E5gxjV82rATzkdp3fN1qISrH
axrGCHFVHqxBK3QsV+umxavcRluZIocXYOLH0pd7EYsYm8eUCkNbmUIY5CyIvYT2rcNTgaLYpzyF
xsNWMzegADMxCX68WayuRjsftByPO0QQRWAdlrz65MJldUVA+nbPKkBAZ/0zTo3zFjMsWnwpscNi
IrGrgkCIuahNGVh7UdMwGes2gW43Tog9l8LtC6unCxunAVn9vhvV7k2iL/2mZdqLIYohKNVywkjW
lUTkHHcb/IO2PgMsrjElgiMZarj9cR1ctlr34N41PyZYrtR8JYcRSFtHkliHr/ot4AiQfgOdmvoK
mXB9PQQ04aes+Q+nEC8bPnmcZ3YxCe+1ICGZ4Falyp+38u6q3US6wzNmRCC2g5CdE4dzZaAHiNbP
K43BxQY/oq8pWD8+Wbv8F1nVLM2hF6SEFiurEee396aXBcoNiE5MI78mAbAQv+Btyn+fjZ6CsnWE
wAjRfue9e4hY/WSjZsxHzBIT7V7dQjgxYAsct18g9+cGMNA8u4PTBEbOSkmDCJH6lwg3BSoTMSqq
EhdWPH6Xmo+/97Ce0gn2c4sSLyFGsa9UGAL2bCx4SlDTlAkU6DWSSpeUtAH0xL7Apbqv1Y315VmH
ePsvVrUibMavdQJzuc7G0F7VDXq/zjxm2V399HPsTLF8M/HOSdlVKWdAQK00hG7eLHE0fRQoRMBd
VZwpj4VZ0KJQjeDsszVOvMeAQL1PAw/N5XEACcrgRWB+j93A2cJYdmghvgsJxiYJcF8NfcecE8bW
iaEzNjOLyvdkx1pB6z6c5VNys+USuDm2J7jxUDhMrcE+EseQ/o9n9a3+IkbGrIuv5YtNGfRiDWM6
V0UHqxq3KGa4DJ9kG4evW9loNQ7q/iggJYUcF5NanAYyllDjlI+M7+IvF+qUXXxDmlCC2B63Y/6e
U84WN8yzOCGDmjMum1wKfhIMzWNb/o7sX2Q1mdYLWW+wCfMKAxCwcisdw+IQRx/9y7VAYEmNx/Tb
S1Ec41yirVieVHNLk0rY5oAYRpKndFX0HebP9zlntL7PSRDs8n0tPCLxLXvOvBnkAx8VtNnDoAPd
lDZ6mmmzg8V6opTC0TbLRifNxpe+uEBG5YCbIU87kg8w19BwoWfPp7kxiRK/O/G6VzFYwHmUprsh
wwevXr0RMd6eYStwoIhyXS5RrXLdFJGM0ofwOu0CeFll9bOYYaFAKgs+qpR3dAKh+xzX8Pc76GqH
3l0ltFh2K9lU95LHXEUYtIRZLU80cgN7K62S5HVFpj3GdCYnWnT6Sgo+cYP2AY4a3gQK3aExf4PQ
2x8aOj7yii6n5KMW1sFOzsG3CvLndW1jjw1z9a+1QtlIa0btlEUCyDvYaKjUwAxT0S6aerc22nDd
j9GZ2GTDh/aMaTZ8ijxx49V3ZbaE87eBmEd+viG+q83C7itxm2fPLestm27q/zBPhggLKTnKfieN
uM96pC7yz5m/G7G/8XCRPEfhf1CViOCMOuPRuPEa1rZJaS/hd5o1Ar9NPqzmgX6dz5IQNbM5craK
kC7maOhxiQABwMl+1iEUoTjNnhIbJmJBfDR9krR3skZozdDl0Aerf0gUW4g4qWVOl5xnfQMDSqEB
1KY2NjiuPwp1n6zyCYXXOQAh9jOBa9eJaywFVmLfJ9BEAKnJDDIUAjuDW6y+h0SqcbgBHSdARfFj
ZfNWndT3duKHCdyGf4mbSTAavyhjAMSbNT9Fr8Gjci5D294/RYvZ1wiuBubk2K1mW+5YQ3rUO7eB
2R3d11U07LgBQf9rJhPc/+dsCPxQlH8TzYb69i6xmR/5xSe7RD97b2WR8noo4w9XokrN7Abt66SX
8y0NflpRGeoQtNMm8VBSpnbXQWQ9BKToWWjzVAPXYje7JjsOaLbQX7Q4vO1oo5X4ZAGBnCydoZKz
pgNyvFoBY0k/AKl6QtD9DfTc4oCRju7ZYcca6KZeeOJSmTKufPMWbf9IY8cILTYTyCtQ8Rl68GPG
GjNhaKZY9AO2OufOK5LisUKTxDwGrDCZ/wwj0HhAjsR5F7q35P9lJxtZp583I7WbzgwcFXNFD8jO
JqhIIfrBYGzjy+gz6AGy9Sxdyl73pfnhTQ8y8CN7fh1JB01nMC2SJL2j/knKfog9hRW3ODorfpO8
DtxBKL6wF5eD90OF0budGrQqVa85QwmRWsA61w9VXfOiS0VgJMY+CMvz0JG6oRqPpxihhajGuqRw
jdtjLeK8TMtv7hlhPCCRmZa9uE4EnZuTVQrRDDdsqHk88T6WZxiKueXkY2WGnqnrg6wvUOnhWLBG
iwBXzq57aLFZnRvmjoRhK8AqG5gnGYTBnBlX+2ZI1PUhw/vUDh40SAZS7RVXWpevQRXdwtW9c6pj
3Z5AyxXNR6lfiCQLlLas8kKgLj9qrP4Cq4RB55edlDPcKvnRme/mEAtCcZMBQF/tj6IMfqfMF+xV
XTbe4UBP8nsCVedf8zr165wD+jQ5tg3oSV1FbkAf9ZujDMKU7Agf8HBgEYmMPQ2R/j/2BFQqEidY
AJgRmaGJY1sZJQjh131J7pP1aNdlMiiF2kv9yNCWyyo0r7wq1eZw3bZCqhp3PX35slcxosQ7DbRi
9/iRhHdbIO9TI7y2BgMw7UG3E6YlSWH7YCnyWYsFEyaoVTPRd/crPgLH4f1e+mY9zeImqc3b+c7G
dnAzLr9SnzRcms0iEKXVo+wyuQOOrGuUJg9NQc5rIptf5llyOdwo/lK8Z2Eddb38QK/ZggAWRe30
+TxSLrT07E/IznETOx6BsOgbIU/tXB9uD/JZABb+CmjaAArptRiFDbcl7o47Z6VDctTYbbdrDhI0
ZBLGmPSS2i2MTIGKqR4Ueaxa8+8aSQyOicETsIf/j3iOjoW4hP9t/4jumGfr6xFFIhSO4I34CTAD
045aTQdLlHLGxqrjaYnya4Y1ejmBIhdMosp3FnhkHPy2PPneo23foaiQuBI28DZLmnw0JcteCGUc
rhr3Fj+6NePlrnVASx+ncwjP1fGZdqV4WR+zymwMUmIxSLAEmXg7XGci3D2sPxN1xzNHtw5pTcNN
ENdOXLAnksms9OtIS8WRXfZYtJICa3fE2SFD1ccmzm46hwTuoYDmmHddkJKA/vpLT0gGTEuK39/L
QUC5evGnMZulEAhOsxFZefS7MLnL13X2VLcNgLmax98cXNycwemtfYI68GiF68NoBIhpVBD6Ek6E
DXSNNW9wwsu9+V56ToYqQpVCC/qs0oBgePE4Vtz4VPUm+P2fyn2ShsQRh7w+ZrSUNi7xwBf6ZNT0
9j+MPxQCwklxO46MdHsS4aiiDafebo9lB/SNdRLsqfu+omNDHfk1IDOhByiz3xsUck+upleraL8X
c/yLJ+HHYf3Y/+E9oKIZE+KrPPKR4uKeth456rY3njWLqw01o47gEmprBbW6WoP9+GBBN2BWI1Mm
sTCFAHrCfOEJ+nK8KQHWFpbOGhUX7w9BXdX1KZn9NylKBjQO3OzkVufD6QGrdCzmofGZBolIDtsz
IayVZimMLSmy/LJRQ0ude5Hj4/PkElOky7dxWgfQm9hgYhqyPQHEOSyDPwFNttqSk0KoKQIJoAHU
8BG2bDhpnVOOQMK1M4lze9pPmhok4AuBgVhBlD77wMRER+1fSCiBYHtkuauwIwuCZ9USpjgFAJAV
DYbanaBXa7Ota0hrj3RmemmAoL+gZuv6Jx9u3oOtCP/7hPI+klVxPxU+5lt/aQv+VxIjQJ0YbwFh
K3DtBWr2EkLG+IN9MnWyJzihRlLBdKFAZXbphuEHWvjSvp+jZUDoH3ufYMQsoQSdzbtH5wyjnVVQ
tMfSJ6E4XIchI3EH8Y0NBOdZirzxOO6uxiSuGi0l+6vQtWySYnYphbYkMkXXbcoO03Tc2jpA8eUo
zYaCn7wKi+dhJBqJGSV+shDF0Rnrj1SBj/+BL9egcLcjqN4P6uFjj0KY94E6+AlvD4tURVWVzszz
Cbgxuw14XfgCQXZwaNpQzQ/pPHdhyNPl8splMVNctkqY4j2GeuaTuxjT+XIlaQDRxU2225g4WEIG
0DSH8KKQg2rlGLPB1GG3pdnGVYjTvDFkujPm+iDFYV5XmA/XH+sDfbJz+lbLb7VEm+pbUkLzKs4c
g+uyHKni0/7fZgpz5f5W8LXckUrIVM60rFDh+bQMXzTZkFCjeAyBQncXg+ZECV3oExQ3mAoohbBE
t/SsleeqwIGmZCJXeTcqVYX5SP6amLCXdUBnYu0lKKH4y2j3vGJ7WOTXf1LmZDc6MBCPeUVg4xln
dDwVaiJ6fl+m9zMFa3K/ED50Vb7TUZwHV4VNss0vcQBDKK27+amL8nOiC7PHWg90cARXctLhsc/I
axpRa0p1/jZ2/ax8F5J/E00bESpKBXk1Ajonn7+TJc9oDt8u5GkkfyKcvC+NKvj3yZ/GpGsvwZh/
KA5C/4lzTNCGasIYbS7aTc5w1jOpfCPnivXDW0k+Ferj+969kkAOC2Aqn2JdYHuT/IN6MvAT2wJ9
w03K4itpIztxlDvgm+q3SnZptiONOkdg4vDlLFSrwCNy5ypXxMjm/Yfa3qTzoYhqbthmegMEXpsk
gxuxSRqa5azozm/x/sLOh9uUyW+ugMOKWzQEYv3byMIDvKewDQrDt50p3hUB+vwgnt8eKflLbBKM
my2mc77cy8xMKWiC4HV8CxBtn5PSg2xa7Cvj8d6B27pAlRNS/aAiMUq2EomwDF5tZtZA8MlvgWMM
qL7sfxH4YphLXwB3Zeth36tfGNbpWUx+RkkzXhd/pJhN3cVCNGYqTw7d5/mcwcM/Hm6LyuNbGF3B
ghyKUQLfgxdCAjU/8wMqyOIH6teRa2gK27g51HnnwP0Pae6Qa29nMpTK/STCtix9M7Itl5z8hxiu
1sOMCAEas2Wi/8WasDLFsY/PrEbv2V9bHPdXbjt3XEplu2lvp2OLiEoTK8kw1icgsQjP5iqWYQxX
ua8hpBknZ1lsXE/aoI4jXN6YpnZHdnyPG+qMmd3NDf9G6l+H2J9NIfr4LMgsAMTHM+u76ibAxGSZ
yrDMr1G6Xk9V0gyGJEU68nNRBMbqen25j3gGeyP7bwvn8Vh2cRZVo7z4NWP6TgQ3qDgXmWLTCyHl
LTIIjYYxoeYJ5gt3IE1r4E8JiSu+dSQ531DnWjMIl/gQB9aVQ4GEQJ8rfV2sMRvEP3v7MeYuSxp+
k9BHyykXke6+0o3Fyyg49PtYfxUW/4kJtIpdRLm0peM+maTr1LkljmJTz4d3S8joP4mOR4XCD8dV
3xszEa51v21RS2vwMGRd4MdRvmb32khPNw1o8Qm5EshUZqibNdbV+8Z34fPEIDCXgry2i8+UXtAy
qkVuWUhnoa+QY4j+r58OS7t5hJHXnEefresmK2ZUKKO4IFeD4Yqw4S4fsnKqxI5YXcwc6yiqmy6D
ne5cns+vN/07ogIorAKGfRvqnTK82sSrqft3ExFov35BmH0DTforWN44tuahCJtjI1r0+UCvm84E
zap4HQ1WLQm7dGB/cQD7vxYyyUJbyvxzwjX4+qA3d2Em1KMvaQbte3sZ/iUuDkGCoiUD+nnn2uzA
o94hahbv4MRATBYSrKF7ZlGOFZzp4t4+EpF0OcCt8K7ZBHMe+n0CKXk4uxnY3N58CEHELIFuIUnF
wUx4SpynjinBaLmlsoCz6gRwhFTmlIcJMD4Uo7+2zpgjtiyKgU/du0Rf+L8lhDyWe7g1dcd1su1H
uP8RS9XdIqfiUzR/06/ovTh1RStrGAArBoOFrBTJJ653tV95BtubGRNaBpW+7BLpGp6vyIPZiloV
LfIuaDTJE7HeJgEjwXxMKlyx6jnzXqgaKp57QQZXy91Vw4k6rWFYqRzJhaozWIo2tSpyhJ8bqeMr
3OdFEXCBAvz7cbGDD3zDNaj/WQIJfW2uoEuTtb3egPNllaKcH/m/sYiPp4TuGms7fHEHoJVVDAge
4l7sqYYWXoBtdqPLrL2xkfR8CJ1DjQ5r/D7wVkpBenkApl+jwv8yxwFE8VlQDASuEezFLKcTZSMy
s4qI6YvX7BUE4lN3GTYv/O3brOl30mcONas7TnzbYdlJQ5a/AogN9Lne7e3ETKqNCG76jbaNmdUk
eTia09PREwmIh3h/nXyqeo4n8q2L3ocxfCZjUp6evmKAjgfGOZsdooPiG+hLMv78N7LbqqwuFJMl
ZZq6+R09pdADt+fFRN4wMmy5J/aficB95Q3G8YAXwY5+/y1WuFNdohOy4sXru6wJw49zq3fUqCC3
N9xzCCvECMTjNlahuO5EdeT0L9EmiajjD9NnLA2Hpjm2wSSqm0P1ZxNKj6UqnWnB7vhy5Obim9U7
PQyv/Brkgyvd52CiEs1Xs78s40ps7CKh+eZRiKSowUe9qUYqpConWFJaJSSz7HIe+1hKUVPfjlbQ
wu1usB5bkfOL40mx1j6664yyiKJqPgqWWNQAwj5ZptBoWXsefIjECgvT0sHIrBSoUKa1ZVb1GLkv
F29BZXhiugg7f8nUGEfhslWr4KIVEUQM4ceVbI0VTJbauXd3hzNi5ESi9ZGIKgEBu0hs69P13c1G
xh5EaGYVio4eauRP4s7Nr51Esn7D7g5O7cCmSecFSl9lOnNkEiRCuI3NRJus/etf8Qdq2WSrGXgY
52sL9OOsIkWhYBactPUQLB0zGXGADajgkFuJvaztuS9xuIDc/A0IfT901fKRJ3FaqJtMS4d7xl/m
5mVZtacxP0MzKu/uTTjtpSkLOgZnT0d9JtFX0jUhml4FyNwBgq+qf/1ax5HPZDZMHBDqDTa1Xbn2
j0oFzb5VoU0W/V289xRJni5Qwh8MsHwiFGzPT+VX7J7RhRNVUd4WKARZjL4JONHs8e372NSRsUqf
xsEbvFchEhSD7iS+Im3tEaaR5xrL7r2bWSfwkcjdoIPlrmjqdJIYI9GElntEbQVja8QEK2bXXkPn
aStNp2eOu7EbPNKFPYU2pdFTK1fd68DwJx6Qq5J4gUMRO/f/YUrXWXds8pV0g7UFsDDUOC9BmD1J
QEQ6HyhKV6WVsJhHIUAqD0jYy0s6w/9SKkD+XQlQtTfKcHdbyl/b46BtC3KYbETJYPL7DiI2BMT5
4wp6yGGlRTuYbHHrdVYOyt06Cux+BOZS4rqBQ5rUwCzy8jheIFPSDqSwsOwDYK+snxws2+kQ8era
EP2YeEsWKkAaGw1t+L0eKz4e9epV5h7CXxqlWVQtInrkg/2lnQp5+vqWGhbB/xX+pyQWSy4LY9kF
U52DyOIZgEFWlOf2c/LDHOcWYFl/LEvPlLKCOw94n/sxsvO7+C46YCmFzd0cfejBH/Grf5g5BDH+
Qt8OWfKHgMNqMhZI8m5TZluYZlfcSH0rpWlCp1JRsZoPCOV+aFLNq1wYDMLb2FaLXhFihKdIuX7X
mjKpN0XhC42RlCv/2C8kY27J3kAD3dx7c/VtdvtwEFrpn1ReA+Jqh2yQcOKZme6BJ5k+3/XJjwOw
wvN8e9tV9CRHQTT29i9+/h1Iro/0gzQ295LU17Gpmn2WQpLoj1biOtQ5KpVdh8HCSwax+BiWcNzy
AgYWAf4YN/AmjajvvlOu2QxGL32ncNKrEryosW+1iyNjMxTFDvQBZDt7zhuUtrpzqjywTi8HDPIb
VI1jTphToL1nLo3prTYQMedyHlbrSyqGWRSGHfGCzW7LQCDJ3bYFI6XtOAi+vplfiQLcvQTgHGuK
/U00q2bU6z+RIfLSa/rWly9+ORY46jkX2HaDj1Sf+U8VXBGth55qU0fjnDCL6kbHeHULcceUeOGn
pMuWc+oQftvm3rW1z/PLq/G66Vm/YisGeyMeGzcWT9cJCV13Xv2Ep1yMjiRXAQ+qzeGQ60Z8haex
3VuU3Qk3SF3BAEIy+8AoKJuQiskYX1LsXttjpDPNAEO9f7XiKJhXZrhhI0/zLzIQ4aSpFV+7scA7
SDn1zigq6Lui2LdwrryUjRdwI+UL4UjYK516ZlDxWZm8LasnrAFs4wx0oH9lFb8Vy6FLYYT0dT5J
AdO9B5G6LyGG0g/b0U/jT90bBIp8QaE9zIlvWbDVj9I/YlVHhdmeark+FHh3MHa3jU4nqbpHzdGj
JSy5dLaLub3uvvvMqdXmMHUdJ3ArI7CxzCkgjf8lU9oatnDsNnqqTotmWCtDo59aaEGWKddBqL9A
qSzUtGvxzX/iP0Ya8CqG893uIIpuvIcm92byo2OuJaatMCYaqKDGVLm0BoldFdxbsUYSSRj4Fnz6
hOwVC4g6j/3ltCgcwZohiZV7SzvQjbjwIciUH/duVfS6ACYkQ9rt7eLxYaGedW99TkSKOxbMi+jj
JomO2OxwRR6+QTKZR/H82fZcqDQ73SvQtUtNmLWFypWMHgNIEIbd4aXxaQTLsjLdj9GsttI6sCyV
mIbyhN8icWmbgP2gi+bytMybTTx7kPBjyuhN24K47UNU5wc1pmGggZZS9+RA+xahZPX8rrzsfXne
yqHRQjSEWmICG6k9b8MrwAFCoSLVb97JmBiOoBFlyDlMeHOkde0+A+cwfeVu0SMQQ49IyNiQZrxZ
sTas1IDo5NvO/lcSHhAY0pkcTsgNZPhyHMUj0AwxKmHJj/F14epigJ/ORQ+fgOr2TYsrAgqxJcdz
+RP1F2V3WaqKysdetbyT74XER9HPa7XhbPxTDfWKl36+x1ac3hFSYuzlHC0mubr4ku5OVo9JnSOJ
53tCp20hcn+M2y7svn7VpB97KkXvEzwC+dzqX1LMweuPs3A0ucW9MOHIKWvXcWLIlQcfUOdSYP4X
IFBhhL1PFoVRm9LfYH8iR8ksiZ/ajS934WzGkkh24hmPBLlrlgNGyuwGhDPmu+Ovzl12B1wKNcPP
B9WtUK8phk7/ThAPsNQGNBd45+sz+y9nM1FOfurBCuM0ZqZA+S7A6Ak6jxRTOtMMnC0wvS4RtXN1
4kCYL+PEaKWx+F4GfeTA1hhMpdmlACh6G6mlfZbIsq+DgYLDEDlNq7bKuJxRqzqAOxA6WvxnqcqX
K33PF/NE/9047MXvVoAjqQUMTJ1lezG2qKQH9cS2XJqS1X5VPCEAU7lI8KjYhysnrllODBqrKITj
01tZ64AJrBQzwrH38Q5P6vEcaYG/7NZqp3RfbT45hxUPXWkCH71FxKmYiKNBQ2h1igC93LJi3F8W
0c5Wz5vlPbrFrnU27cwiHHddTJSL4+KEnJpsn0qU5JVV2YfQKLdFXWh23nCVJPVbYiPKoHFrN/D/
7agYo/1rISU12e5ikrLoQy5qVftXlnYmy04Qti8lc/7iX0q9aZ2zTPoA4f4jv5vYFDBk+glk4W7G
rEwKjEYYWWngURJQgHijgxx5kBtzR6147uvxA6KsN165DnkQ/KA7YfcEAKFcqiudiHUICPqN4LgJ
wv/NRxA29Z51+sprrsEhaifT6ye8e3K+JMSbFOcW2HGXa0bQvawWBFOfr0JwA9pMUQaXBmQf87p2
6r4PVJCsnPEmqw0yHTLxfEvZbtIYafP4M7Sch6oIKyY1gidCzQa+m3j8Mtcio7KvTldr5fI9BT5W
GPBsA61Kq36Z5RkjOLy6N4J40hoc6ZYNW3t5ZEE3JylRtmFYq0+1c0YUPSTqyL0uTmrdq767iv2R
xXugE17zuNy/uf1fjZTYh6EFk1ngTC5Z+9xWNltwTAo8zyI1tH7DuVi4lnru0rfQo4VbClpifT2w
RmmXrAC+eM5A3vYn5Rmo+X/zNjCItdbMqeioe7EvDtMRzJ4kQEmPsch4mbE3A1rac0vYHvUI49Me
fNn3ClsWZjWcRIotaPeQQ4mmV7ZPum48R3SMr9/SrorAqK+Ckq7h4fsGX2eQxL/9Sp18fdd2aoWa
arqx6W9rMZxTLKB8vxC6OgyJri3QBL7gseghqUX3IIBUMgfrBzs9ZsTF26MWriXVerL8riCGNUyh
jyEfm9r3pIJqmJfHRS+ipv4jx2QFjjri7q3VlzylXk89MIMQAaD2oH8U+sQVLpNvyE97NOwWDBXC
cixrsO6KuHPNiCAgPvHrUdZYRkTc+EPIKOGvMppkj7ARfE9R4y+Sflv22drVt/nqheMSNX0YzgAE
7VkLEvwPL6+O1u8wmc6ZPX1fxOe5G7GawrjrvZILqFNmCiVSHJ3Vw2o/9wUhp60ZypIIWyjVuaSd
IeZLKk7s+eyWNe+WqFUx2vaTbJWXnn/Pt5xIxQ4pD9Bj8mJKT7r7xPjDp+5o+xeYe2ZwSnrmuEzP
hoJLQEIYKEyDWS026CHsx/Wq4AP+ClaiOfTkDjJCXli42/M1mepGRxgRhVyC27nhSKYkM0tOnsFL
C7af0NRos63hsKRnT/nlexOkoUfAqu2xz9N12ejxCsynjXl6dZP3zbNFIQs9mjicKbHDdF0OJ/zG
s0+r6XKT0oadoklAf8jfrHQqrtP3vFa/GywKEdpWnrPu+8ivuEFWKLvXCGosGUwDQPPRsGgWSEcj
l5qnpHATuQHrmefQFWzLS1EXkd4sUHADCp2zOMJAgY+B02vqs8QQC5Fghk6x67sHc99ySKSxCW3n
H5J3fRvbReESQ7AZdM+ZdFNsyJubIfk1bPUrOH8oxxVD1Y2HcBZ8owf9ULKK38TsQn3SN5uDkh56
eDW2FjYMPCQWSkgcilw5TFQHZD5Fk1Fsi33mgTWzuCNxjsC2/pT7LPkH7bqOUPZeoxlTZ2WJMkoI
AW9NlU7m+TxoEi6D8R67Z5SOSB23TguhrxYCQdo2NzXOCR8c81lJ8q2ny33x91NFk6zIe70v4AtJ
GZaS43rJpE9uqDBBeV1OInEUN6HrKrho2c8bNQp3ThfBun+6vjsBtyHnjY80r/lxkma+2aM3+9Qn
jb8Sza/k6HN0/oRZjWcueEo+0iEWAII4VYd4NmKgR6wojgsqEevpa/47ppQ2IyS3JYXrZbYzs5Cm
wxMaulvwOmNXb/wVuGfrVHzEz9G0Z0JKjeQ52+uPc2cgTT7zNHyYtkT2OkUQLw7g9sLIozkCwkVW
yuW6wzGVM4c4HvcLULwYpEOBgcEpQ23n/AOSRUcFCcKfJveKZPRLxF0xE+wIRioTvXmEXoRTBv1j
Rrm7AxfDTHctteNnMtRl1AtojiulIU1LP/ZgTTRER21jJ/R3gpSA7kt+zPlD3iemgYKxLOCPWMO+
hrv5VJhC7pXqM7I7Hovhp8VUlfFd/loVjRdSDBuXYaxlEW+xwhkynyra9LKEzLpMB3ib+3pmGJ3C
jvbexFBBlDGlOmLgrSejUQ73XkKs3UzaLN25Opp+aACO8c4DeCaMzlbFatkmNvQmFvQA3mWwJXoc
k0i3XaN8BJ51vOwoDfsj+42e/DzG6CEUyZ6fzzELpdK0UsIW40bK+9MdUD8eltW/YPFaFEr1FGrX
7ByfVjFK75y4pi2fai+C+TV3J0xEPfFpaX7NwjNYPItOvuLYTX2PyiBd6UCMxkjxoVCkbjQFkAsU
T4IIXH32FIQLU7SH5Hry7tme2WPS1FbtMHqkj8u2yNmKYl/3IhGvNI99mdTtQSIdBz6i/GVRWXSi
3jAFRUZHnyrMfXd152fm0FWjWF6pnG6dRhp64m0EhgARhfhTvx2//dTT4kfJi7qF3n/6G2KqrgSR
Lmeu9B2xwHNGiwHgzn7PlaLoHczPZKEmVi2EY+OMdusFDewzlSDHrhERId8RPJoRx743STrUQ67x
VWDfI7A9HsTEeQCFH1pTGSthrDPx1rHfTMKiwU2pjBJZNzcEE0iYajvFbbEcxieUSV/o2o3xuSLc
YgqiY0GN+aBUhB0Nriip2zjQRED5cKBcahb31qFIb0mtD0onebVkxRehc14mc1J3POY98i9ltLZX
FsQsV1Y2LVo/RLzHs/PuDf7fDCAxPe97nHge59sE8iQ8xoEuBFR16tBdhkRgFlAr6bs9xz4k0tda
X3iFEFKI0JZZT7yEDHskefXQ232AUnbLJSg97z1AOTjaO8s97SoYgv6WNxDyInPnEQ9I5wCCBaXN
lXpdJ8mwO+APSmx9hWGooBVb2BWaaWqy3dbosFaUUYn+W1VJHgrOsFHZ5Os/AjLDrauFF4xQxRcW
4tJE/tgf2nFQIsXRYaTPUXYRvJbg7KUyyXAcY2Tr+e3F9OKgqr0KQl1jaSoqwddgOhOqhcXLXWTQ
OIQIvOSdP8BHtjaDOeUEzsVsdM99hgHNPOfj18B+QRH9NaE3LTZ8+I5DXJ3Bnvm81SQ8Fe9R2tWJ
Uyx4+5USKdLEBt3peoHOmvhURcfxPP1+qxvGAh6euxfq5HeSp2gYsnyF4crHy6U/PdwQAsZAzvFo
d0c6eO/cIcT26U960iJBrCY4uAqdLzptFd6TCx7EDoT9fX+Alhz1xwbuoWIhVsvJEZdbkFSvEu/9
gMAqBAD9aTi+Mztfy3Q9UQVQJoh1ajM39SVmYYNF3M7BUGPvnxMODFyE+yuzw/m5BFNfzud8iXBF
+10QyH4WFONE7r51JFfPTMOlYiGJa1aWMdvUM9B/jszRJdk43Nysd4Qxhqsn+E0SUmDkJkOW61oF
7d/YERtm1MNV+rpO6JuILIrLAGRDQPMjbpdDPc3m5mFR8CjWKwl3qT0W45qdK+xIn9WBh1umwgNC
T2FFsekD0PdJ4FUXSB4NQFXL9DrdwXSz6fcMuwGtya/cs2+5EoFOpaMDRr8aQkOhjSFhVApjdZsl
V3pxaxms+TNO5VxNRmPUhTYti0xpowPSfunemezRbv1LZBFTxsaQorykmyNa46ne1Kj1vyJHaGbC
c9Zrxqt3XrGbPpb+/wt2wFMYSnM1b+4eAv5TlFPvcycibxizZ5sbPUCAY8KF/N6KMh5DgNT4ET51
xb/eLCDeEnRArFRMK5iA38pJVUnoYLCgOIgqyG0PLKmcmusPaI8qqRYayCywbfHD7e+X8h5c5krg
ikX6n8cUcgqTvH6As6X8R4X2w8gHgT3TUpcRUcYlPLF241ZBrLyXbdYtKczKiPHGRbCblgNiaEaz
neV+lizGmIF0mdXj2T/ib8VTLSFhPoEulSNOzSJo9/kfr7n2+ljfC/wK6NCRX7wKrXjk/na8tP5Q
Jl+mBv9zqs/kl8Xd7GjyFKAv8ZTGrZlIzC4uzK9Uoj7YFRdWL0kFKKJOJI8WfPQ9FODrRuxtTx8B
P5oplkLbic8nn2rJebcBKqNC0AxukB22Rhd8R4924S+1lGKbOgYixMAM9vqoheTkX6R9G4T6CXja
TsqMviKmxU55x9IEb/xilzoVvHxytz4C2Are2H8wh1L/vpOPNwcWxOp0uqrM+SJDkvfU7YKb08qx
79mNzx5BYCGxpJ0GzlrbmDHgOTEDGZ2+f+XU1DVuWy9pbdhftAqXvB8j4nkM8AkgypA8cBvb/JWv
BrTe2Jn3PYVRXkpg5phQOaXjnc85EdAVJP+RF/IEqONdRFl+8OPQm8qvA4VpoUXTHKLKFjLNK483
0MT09I13PUq2qzFAYCz6K65zuD0175zmIdmIWpHOnwLVoznmLNL9DyDJcZ7O2h+yL8SjxlA9JK9S
dzHREOeoy/nnUcPkvb7v6Uav486irqSLe/WXckvPcd57w5UNIsZwlDQPXuSa7iR7r5H74WQhOEiX
evi8yBUIzhMiXjFTnS9TfOy9jWiHR2+OMSLSW9T+wkrzBpxHVWuUZ1WfbGidNu1HrA9dTOlmxUf2
f6e4IAvta/Wt7+dFMt31RrlxEIpTaLt+JFFK4a1Tp+7K/EGOVAJ1J1BG88PZ1NuUe873AbVfz6Av
Rp+slGIpAFvPyInEIZY8e5NSo0HbZnkSrUVehfzSPiZodfsstXrxLSYkc9ZttnVIcgh9wAEAdNTl
DkruO4ysc0IObnZos7rGm4VfXh+sY2inya7Ib4Q9aXaVxNHqtT9xm9XdLRmRyu+aenhnXKjWrCRW
n+UTdBRlmTjXSJmR1T0dsFUZRNiuMMT0kliYojHVL3dTsvTX4cjHB+2My+Jz+BFcUliP9OD6QQn7
3oWMaoGXZqENN+IqnvtRl7FEu/yL6QEanJt5yI/wT4q/V3aoEZN0a2HlFhY24qfhXbbuC+PO0pKG
CtDz0NST3Rt4hoOjlY61cGMTnVPI9zoOHnZl3LCDv7dWXLn7gtTcH4it2NZOW563NHJm/0H3Zh53
YBst9LVAdL0RwOWlHqgZxzJVYEBJf+1uCYLC8ZYaHmllRT97VV0UBzFL8IsmVAjyY7v97OyO6+9Q
6pf5obXMADF6r7uXKSTP6Vf49ddPDrjNI2Z9XAp56R9tUWjK7xfXazSUdJ6uKfJj8Npisrj+QWuB
Vd39uXImqRQNbMklylx1mewcVGZEIj6Fv6lR8lnPAU+31eVdP92FzTy1PDWRzrt5iPfvQCOXri5U
hRTRWy6dRzVJDxktNHrYp2d+7kQ40EH+MPenx8oMnZH+ZrIdtugJBNFxdHPTtoVaXrtl/axA43C1
jhtpzT/iCBENQ524piOSyXRxPo3L9DKH9pXKU6XJ3q2BOILzHW5/ZBD1NaeJaIzAN8G37PUQS172
HrflQHQrBdKElGyfbUS6uX3wsuor0qeCrY9vYBVT/gb4aZRXjh4h7I/omR5xLI2ns99ZVG22gGZW
/tuMXSn1q4Ku5JGGnoFglCuQssmGdit5Vp1hjujFDZauOQWcaX7sMi6xMw+8EJi1ZVeHxw8df2sh
jcxyqu5SUDqvT83IK0j80y3kGowMYket8bNs+W9VrITnNihMSDfdYE4hmXdvq+yIZNnfj+Fy7jib
p0hRwYzaY9MgLG1O80Vn4E9q8VEAmIMwI9yZgjzafD3+gdXnZtVFNoDaugldxdQGaqnY1C/whXnV
Da/VTVA8+DroywOfKfsfYPIlcbHceGGoM+Kcb5Zw8m6GIXF5FIlOoG/Roxsudpd1Xdl/yqAdxUuJ
JEA5EbR3rtTgpnZyNYz73iLZgb8DAslWqvrG51BtEibCsyP3W4nJYrK2o+/Q5CQPNy6rTZn09G0m
nIdUXkNYlcNRpTiMYngo7ms+olH08cN4hwXc96bxkH/exh7YVXKrNHu6YvMP+b9AGhBl83f9BPkb
ReXP7LeyitA8lCvyFATp2bvOLFKeB8zWMnUqPVKFGLljh77p7mgsix4+BJNUk2/rAgkXRXt2TVHr
yVTuN/g6iNOooxxl+jJGrZzyP+LCBFjhgPbnbNkoB4KMUROuGghMt+gKYJSRbhJbyRqRKQTRYZaB
YgBs7PcTk7un2YtjvPTy7C6RJYU8R9W5jinh40agz2tnNEPK3mOCTB9yKes9lFykGry095moCIXy
rIa5RXTkGbtT2g18ClAfIr+Vrj5MCpxirR4kQDG1PC5tS52bf8ZFLD91S0hvGpgs1sO8+C7tNOpN
Dzr8ts9sNcijfKo14+e4ur83gF6uel5ICIjsn1L+rCJwAXRB8X7mymsFSx65HxKMzjJ/zpVRNZCY
+bbLM8URhUwlySFgixSS5KFUn3GeaxfMK45sUBW40KjbUHi49+BevGeEOmiTs3U+NW/GDq8eJmp7
gSAl6CK/fdnCJwA1rYe+/NeoXtPDygvilTBTt5bTQvmQLAqLGlTTRd8wrrW6n3d0ddvtZNo4oK4G
+WWTRbY8CKIJKYshXVbNniHk3MxOrzEz0SzH/OcDp1n28It06qikvfNuTsz2jVIOfasMafPmpzfP
xWs5QdOWCtk0fLnN4f5aRUdV+tCTR6OjMG/Ms0HtsZaJcUBZdJ3FLT0/NlZ+x5pPhF3/NNx/ZP7j
pwfGRzgOXNLDQf7sc38zO5Q4qCGuZL5KKYrdR4eU8cn2ByzsGtzaJ7n3nxjjVe8DvoBkMvqUwZWT
rh1jqxIK/ejCnL+hu4YgzcP7uGSHuVk6HqgChEbC3Wr479/tUTGWeUW6eneS1lwBsfcMvCikyDi2
MJfWlpKAZI0nF3R6ZGzJCVkMAGgwg9d5QOf23A1fQZ3oMrbhGKqr85ZoTHApfAeSrFmzXFYqhjVg
IHtihyysr23IyZFnFui0ZN3jeWFqbjJWuko9YMiEc1dCYWeNGpXHSgh7FITt3j+ZmUvMrzJIeVBB
uEfYt5tr8qeN5qNVdsNJAGIS3ctQOPB+AiGJ4EV9I7pGgIv5U1xLMeZSAiVv6Fw0D6uh43TLd3DH
uxzfkpTbCcI3q5E648FABsmpA934PTW9mm6vtVqnNYxvU/l0OKbI4UBqMuYmuOO4yCstWqXBW7AB
p2IvouuzwnbTgxu6ppLIxDTcJo2smYu+d0q6NjS8EVPR+mxzTSkeOnrEChnYxNc3T2sRaM4JcLW0
ucYfMnW1t+N2hPuzMxJT+DyobmxqfQzPwbjFP4xrPUcwCP8fHO7RABIhLXN17HikeYPvWHZO8hQD
d386pQZzQ7KGWckZSLaszz+iwl+xXTgPwU2G/SygHAcydcXrIOhUaEcuNujfyclfoTHmK/UfyH9j
/cJm5JfMxFyXaOG3ihzpppwb3ZcZE9Svsh3NVCWrwaoAGq0frpc9Rxs0aI241izCj0oCP7KW9Dkw
ceCrtEYKK86xDU3vnV5CAL35fBG3whpcem9y7mC3pm9ILfRp+8DPE3mhIwwKzmQp1PYyF9W+KOjy
w95yjnWOm9yDsioURdCOivtzFz+P46kX4rxDjhm7KtCrWaTzIblj4D7opOFYf1ef5oL8EfJztHu+
oBXhDyxf5zIXy9ncLiXVwuqmpEUjNHU/tvUywLL4Z0MFKT0QU5p8JF/xU/whGo0no4cowxCyNE+T
CWyeJSVm/qx+TB92ofM1aZ/5rvY+aum86ZSDSSrCV2AqsyL6NNBTXPHIIMSGSL4wMiU2FSpV2OR2
3fc775FCaG+sd758kXoI8FF5xZCn6WTykbWzkxe8HhCWl9lljAhi30t8UT4KA8kNH+Z5SDr224n5
DoOO2A0Zam6F7AedM2x4bSeowg3EVrQKlIgLXP+16SQvrukfZFuj2dWQQu2puQihq1jUBxBRH4ql
JI1VyqSSWfrwc1VbLpSnNMrac27hLl5OTmxxKzFFIBo64A9dSX9aiY9Do7+qjlMjI2+Wxdh7wdlp
wKj6Ils+7UoI6sl/0ROpwlE7ScOUy6H2M4pduu9YalNbpK0nJA+rIHG8TW23tKHm3h/vH7wA/Wh4
vFFRKF1p8qb6+bFtYmpn3farKRlwXe8a4dGb+0/bOm2FGz216pXrU1qDW/2wLJqy68VJETwuSXPf
2WQaryI+HvOeB7ZgJ5UMvZyJ61Q3OlGLmZ5wtW1Ip3duYC6JzysB2zaT50gND5u4WeHJEH6+eJr2
V4GhKawB+d91nBHgQ/G4LYnV59qT8A/LJwtTVDHcQ1KGedFPIxeH4cgkSMqmy1KhIveFPkIoNz6A
EENAJa8OEP9Y3V1v/wlbIhh8oGlz3hgWPKVLeh3lZQR4ifS39vrxsZXjhrulo+lfIqknaxjm79kt
DXGPiBE/XNnEp/NWQJJTAFY/zt2aCrfFCrY4i2zgvv8+S57q/HN7luPGIuZ1+1rStrztQ6BW/rN9
H3/D0+LEpT/lwgz+Qg74RhDJHCbhVmRWhsHxYGTNjUYwazUqDnCEYMSFDnK4G0w5aTR1y0qzZjkR
auZtvdHjN2NXaTEZvcZCFIYgYwY673dzpPR6YYgqGFpSR1Wp/HL9zNEOfYFYlF336W79xMwa1Zfd
O1ty0KBcR2oXH9hEvusN5TCv8F+go0DFbwXq8C/2MUfWTi0drVsg5OdtBVHYEVTMbJnYLyhpuCIu
bd4Y65YNe3ZZGg2PJcWeAjNOi02rfM3/hE7XU5CwDZVuvBlz6nQ2Y8k4sQPzvqzCZv6bno67HEgu
QMsBuAFjImt4dRtZ6H8BR84DoFzfU6NXseTmyOKynH8DojXCibhy01gPQknBNAPKBvo8tJWB8s/3
D8OTA7LeuKyEotfQtZC2+xtIf19Nx99h950iD9TgncDyFdSkhaumm2rhiRBDM6dbJfFK/uxnWq0f
4gmZNsWKIHTXSY5QN34rON/GzI1PIC1AILo2g9VTg6i6EbYW5f1hBUKwVdmAyYTSs4rJ9DT8g/6P
ZQhkkTRv3G8P5BRmxDr0fxW0XS948zBtBkkraaH/X+8a+3v6zzm8j/PN0Dl3/ln2UarUqXigQhPC
wKn2LrQgnmWJenixe6F0zCH/8sFM/v30M1flp4LBnh6eirk4vUpLAdxAFUJw+jRc+hGJ68XtoK2O
B3KenV6RJMU5Z0lQZfpCLocZS4/aXbWf+PgVCNCcH5LmUkxZwFPe6a3gEysHQ2GK1CD0dZWi/ue2
adfnQjWsyF/m+CSRo6wVMv16LEh7RWzb53GoPt28udDXleg26p3BbH9SOqF6FH4oypTYl01bO8EB
s11NKYKjJsqn/1IEYlYDILLDBU7CPzA3LnkyTYANHAlfhNjLwmLLgKkehvYyHj1h8FxdtOZmdYfu
OeFSOQ4uNTVtPgq9AKRV6/oScZg5BMWnCfA9sLi1jJHNh5OdPx7YLiXmvS5l4tr4rCPpJO7ZXrR5
8NbIQOjAKeMIcscYLmVnJjYurf7bu/gDdssbfzuUq0mayWe8V9tYT68Y23mHrfWvLc2mHDxYtJKZ
cksdNRG9nKIfJtO39jxHxSxuUiRnAIsVoC8WS2wWMrFTZsjTD3Yp0lAtQZ0jw88qcZviJn5eySAL
Y/0d+3db92ed8gN9r3ikNFoocoGB95vVC9V725HjDxpXeqrgRNHAC3c/zU6rLUWogqsGB7lZTorn
Rx8hhwx78PHpEqI4g9BYNsN6wVcd7sTCli+dLaENzquqMNipq8xkab6TabcuQM9wbNWfWpRz7bcc
EfbbeUuA+feplFH1rj4F5zZ3HXFTQIqO+S1r+75DKhFHQA+SlIhmo5NHY1V2ykmKivnkZp4db3HD
LyaMGeIQ0ibCIOA+J2OF6wQemE4BenyS1+etdwBfRlTkRyOfrVcHKVQ5/8xrQ2U37Vne2K3TeiVw
FzDrz+XdwuDdEF5qVnRUctbo1lQqrIPPhQvPlavEsZvUPKZ4Uue6jfEan5KVV/Y8nZG5rjM/M3tM
6X/fp2dEyJ231CnFdexqI4X+P6PmHWYycoPR1GCGE7zdvqD5xN+ooMyVR6leWfYHgGj/rULpKWsD
SqpoxsLFK4OcjEP8akecm271W6UIs0RaLWNaUMv0KPgWFDkdIYa6PECaXpgZ7P6LMYQyrZsuR4i+
6UgfZ/Yk62Qxae6PADNeAq7yUucbjKBGTcwQDUeB5VVaaDgQdF499QPunp3lpTQ9q7sqvXaoBXyf
OFv5llpEbWQ1LWzJaH/UhoYNte87+ycPze+Vq7P6jeg14GrpA8V1+Ok0XkiRW9NUJO7WwDkGeN+C
zwDN7DILnKWLaPM2VdVJFSnDCSFzLaYcEuMsSbjVwm5vFw4pjosCUQ/3ALazNq13aKNPKsgDjb2o
GZnxWzaqaInORtc/7jJx/QLg7BpI8liUzvbk8jjIsWYw9g82/jIGya6gTE4jWmaaaUrladZgfMit
ZALBkGTeRvvZ3Spf8zhlLqhGG7WiBWYYtQ7+Jb9aoEE1SevOP9PnM3r7fk+CtYGtQXJU23hGEwlg
0P893a8VjpJsaWqJZzwuUaEVscbdHKwrFE1Y7XxfYsodsjmwu3FU2NRnIOi0cw0l0RqHVxcUb4/k
Wi2QNeDKT2LUuz0yq5yiID8nT9jBxE8Uqk48fRfnxPUwL9xnkhNYsQok2oXNjolU5YFAh5HSdZuH
1+18Wn+XmVAHmi8X4vCzX0s0jWxzEQUNqvRBdp7FOPKxvNmivoj/X0KwZG4ioHWG9axFUhbHPH+R
5qr8IE8WXr9dKyAKFGM5MoZHayYs8eoM8afYUIHeSmHHeupnEAXYLjM6iwL+KULHNdbNR51DVnWK
HtYMcsPhtqfRCnMmtKYEL8dkttJTivzReL/+Sfb36XHyfkIDL7z05vkGrzpKFOuVd+vsHm18Rgq6
a0SUW07cyl+8no90Rcltp6CScF4ukvjEdN1ZeR4M29b+Xs47hgITWefbG3zLN4O2cXGWerkjsYJV
RSa4RDSdX5y9l3hM4gZ4xznHhUEBCq0XsegYKXOLAGmxHwApwm4yapL6ia9KGaiXN+PpxHdcCLRt
8e/Pa+A2md/d3c+WE59M0bdkahrS3Q6AIRAGVi51lq/VUyMmBz0cFiKpkIsfV4/fanQhyriJ9aw4
GNMAp+fikbC1P7c48qBMQicjCWFqbwiqcViX/2nxknDTccb4fKdrAoLrHFjrDJXH9IBaowYwqnWe
uj62K9w8V+9H4LJw2XBvpdYOLg83fNjkjC7ewpxoA0SUNxD6A9ldrOl9BrJG6jwxwendyr0BLsPk
kO78MrYmcr1pJ1O6lnTiyCc55MO1O46pksC0jRD7uiVEvxcAVGpMZ00F6cyyk08QyPhTH8txLscd
n749g1Qxligup51s6Q0uCV9CWJEE9NxQ8K/z0EKOyopjkkiITGeSAJ+t7T9zNEoXGs56Mt1iLfoa
2KzMywEcS1LIFE99WhTN3+7avqou1VTYHE5xN59Od/IEwBJaWALW1YfMWodOPiQOwS52jyyybEHC
kbv3UlZ9MX2LVXP1vmbaWRxvG35sGUp1T1XFrbZvNdLHiZN9lmpbJhlHIc2TZ3aByBdtsnbs7n7m
kjgQqL+t2djO9CUDckLm3RLw/GZEe4WmrR/oKjcOvcER00vFI+tLw12Qbu32tnqPAY8Zg+Fvi70+
0v5KutI1+31DLIMtj0uljv3Q3DV1V4Gg2LK+2gql3uLMuriNdoi6PVNMVpC07PhzfVNwAklflcz4
NuWID/HAeKVlXnfep3qcmvp4SCFQGML/vDQDEl4YKZ/n4DJJIem3wwZArA+Ti4OMrUIPVL9S22az
rzAI8VvrKIE4dMtFFZB2gu00Cn9r4smaPZt3m9e5Y8kpZjYUYxar+c80S61fXXrYzNmbUb9IgU4U
KAYLyIbFU/978VH/F4/E0hztWmNwkPoXEM51EZAAI9LnXPOYmGuNnFijSrLVXJHBoe9nqGQOrjx9
NKh2g/BRlufAPBOZkx3ALz1YGKLghTZdusPrSxjMQ2HfP9k6l/eKWpjfZZsHmlk9wnM/g5197Vgh
OeNjqyj/7+lCumFPxoli0MSDibvzjov2SriNZEgHh5QnBHBMjZmIOj4psWTkLZPKKkxfrokYLYDd
7Lt95Aq5k2ZfqY9nz38nrMi2qx4V+U0mLOuFOolPzB83M0P//D8nAHJV85xYUdCv4Z2OlkrDz7Rw
yIs25d8be2XI+RDzU8OI5rAx8sld1q6NiW8CtH/rWz8EE90rh8dOsGXBqvLa/PoTRtY72UoALSQ4
K1IUP5K6tk74LkUuCjMVsbyJgEnEnUMhZhgLr7wMCVcgwwWerikQp6ypPKo0o1YGV0DP4HGRYJhu
8xe6krAkxIHFWH8GSokgdm4YVPy0drUmKfkrc6g2Q2rijLP0WTKXu72smy4kC4bnVwMiQjm/RTgl
D09H1LFBsrz2+12WStOlLn+PCRHYF1mXf0VjNBDSrR8/q/fYoto9T7X09Sk7qy1RCyVQwTLupeOy
7dx/VPXbRrc9f8jiu2bmpPVH4KcPZvp/rhf9Fht3HBCTxGNoMGFHQnmQHFOg/cS3eNTr6VbyGHvT
pRrzlVVKjn7ksmmMSeRxbynEFzKct+2pkvjskb1s0hLRRC3N3MojNqaPgKmQHfdSBlvYvof8N6Ln
L9eJg4+F4Yoci+g91rxUsuJ30wxgwLZ0Hd+xZ3o9zwYv/wm0bA8g42RzmOZrzCO8FLEnKswL4dMn
eG2q22VmID/6tMbPc1hWS/im9gvhtBREs03lfcIQOpLO/wVD0mEOZV8KAOY2ZZ3DRmdzHtzoCNii
jXaOOu/lBo1lA2ujVd4AyPlhPFS7pQZMVeLx7y/oXy3JS+WiKX/RQJGy7dJCk2Y9yffmmbBXrf2t
WGvW7YjMiUxwIvocllB/pHrj3Vn8B5tGO3FoZNlmdz3/xG6tapzNklJjx6ig4jOsa7JOJhKwsAXm
0mBhBKRFvE1Oyw77nMhI4u4OV2BDIK1exz/HP8qGvR/q8KKlhB5FQyqi9FY2xpa4vlUQ/t7tx891
A+tvxkz0HaJlWAEwm7QwLZT10MGPr5VLjY7Kzpu50yO+tlch/7Dd6un3eVsmrSpUnPIJAUsygwzH
ecV1VWrC8HGcdp6AHEcGrwWvNE3H+RMek3pkIERQt9pKcl2ttjefZrw3shCBB2Fef357ZQQ3jz0S
C5uobTpKsEYg8IYIgDevVxrPbOaPHv4j7w1mdb3IAAM7zlWUjYj2/pYpPqKS9ylz/VvW6GTralvQ
9bDK4tI/vUT/JYduu1D6rskDeK63b4r/ojLsJgdclgQP/RMRxRZHHkusC0rntt2SC92yz4ENhwJo
ANhBO2oNfYCApfjcgcfxO/dVejKieCfxUIDtp3++i6bGwJ4ttd9HTe8qtaYxvjzww7+5ZVYUKGcH
Z9zOrMAwA0CvAzx3k6jFkwuWKVyzh99w2kDjri2bKVX2RlHmJG86z0afKdrmddOlpNXook/NR0mb
RNxs/G1VWlzG/w/ezdOMD2WDbhAVEweLwrUuPhEhlD65cS6l7FcRSoY0JrJ47CPjNbt+0SuCh+FJ
ZVIqrJkuwsPJNdmExIZugiDGl5HxVxmiS4XIMf1Y3CQ7FtUcd2mOvq1WVBnM+MFBFjcET6yAl0P6
9T5kFYvaJpvVysp7mGmWLueTM7MT84KBSBZEnJef1sKIBsO6QOoYdWId5gt3iFoLoNdwQdt60TRu
xjHBcodPhzfea2WqBaGEtCg4siUzRtZaDV5a99dMjKhHQnzW2dn8HiY8pZL9wlaIPHNQW2cDPaf5
d8ErlBywsn95uPLAaiQ8Ulo9E4cpYVWBQXrsQmcwrWk136jIQVp6OcEAxzBB57prAjGMTrlJTD9C
swNccIDcByL2ILMc5fxkcMhW/7aaJVDZ6mro+Des8sd5vIWw9Pc4bTXe8V+eZM+APqIfJ4nVC7Rp
5l0+4mVJ30YU6hnGpyKGWeInG8sYrIhNy1qr2GuoNNUOlFIn3+U50cicynDyZhIv6UAJ8O93GR9W
yVPRvQxLb1kQGNs/KOJh1reaNCd+vjB3bZljO/+uOuGk+G+9PTBcRXtYVkzX4KCye/cNVwY47zYf
10W6HNL9nP8dwTmpGEmtKQwgvqV3XOnajgiLV7qbvTKm+ykE+KDfJZhXeglM+xcQV9by5vAJ19uc
3a/NbnhCwDObVdwgtXyTf1s0wYp3jiATxUUtT57as2Uf+RUOXQ6DfCeEpTLiTdOwzdgaVytNifUd
smJanrheqD+oaY8X32izsEtnm1e1gNW7UfHrIbrr9Wa9++BkqXlC/Xlm52J2H6C4HmTZa10g1MG9
28ToKJR7LvroNUMFkczSCgcI/i27KSs/RwHvZRDZLj8gDMYpoSLk8Xzoi4x83f0goggCFyAooHjA
8r7/zGESaFPhOVbyBS5RnYsvyLuyVdVt/QJt7Pdq7OLA4yETJYyTxTpIPx2DORh7iPiX73VlGw9y
+8tKuzyqmLL8z6ilGsfi9wLyh45wclqi5b02gJdjKwRGUnax/1jqBwn4Ew5wtk2AQ6xk6jW78taD
HHh79moRtjG3envU31OgSh25dOFi1fvQqRou519yR5NiVlJo8oPgmL4BkYJDOV/69UyUpY36TnW8
I9xxLfhcM5phzPKn9zgjh146vVQTdwVuxA/NWD6336vkjuK8XYgLThUktpZBM6eDpWEUEUmXF9Hy
op+A3uQiqmkd5BwT4ynGa4QjMICKiweBlrnbKrSEHbSrTaR2dmKfKMCse7p1poqkUi3x28MRfN6z
LvedSA0JSqjWGc1f+Jy4XMX/neS3MiT0wxnbV7AVREGO4q82EnyOpChxF5NkXlMEmxmKsQFVR1LQ
ABB0NuCcxcQmc1nUhEH/jAlapwvHu5iSpgStG0NRebcHuAV7MJ1W49CyhKMdyxEOM3e/6tw/bmqH
kAnM+eBw/e8AQ2lq3hO3NOItXZxGqAl4nw97VyC599krskcf7sds9SIyB7p7NWYl5ePDznQBWDTl
SnkbaUWcgtEwXX7233vtW++Ao/MqW28SQ/Bqy21NX8p1VSXq11om4dpNrPDEhdCKRrMUzcg20GDj
oionPnCZ5Y5H0U57DbqFLiNO3ufnLAW57epBG60Syepe5S0hRGEhiRyc8p4P754pR3CP/b8EjfBa
TnP8UCmJz8ofEs4NFGeE3ayZj/n4MPmRttQvWJWHUM9keZIi5ipDeg7mSdWihWMy4hDWFo++MSTw
Z9FT6rTTilfBWIZYDSbfD8p3UL4Fpe2rvtACSlWlQyS4Vv/RIgKwSB4+R1W9edXo1psOXxAfd9IP
Xia2g6cEprWZdrLqj5NmeU2F1B4sc8TXJWObQdenAb4TpylcMVmfOPSs1lsi6rPFMrAaYnYphn1R
SbmT2qED7j8qhtK5G6J0rO/FuMpAZlui9RDVakSBPCIh2WyZJttcMfjvyZ3svCblwWBotGsN5plW
NKRN0qo9m4/WZ7EkzcwhdV+m4TxCOYhKiNoroy1LR9rO2MRq1KVljt/LRZiQCLvCZ3wxIAjFytf8
Q7YT/Bp/II58FV8HT4KpMXp8ypNQnpM5tvgCBOPPURa6H3YT29emFYAss1MTwWllpcYjJcY2yRgn
HUiiCUWvp4tsKm7JfLCD6B8JkMW6xI1c7D2O2Ui9/PqKFAls0moVYa0gKY8ZS5QIjzOOqQAX+ZVV
YV27OhptblItbcglTxdjXpZ7PnjvKOV+jbz5JWSxlDXFMUaw3jAHB47LpDLNLbJpuiZeamJSQWOP
E9Evlozd5WIY3q+vNkWdx7mSBh80ZRT94WyrZMA4a+JUep9ragKMV4oR/qUDpGelA3R9+uD3asC2
1NYN8WQ3CkMlUpSSJzyVd+Km+LGUdvU3Xm5yZvwQxdtzkwhX9TTVFkAKUyV+I2unUp66sCQ1R878
gMiEZ5FAupGWXnrqUQIuPTsZQgYLDpPCR9eVc9CBT9YefeIwVv7CQm8GyoXrcUZkYMi8pSnzswaI
5gZb5lh+NgckY7PvKDO3/UH+gNFt3GKuu5DNRebHXgfNATNus9tv1QbrlHVMUa9FMxo6rL9egZoc
fr3GEF2byrRk8MrOYOLe73IwPU3hlITqZmT1Fk30Jo5bC2VGovg4gmP5A48xVTcj27xq2pwbjKsF
I+mMEek85NU4j+VWYil7dOSAV+5IC9d9MZdsywHSpe665rDveAQzK8KoFmSLO5QeBwga6DI4pbkK
lXpCF9FhmPHpiPQWyZmKj92ZOJVRaFNHfO3hCthuKIUD+pBpLmzzWY+j93uV3DET9MZdG3NuleQQ
9hRFzJVTVuyu41D+FgBO/o7xhi6x5zRX9olqezw43tCMeQESvF+MDAZJjBqg0zJDXO7Q8zVWOBzR
LXc0LRll94ZbLuzQCJGocweOf7sD94oYw0yY3C5nkMbrx47/Bw5ojsXoQhVWOTDj9jjOpiMQWU+s
tHKdjAdAyE67B8u4SLSt8zrmWQKRQ8RsSaUoVT4l5cgdUcjoY1hOLbEc8BEM0rGcpwC9JdrsM1RL
IqAnwr3FJpQvV4fvVCu+EM/pCbm5coibLR7Dr2rwYZd6mc+tkA3yyBW0VGa4XAtzS1ELrz/uhW7k
FGzYIyTSKbagoF0v+ygTdJuuecUEOT+fe++tiAjBrzO0I9zArPZSg4yJuyU4p6Q3+XAK1SbtrulC
l2F0uyesqKZK3Y6tWj2Y8t1R67huPs3c6oruSGbB4ZIgEg0isXsFYfcIBNmB6CZQiCTWf0hjF++m
gvZYG9Qx1sSdfNuKCj/AtFuBMAAGW/seeJrKclShismuacZYLvbsUiXRn1fat4HIHLoPo/ZLEmfU
lNBjCttdf0a/XLvR3DjaK3xYhYF9ML6T3R5pKFobtK5Nlt8q+PJ57AQ7Lcuq3m+QaPoIMUNDZozx
n/ql1O8jeMnm4udiLZjSYgPfQsmBp+RsZtkQN3mDNs0Ffgb0YYush+d1EpO5RgCVFodw1S5cedts
uCMOxZ4c+hLV1D0sdjlTT2ZaKttPkYt30NnAPdHUYBadHM/VL/Mw4ip6boaRzh49lSFvtO8ypYJb
QOWJDYJddNMJMsWVYUApol9Ig2VZchoWUScLxzYSDnXswFPcBtdtgaADXdrc+8tJtl5Az37/k9WI
1u8AsIWYFldEcCeibY4HzWf+3WBzgxUqL2yrnaMol3mXIEfe89OyW8AQOLD2PXNyeTq9e9MZul+r
cSIPWkoAMfulUbWGCqYNHns8leQR0Fscvaq6wZzYkL2JjniAHlZmxCDyBheHs6ifeJqZY4AcoVJW
/2WNjKaQKrz9rTrWCPFoRMox7ocLl4E0HaDxbU22C7sZBtB6xvqFqihKZwWaACVEsbHwhTvqwHdp
nehKOMVzVvfIiPdo00YAkojdfrF8tlca6Zz2yyBUBnPx2dSdngmgxPB+K0qg70wtO9M92ZOY+Tg3
svsgrPJq2+bGUnDGWmbZLRDq1K70XjGdzngEmHXNc+KZ5oGYx7inGc53vPLLN+I+hV2kxCeoB3JG
X7OH6K6OUIAJZbDDZk0DFInBY1LChUdlltpP21kxxp+/EJHGXB9DS3M+oK9uLML+1KMBjmqDx/lj
pOmPb1kazaiE2Hihjedx8tc0iHXd3CpZFt7g923XBSunATtXr60qUrQIq3KL9LEfXlCGDHDNSr3D
UzYww8wsxnx42vlnIxaoj8LW1iXEYLwosKw7MxEbmapouol/0oU8nLrgT3vO36kNH2ZwO6FBGDPs
We9kKANEHXU2BkSMKmUavOzvozWwfXSQL05fanf3LRZai/ZpzzIj6fOVv7MA+zAz03DWX/3o50ug
+mOLj+HQPvOm6H5LmbVLXSdUZqqYo+SWrjkrW7xZIUZpnpWdtdvd5sCupwWGVS/yNfvluf2NGBwD
JOBGemohoHUfAivL/PL808t1wiiWw3nL3cb5ueNPh/Lksqk6v7lBQAjX/Du9L8rbJYuwqROOaTTu
MVsWm9HxtGtiA9SZHaz2ZUhdRbVuXh5uz4PEE1NSsioivvOZ36Gn3h0g+wUqlbo6oo8vLARecv6c
tXe/N1SjAn4ACrdU+3dEElX6jpIqVzeppUnSuGW9VqZCi2K/oKapr6xSOo0hro5ovIGdWf7LbDmK
SwMp7SOEyhjG+J06yIDaLJJ+WTLDFMAHOmJr2RJMLqNv1Sd68eqSb9QOdiIYnGq4wK2H3k7RvS24
UxGD5z7+tbBcQpIV+wtBvXEd52+fndqlArETm5nz0FC+HmgySXuEbhabxW90ECC7CU/zI+pjdzYj
aaG3OAvLLpZTOvBoyW8BU5O0yvw+ypHMJjRwCYMG6q85+JXls2TjjYY+fX5yhDvuSkTpQrblwXeC
w+RJbDVfKwSWCQfZSrvVKp5Ux5lKkplc+xDg8nSvA1qUgiajjxmy6gI4tlDEAf4vss854nF+4m/a
WMc3xG1MsyVJ1xuxIPAc9LsxNONYNmriz7FFBaWmqfetExUuGMRS2UOaOql901rPZvAlpmFWaYbp
JZZxg5jLHJnPi4Sv6OHLdWftUW4wfrKFH7psvqyeaJHRt0x12dbiP8aJ05cxOxomZd9Qtgf5BHj9
UuXiRnOtkANlkr833WFYMIFryammh8PAe3kn4nN/yHYa8WijRYsmqUtMjiH01Hhbhxi5SXJJMerS
NMKYWPqJCvlouM+lt1TaagudA7SW2bIGdf9Wz+ZYYsekvY68wtNPf/frEfV8p3J3ngHhz+9PR/Pt
dDhj/5vB2GVFVQ6u/h8EbsuzhsNVse3io0f3y7lX2+mFJE2FU4B8pJHKQNSNsdteNcrFdg3JCdRE
fff6vMnE5L2oqCd1Ul+k+eGjuPJ8FxZ1jNU6LW5Eh2/Qa50/m4qPWl06yzUKudNK1BMeNud6kBfB
dA6NGgw4lHSgO4XZqnePPqxinzrOsG7L0rHFGi448dzyvFpnzIqHVDgaYv/Jx6Jl6VY41nFOIVoD
rUsw5kC9kdOwv2lJr8mlTC+a7zxekjjrwukqv32iBd1pryCef27E2bPuBP4fu4c/uj+PExxEbCBq
MLRpuBn8KH0rORb1TQJa1TDHRwYH12DBpw4xfMKnF/pmSupMbTWeEZSgPL+52jrkmKqzB6L7l2JL
fjQNKlESZTsLhehoC0ScpmVOnn833A3nhlr6B4ZyhkvAA4xXbVGftY7Qwrwsf2jk3AA9ZIVZszR/
xNdSqNZq2QEGz4XsDKsLAQCxdy9NhpDfd65IKD83TJjB3/ac0oZiNtseYiObVTIi44tUIOerI0u+
8FmSyYX0k4LWcCkRFEuSvT3/QVXMqADOla+p4/njhpFFmmklKkrMFpsDptBywjwk9WcZ56MuBBNq
bEhfpWg7foSzydbLpLlFB3d65J6JDLRVlKtunxgGnYHnQ692MIQwxVOWMAwkQPh0Pf9GGNZWG1Vn
qXJz3d8NKW/I9NBxNO6UQFRbvtljuj4j4gWc7AVwtU//y1dSANp/2TvubCr6sW/PlwDpfoclJpXf
bEpxOXDf+BoY6vI/s41IO1AYZC0Cbf2WgaQffSioJ0WjypX1Nk/Q5QRgJliYvG4sJp8JfAYynoeK
l42fSfl5xSgFxX2kDRipHNxy2gJ546S/nCJKwA3egZjhQxs8oOO98ddckKcsCUo4KrB8AY4tb2k0
3xq8aiU8Ioo7q3fH+UcPY13fP65nymV5pFeTk7chJ5d+r6/tOuY6uVszatva+wWUXKoq64DV1uJr
+yCvHLyfmzkG9GBkQcZRgdUxyfh/p0g/MCnWF4wCVm4wb+xWDyrYMePA1H8nym0bev2evL+b27QG
M5QyRxlzTwise16CyiVTVHHvha4dJg6P9o2Q5J0Zo12x8hX7I7zjwUXfnjYv9X0GINEZUhPBf+IE
xLBl0kP4JU7sR8m4qOdDjwshJ67/aHJeRzM41PTe0ldDkQGVWlJZsZfTOzUzG1LUe0kxzDPnckVp
NDxgFQu9IiHaTfsJaD9DPGCf/bqnEGT2OnWWiGvpGsiVZOFTTo9KDorX/bRiBbt1XqsWcC+uy5Hn
Nq2mwjs8BtHqU/ZeJH2HuWXV/zF9hXpp1q18NNqL347iMNNNNlfKuHogrROVnjRu8jHLdeDkhPfN
qog7VFWkgcOY81gRXDQ8SqzidVzH9d2/pIiiSxnBpv5FM3yxfJAjVQt8Aukaez5U2oUdVnp1otqP
D8mEFpjq5xSOFnP2xXcHNqTeM2+x7cV91NaAt5AWn4HVExeSZbMuxVX9VRdCjq9JAElyiZkSSMZP
BAE7p0yyPwvnSkEhjt2PNukrYbMo1/ifpEavEvO34cEC1NJtF/3aSh4ZBA8LxT3UmtJsYfnPKHFN
knzvfaPXmIWcTHKfkAb0gPf8TDCn0RrYcL3RKELmT+Zw3WeOyhufI0g+TTMASG+FNo6N1I2NkFxd
hquFqwM+w43DDOFPbNaGV+IgnkBHWrsW0f9vgcENZVDXXcikDpst8CHUokLotBVRNHiclejKkPc3
MoTipY8YCzAXQty1gdklbZcIZ/e3kDENc4PjQIwb57urWZiYu9hzGepeO337gHy2z/PFmS++Gsqz
kKeaV4Sh2EG/LCBTOwD1rz58Fvb/OQGRNgGK4S3+sSLx5XuqSoqXG0Ydy4lVGGv3QC6xhR47mI1h
t+1TisFoq90cyUfuOplBrks0mXxMCRujXmYbJW5hr+x+UZGdZT26fjrZyHUFbzMiIMYU5+0+p1dJ
ud9qaeUWaM0rJgYbfwu0499/JMD+7RQOUvtovqOdOft35Cp1bDC1vawKD+jCBXEpTi60HXuwzhRT
KyaTbeMmJ5Rts3Dwl0WWUoImRNrT4sCMk0XMWEVbEDgHz7G3lgzgNJDrQExTadwA7zbnWL3+loY0
PRxQXXupswxhH/cI5OBVCFueEEWYGkqJ76mbvZklSl9o5mtod1uUnoJojP3NrOpdYlnpelAOAyQc
S1DNciwPjHTC/O2gk8fvt6teE/ewDm2BZl+0qHE4wQQSugWjU9afZ+si48mAPLopu5RfVkMT/A5E
J+tNWtlULfZwajTU329Fhp0lQyX+uxZBmxBT5HLzFf/BDAbo8UZh2FhleC5XdBUKe3eHt2zgUZgT
0npLpw5m+lG/f6KcGVfgmQf4QAh+runaZyiTnrb2RvpECpMSsVkNAmEKswrQth02aIIjlZIX3Brg
IL0/JB/Yxp/GKrW3rKjPEx3EM4Dng8MdUnM+iJukZ0zjRdQG9YRWZ6gXlrjjkAAeL0O2Gr6T3oHb
cP6ZT6F57Ru2+RdgPY8SnCj1BSl+tL2S7QnTu/fF+IccQGTT9tZJDEB9Net8zlPhGYDea40sTwXo
gZfFcHDO79RwZMcVXP06CUKWDFclNTHVOsQLelI0cXq8sfyid8BNppwRCVq51sOBExWdIQ/xPXSt
VCOM9Obcvp0RdJOcN6agesLzP+toApEuVuA4UfK87kAKdpTJ7ULaGLRDTPnahytBW6/DoWp3OlDT
9nrKcslghP9GWQHaVh81LF7HcwQsWAlC6QNYRNJ8lz8tiQssCHAxAMcjgd9snB9WVPwQPoZF2A5g
zcX9/+Y2VndnFSWdwR071VrVMFWsa84WZjUlDrtdym3gbwtEcoWNAdApRWiDhQi7aG7Ul/5BaSRk
0Dlvi//FGqB5vkQ9U/7RuzGjzqtuPicepHnNHXGAcFoRAQKdgdoY67llvxA5/Ni+VKYwVzzTvtMi
KdGuRfbG7jDpDN0IhACNOdZ5v9fQk0Ka2B8+jEmtRpd+stKa17F2XA/Gav/lbkzUOsqyG6whvtix
hwx8l1qgiSfJe7Yn8K6UQI7FxRzB3Q1ywcV59ej156brAB2D77CKbAj4AOC0Bf17DUh9W2HdAaoK
ilmHB4vjph8elH6EFRfFCRiVPcC0qRldizmsZEO/ooHPwu2Ri4ykZY48joRIvypBqYhLnbQ4kQVd
HlhVGPQuN+MPUxG3SkzvnSSO8CRyEhPQda43VNQgUyi4c2xjuXdDuUNh9m1kViq0Sz+TXk7/cMBc
QQp1qwdFRRZnFxZUQVvxH7e+G+fadaKIhq2jv7gIVzxQvGd4ngc2zzflFFWCoqJyxiGb9yem19VG
PAgzi1Z9WT27nEHrbhnWvu1iSQHv2vTb80CqrYYjklQP5Xhj06H+9uJKRYCHufbXPvrQPx9ZiO6+
JW0qSpuAmfxPQdvdbCToPGKwokSzN0iI0ysDM1grxmGiZX4DPN45exifZf4m3zL7Bt9HY4M9wIQo
VvKpi4xh2omXL57Tuuock1Y6Unfs7ulQEe4IrDtd7w8zXUu+i3fahguhaYsyd+dkRLEdyqDvwb7w
NZRaJJTRSCPAeDNNMzDvWVHxBtLiJbxQUXnn4R16evrWS1NcM/eS96EQe7pd0+4DNIqBSgLo8KmY
m0W43/sTOdIWidfyv5faw7OhUM+Dpc06mvgLRPqU94FxbyF+k6Sg68wXGQlp2GQ/MeOx+nkSuQwN
y5vNbIagVp/IQ6mUrMhanhC3qyh0D4G4p5Tq7AoGI6bQnn4XzGw+DvQ/DHAGYq+L2LYDqmlmlMUy
Tg0CS4A79hDByDmP0kdtfBCLfC/TY7P/i+ZNMk7xpRh4kYSs8rnStRcWDEIqe0vt9jGvw+hYzWyr
bNfdtpRbWk/fhcyXXHgI0rnVQBzDy0I5/zNyEcsSfGmC+B2nmpIMeI847zQrniZzRPCf6aoQmrFi
/FdXFtRsktasDx9vXUeZbS0AWvmcCDMAtKeGJYNvSQga8nVZ3bJhkGSWoPYLsMlv14WpGKF7Tuyy
1Ydh0knKS1kFMph7+kyK6SoG5Eal20y5jx0gn/nmpXaJFR0GJ88DrwIH+JgObOV5/h7ra8mdE1U6
M9plLhnjnGYBmIWvjFAH34kEeuyYkmvFd6lPFdmzkd2SX70pYwevIn0/UBZ3v80Qu/oxUCoNlhQt
Uwcl/gWqEan+Bu/TVpeVruOxM4eh6KaOM9UaB2QPQbjBIJIF0o7H/t9/zG4y1u5wFVCq+vbEP2x1
VEBu5x+kus75XXe/EUl0ZeAfRjTnPapxmVJL8Jauhu/7wbBnxXfBdPmJMIgfoM9vGM59SS0FZ1Ox
+gezjnYRiCUWaGr7Ck1C7qdBNQHWQgppDoi3x2tUaumGrkguftDjTq4Y7uJhkiXtOrF3KRkD33C2
MPqGF3yxoWjLIlVluk4ZNiCLeA9rUY5QHaUPbCc7ztdeMwulwtS6HiMNBrM5b0e2goLU2mbgav2Q
Y1MhnjNvSdcEsQmM0DBgmQYzehvrJNGztprTIeVR/4lGnAZbxwQFUY/6kvx2mPF5ZIo/wiC6/4tB
l1Szg33k47CRxu4f7THjtS8yukQBS1hPxR8nVKG3xefgwpxIdW3/MsY+vqXLT7lDAbqgysiRhy7V
l31PNvlrx6OWoaKwcVFWEFU7yxbvzPGcLZ4Yz3hmQwMBx0Nn3/Tqt/4gvh5ytvEAs2a0YyIxsqM6
Ak2so51nkIP0gBUZpXOYHd9BERxXEyl2jUtVRDvW/MEGGS1bjvWtiUnat+/Y7UlGeefLIX/R9wcs
Y2HN3Kafcxh6BzUjqHj7V72NnmA9UFS9kHxeUQih5DJypc3Vs3JdWeugxAY9x+H6WllAWZe9pfIu
QkLgeKm6OfMxRuW0ARyN20R7qm7QeaqHU2FsxWoG72jsBvWipFGuyrU9z4LIw6ftx7z4qQ2IT1QH
iN5IK4Uwz5W/1Z3DGwDR5AsA+H6XJRrqKqrQQRBmJNENUndXZVH3+DDMPH5w9J7mrPc8CrqxXBF0
SlryvJ6LWDZkRPBH1jEYP0RjyU0cX2q6zIuYvsh+gsSJb5bwqZi/IBEQ5ZtllDJxy/4OtCi9JE2u
WuFEZnf9LGw9TbLOHU7T7UMIMWjbTcm1SYKuIkw+/TsEAYHwUspAfMnMTDtqOOpiFB4Xa4RC96tq
kk0pVrb9p6IPSAfx9XzBSZMAbBu8ahtitfgxQ3p7o34wXUlhN1lcX4rVZ+hexPekpf4ez6Au4Sts
mGwjU3IdKqpgkk/FMhuwl1qRNn35vhU4+oH7W7u8w46c7xYxXCCdMp+wMMMENOBlXuZ2LYBX8Y9V
2eUPZToMykuT9nJWng9y2jskyyTKm6hcRVjuMrQFDLtkDmwNdOOckhtnyKW2X3AfcBVuCVln7jb+
JwGUej+8913lsRJpsDb+cbig5yu7FZhfxEj5CoNBNl6LHvhJ+XMj8e5d4xsCDfZc1Zuzk/REycFG
NF1UcPGDqcu9F/gO7czUwUDDTCsuinvWW8xamR9HM2q42dg6QFownWCt/PE0x2Z73mYdg1y65zq/
ut6fJiU4ewHdG+ki7Fv2q4U4U+3GLKAR6cD7YJHGTcTEKtcMVXpfTrQBafSvTA7h9JfjE+TVXzcX
sBeP/Qx/mfBO3/IVjxR6UYApF2oxkYyGC8yFkx/QzanXK3HSkTrA3Q268cZTTLN9NOfvTP1wuGKm
s83MEPmOLrOXCulQGHkhpqgAakZvY0aJ0eAi8SuIJmv4G/2qiFF7BFw4l4kV48zUlp39RBopk4gz
H4eSfvhVno4APl+of8X5SMoFFPwVk+ZVTS3otNzmBXB4QSSca5q48LyBNBpS3TQ9UlczG9oIZ3rd
8oA7MOdE7FJdNCt0fJTXSH7e5mXA+MafEZzo/4wlEcSY23yBALKNCtVN4o3Rbo6RPc0s0FtEaR0x
m7BdtB87AtUHv8nAF29pGGxEQS6FWkYn//9HEowRcO2TQDgPaujtWB43sMU6MLOFjDMfSJze6MIm
iquBFBF4bwObXaIkuhoMCMdJP61suvpy5/4T2Wu3Q0DrW0Ja71s1MMDwwtoDnBCdQpR6O7DDU8Q1
0y//id6ISLucyrEIW280MRDySv3VLa9jTcVr021gtr0q0q9IQCkHkTyjRAIIbvNPKBLXU0IMEIUa
YWT5Sk8ux9Hmh4qQwoynhQ9N8Wrdri/d85Dtm6a3GALW7v3roJkd2/ilyyjkLM3b5oQmHfP6g46S
AQ8yP+PIOEUySJY/3WH71Vb/PFVQqmTe5Xp4ck90DJWBNZ7ikFoXhno4xJv20ydU18fxr4Lf4lyy
0lsusKiSRySBFwy8wjFl/aI+kfFuTdHVrKOkvEGy6ZwgKlHDMXNCjTN4NYvdtQyN4ftIkU6AYFXM
03MhdT1bFJ07W+q0umprXh4LPU4tHJbP5sao2FXwoa8MADgKbq4pU2FnttFV2z6/7dj5yifAh1Cd
wnF4Ln5mRPsshyiAx836iYn9z9jTJmmPUYJwYnCuIcbV67OMda4t+X4J/I+AtaPHWrfmrhNIV5ZY
sVPRCwdn7a2UD3lQGfmfBRGqoyyYLmmBFCAZITZuMX3LvP6zZ3vF8WIC3h+0ijT3jxSiqNOnz3MR
86OLZH/Da1mjo3HkNVo14JNJ3afT8aGLSRHHTR4ZOyRchztQlTux8ExHdwFQaXCSqO3Sgm/Hduw4
mkLta4QfXlup+SFjdDSPwhKiV9FcY4kC6TlrxReD4U4JP8VwfVOAnp7LBa2D7jTXkkrpEfa/02gs
5a00NRmubVJADsNcyiBsUtSDbTc0gwMEXlDmwJmjj0akczA8xT1lFX2mn+GT2jnIdFpzOjqp9aZE
OZJiMQXGnZguNUJZy0MxwWkTTvRITehXFedwgyu+Q+yxlK/cYShNkJc0LF6Y2V/JM8b1vAsOusKU
kfYvQFLfS5eYg/M+BpVRLgwxP5AK9AsCDi6D3dGFCEoR2X0rrVJ364UGtzlZun6A9W39R3B4NjXG
e18RzOKQQ3hGqauuwbkuj4BQBv7k8VRywk2ynjU9lLTMRZQgdSpS355RUekqO2MdvzcyCGtkgPkT
IXaT9clhDan52xV7gHm4xr1UYxaFlwsQvvIHbECrBpQR2vbdemP4MDKeLpFFui7rQtcFIedKc3+1
KFIomogyTA+UGMerCkQ0yoG3WrO6tZPAPxdSrN0TOyO4NVkst6tQI5xoDnCmML5uZ+LqWoL4YlYu
Afb3ZhBcLzhBBxJDRWTJumDYr0VJdGBdcMfTRs9fI0TKm70d+0MAHXJJZhuTNz6nOoUiX6Xfgw6j
Gf9utsLL2Y/KlpsgnfDd1pqNnOF3NdyWe9s8OF6rmf5X1H2TTG1X5ifBg2yKCAM36Yc+uxPoXtb/
A6RXSJs94drRiwpiNfYCd5ngJMnQYFq5/s0TLzT5kTmGKKIXf1cLsKKEF95pnAMZZ1eDovKdonr9
jKLnL4Qf/m6F/h4jw9+UwWDOVJro1z8/E2NyJVyWY6os33C9usLt6kO4JO41bltnuZVMwI0Xp7xO
RxyO6tNUWSrJ1z4pIrOG/8HW0MGdEfhk1XdBxQQfNBuLDbeNpbRpMMywQYKGW8gBJ1pxgoNj4x63
R+o5rWxueRmtSJ4leYxjMI3nydG2hniSYQL/FSQBMawWZ2sJ9dbe1NaFC0/xJlrHqRWghbrYKXDY
0dk87I31MugBMWbCl0VFxecxyNXEc68yEvEYSfRLGMAE8fIVUNvm/ZVyw30mD5o8WAJ+YHOMFzBZ
c9njw5QI27W2cLqLJ2Azx0vKqBOMnfGcgI5CO7NCr38tNgLyZu8RPRJmzauPbDl0NsNDtMtmRcWH
N6AHg3fTUx+af03FkWL1qg6m8SwAz8YkeJC1xaZZx6Z+1oNX9XSAP46fCcR/FaUWcV8w02WZOFaN
oK90BHLzoMEF+/FDWGXeJq36oc/0Lp7vqNprZZ10ifcionf/TRweexaWnBuYFCLfhYqAKLLAjaaj
IjaV7q6RVCpT/rbSyAyNU3maG59/EFzaMqnMEFZ7Ea3NSvEorHQQ5f58pxPzU19DcdAultpIKyhA
D3uq/JcFgqjeuMXafY6iE/iMa6RBB9cIcuke2006p9EyxVUYsLH9ubunfIEuNRUmS19PDXkFRwWm
6co3Ocumy/8V3opnzkez1/zVjcy8fotMTlCQHj+WsECYl9/FPGlFXuQwk4ZfWwtNPkqzK4PD0vC2
tUi/wVRuXFUeTCfAF7y4dBSn+Asw3ZqZJVFuXxFql/LwYAa7w26JJfuDRV4KkCdg2lQFdB2UrnwJ
X3VuJ8Rrtzp9E3L48aicdhwPme4qxWwfY0+fEkmvzsdVT4Tdn+aXB+iweFWG0KeoKWQyaaAyjNjH
HG9iRpntWZsqYDygiOUAVkT/WDZCB+tpDsalZTzE9zhrtjVe2nF/0xQ6G9f62qSx+7GhXPyktE2G
k815LhFPKYRuCGUXTvs9JjhI3Pu/7iKs+i7oAkt2LrXdEmyj+jy2848cu6slRLrrjh6P7y2dLpRV
uQimLcEUky75VQDdV7+Pkf0F27dq8PUGhCR0PERPzWubUF+PuPQ2NW4WPlFUaQ4iVHgmfsI1OgRA
8Sjqe1c82dNReT1JNjlSuGVYBsLAjEoQhXVPkpJITmCOemc2uUP+dxA+Z5K/gScEwMDjq/omnUlH
ZjsP1T3AHKs+WC0CyB0VQUict0zavT1yuGOy4AaQna91vyOX6N7+90FWmZRFvG9ZaCdRDr+2bG3B
z9W1bLr6TGTnGWSf/AAz8Ctt5BTESeKYW2ItT7bNGS7GxU1FsiIVyhMkUJHgCkzRs+SwAjmgwTIp
eYOdQ2Z10UnVfR+ktbovAJc/zpHXXmqt1Jg2zw0ZqepExLB2So8gXPf5ImSjxQ00DdxX+n00wkte
pFr81taKn5TL+HIKajiMoPYdr+Ok8jh353yjPjYr+QmBtPec4P6Q6/chxqm0qfeRByRqe+kyAwzM
JkH7mlYNMqqRnrtjo8ozXv3+fKq0LofmPC2a9jrqFFnsYIbt+E661uPQ/MNcNep8i9AKSMsox+Kn
AlJL5rfdjFZ4Tiye5OHvPczWOEg3WiFnzneE7F2TUaJhZdIz2M0EpErheW43jzpc88FHBOYw9E0J
XhnI0rxbDeuzLKlUtH32erkwDIKv9cd+JDhWzUnA0PoakN+fYZex6eUGcztmK3UGvMn5YXkyXdk6
WgdB5LxFL9zGdHB2frmaJu8TNJsxGuJ3xqFPPf6aljBWlx0cp0fP0Bv5/nU+t82Zz/KGYTmEjALs
0fSYj4kAmbEas3rmzNumsyQv1rOJ2SaoJeDkTSp4SrAKAA3gvr8TySQiD4HgncTQ0C/+l/shkNqM
sqIOJEqXN5Ur+S4YN+yk0RCYNkpYnk2sKk6F+X5tLA4Gbp/fcQD+PCpQ/xFoerYiqpKP+OZkoich
6fnbgT1YHx9rQNK5jaCqtZxG6cqwuzoVEB4BUK1jw0w80gJ5VnJ543U8gyKQDSTX9ojqc6v/g5Ob
xVlxVtvZEMxScFtOfQfYyh3t/vd6UqceHQn3eGXeLMwf3KLIBEvFar4t2jD6kQaF9bRMY+MO5hY2
yeHJoeCk8yDDjodGxzv2XveyCDbNuSo1413aO6V9ZkptN/hlZJaCXutQmynKRKbzvD/HGc4dMYmN
i8SR3wTzBE9F3ulc376bgl1Ir/Fz5M66vZWYiy2aABuIsivtSyD5YoG8h3LkF+IfFBN7dqFGFiun
HR0tX4irEHjxo41YSulgxzX55qEoT7xc+KBS8OEWcXIxONzWY518BFILaeekaURrUEj7HAnpW8Zw
alcxu3zc2Up6eY4g7q+0xZeNjF6a1aAuRHmvLveXX6gcrLPme/uka1AUsGfG7Jxz7M2cQrepf6cp
ERInHt8ymHipb33x5KziWFvknPMJX9Gyrr1KH2hzbooflTm/uvS3/jjoSSfsHPJ/QwcsnxuPvgh4
lA46FVqmf9XMrrXi0Z/WXbz0cLRhTZbmxKpp0RevrKyxpd6kb2O1q9/U8fTaA62vYk/ZXEZLFY5U
Hfa+z/u/kSwNwRyxsXkhZ99mGWQ+2R0qhQDXCRyCPsz0L/A1C5xlLu1C6V9UGM9xEMmLc2OQ5gfu
1pf2/5AH7501MnFuKbRXc5a8oo31Zajq3og5LFL6nEx9DT4LsEfUxOBf+u7Z7k/xnbHoUkGN9oQw
AqoJQVAUa2JUcwgcaZlfkmEm6maNwviDDTMgtKtcvdoHYR5kSZwa+gg3l5H/Gbn/GbpyQRDnJ2aV
L4QF+ekbtiSA/9LUoQ/8xp5a3SH5ueD25REj4Qi2uvhTcqH2UxKuf/+lI8PH/ngpNAsWJg+7TQDy
9kj1f2OHPRLzHUbZeeuDhPhkiDttJ9SWLSk+xj0+uqe3D5OEeE3GJR7NJIZUW88oC9gS3vg2Y5Ww
QAxxQSV+Tx+IrRwCEEsp3yZGxrLukGTD+42YjIZGa9s0eoo8uS/STZgGtXm2INXcuinl8tIFgzWu
7C27RlCCkOESQsMi0XkoflTvEf2KXbK/snfwNFMhUMaQzDNCVDGjhQFZpN20MFrOsY/oEqMypEu4
2HFH1fSr6zuqb3AIwmZDV0szqsM49o6zEQqfTMWd7b87ukXEwtt9UXEkpoGIbD688v5cdK4CyP5x
bF26oBGJjFxm713twzB24PikJ/gHYCRJe+L5XJpPehx9FmGr09qb0xhxdbcFiJjVe4i4C3TGv3q3
UJ9NMJBSjnSQxctqD/ugvzw+PM+88+R4sYTJzU473OzyV+wlLnHoBtOyG9fhcGhPF9IYws3K+Iqo
SOJUH2ka/p9A8Yqxm1Koyu2BSsIyPVoOLApg2PpAEwmlKXei/eir+EzgJf5XDctzSzgkwGlK65m7
fVmqspUR24iwA1evdJXuo2DjMjTZem+VYU80PS6palnXhJKFqfbDf1XbnOumwm517uBoBwS4vcQ1
gNFQhx3UwS5o/fjzHeb6BAJ/0cEkXZKHJUAxdhtGw6cisRxNiOEBp7lFIsBzwLZQlyfyM+w0+tKz
LiZ9RLK7SaIwAP8JFTDHZiyyJ4PQgforaPf2FBA6Ruj6cMSlBZgLNDE6I0qU+hqLBvhOfoj4qHF6
CY0nvQVuKnDBLsgStvxrOIyNe1r2vOtlv4EmZPOJwJ7hfWLNs7HYHj+nDNhlkRnf6oNuxY7gzJyC
aZhCG7CnTSIhFesNQNo63E0FjUtNUsxYCtHsFJuclN6vfe6GaBOnTdKKkl00GZfjiNoAbHcjFFX0
uI2t7XdP+FhVa2Y1J1kYgUpoIr2R+Y67GAFA8kxR/WmdUPiqd717mcsdwyJ8sbP/iHr/A2lxc/Sw
LnzZJhT9j1bzFL7Yz6vy/TjPTCzWL4z/JfyQb49f78qJKxzpc5fiOEuortDYpp1RI2OzLjtODsGt
AeWBXgfqlqSojwTLERp5CXbg0/2f3yYQ/YebCo8O+bMAy07Z5R0CieqioSI/ARNJ5hsOcm3U673a
J1ShoukjZIQEljlqcq2XM5WQNK/poG/gKFz0NPt35rb4I2wegkHEDAVtUn6djNeuELu5NdehghZw
lQNAPDS7UFrj68OoZry7EpOUxHZML2Q1TwotN83aVaECsUshPNqRiscDMqkPCOUzvjtV6LImMqQW
sKxHH2bUmGAUvfprq/k3l978FH12EkgE6D8ZJwTu5EGBnHWE70NQi3XWEm+Rc/HAUXoWzO8c/QC0
BzIttS5Rd/W+rcr9zKG7q3kHzLv3yQTHKHJtMmWmP3U6pIQXJb/CqKKOG8fdDWT29iipolr0I8YW
lWKISLP6TJiwefW8scHqSGKH/BD7P3qwiI7ER/Pdl0ODhY/y14iBrybGUP9SVzZdcNckISI8Hwcp
1SMgbdSZ7+h4BL87gCYp2NxY20IBxEzcry1xHx0W4h0kr+3uGBGkUgA4nCTGIgkj/j1120w69DGT
o/zqCPPDChoAHkQ+Lw2DFojyJZQyDySo3XP9S6Il6VtsMxI4UOib+2e1bMpo9Y08bK/F35ri9YOq
5wsetkOd5PpMa6tMpTOXmp22OEwT0hu5Ao2mBni8C3oWRbhdb6vYGmdPTdQHQBPw37jYbdPSkNPz
AwzbYjgF27ydVpr489sU4So3r8DyAh9Cw5CQRQ2AU1JTcqz6QewtXskFqNMVSX0wyhSVkmQehcZJ
4k7+uls/FnNosuhtiY7DSIc9EuF2bq1KYB9TUFQy9GIYLOE9dkWx4ew27lM/dlgVA0FQlRN8jRHH
w8e48tKdYv6HBpc3LEg5OowwV2dFhCoUJQsGKH6KmKmpgnn/TM6p5dZwP2eWwCovT1KCS89yKecH
CMiT9zIxUebGfOa635Om+LD2osl1gNDAvmpMlhjDwzqMiIuoUeqitrXQAVTx+0bmcJ5y030SSnMw
vdH5/WrXMf17ooTOAoXDeSRFOBjqMc0QHIZzkp60vjKUs+32ErmaUCvIYknqZ8aUtFpzuypiWe8g
CrNGHFHYHpFWWNN+SVTcpxQdUo1bl2O+FQdZpc8ws/HuBl9dEkr3d5CRouBKA5TlCSyUSkhuNVtm
ZBqP4/0YQjfqfahDASI5gW0mMxBqv2xzD62GleA3IBG8OnkGlwiE2GsbrgWFjJBzpFcd25xLlCrA
N8jXIyXnRSJ+l1exyrZnCKApbgcWDErVlRMGY4nSsvi7p4/dUoyPbfnK0qQxTn0KTNKuP61UQd+6
pKFJC3vb/QdTGdWjGe/NHtMmNfn7dqXU60OUz+b+8PIZOUP6VGgl728rTKkfvC7aZAM+HODAlAPV
k1/ZXeqd6Go+5qMFoa/i+2phBZMP6lTrfmAKZfnBc2Sr144+Mkbe+AUPwtxjzEdLhtsCFYG+5z8K
ilCNgnCMIt4hdVXtf+w5kqIqvt+SMhmTuYlU90kjI8m/hi2VkDF/0K9Im66qc18rLShpHma/cBdV
KPP1Pnz6wlXQm3KlLZwmKzrqYQhjtGOl1KjYPbA0Hz+1CG7mvf+atmkTsZYCDNsKgt2Q19NduqOB
UKEZDt//hCJmwTarfdKuW0XsXZi+OnUlHLM7chiel7CIdWnojfgfsYGUnlPPuaS6JAMW9TlRo1xV
boVS/LSg1V8/tfwdIoYjsLCuCberv9kRt1YSsenvdVKyEmexXzJaDknTyjmkyCDRwFUeJ9hSPxWa
UnsU1E7hWy0rAOsLp15ruZX/8Pj7aKvU6X3fk3Ch0hGypL4rJZ14cNsvut/ouzP+ZJHrn6RjBHDS
wlnzbgMMzjcQtGqHX4bHy+aNrd1/fvJEpzA0uK/hrKdHLQznO72JU545qm3jI54SNJjJfNUTFkfK
1GCEw8uQ4ERfnQhW5xjG6ElesE8KC3tZ/PNgStvfVutmErHIHsqlmoV4oz5r7RESkkFSR/CCMtOf
uhYMf4Y1dMGY2XHVxg3K/VxFZM39mYqMtw3rScgv70mMWX1xGEXBodYnkJ7jFEmi+/93Jny7/hgH
BwjdYRt439ce0Dwm7PyNjR40FGXsRQpTnAdqvRc96g7Q9Nc/notdM00TcoyvLh/7o/8m4TTuFUW9
Wp3QR1lmK0Dan8kZijHgsektwO/QaV0CEMC2Lqh2blF5Uexf1QLR3PCVRcnieVGyQOSGRCBaO17s
OcDPEABC6KDU2A4ozqiov+TRoFEO70WXtxMCqnhl2pl9ErlK+/LKeNF43In9juxIBsG+cGKoBumD
NWuPdmvDjRVezlDf4J/Fpyz2ZUfwh2Nw3VIW5/UMJo51U6du9m3Y0g6rzzACq1lfT/4ZwdAoowWX
0bWJLXN/rbYt26nhyg2guAnUNh0VRk9EPzD2D/Cd9CbtIlNds/+qGdk1wELTtQJDRkK3BnJxLzOU
m03rVI6JtZTRBVtm/xaEw9J6gdGZDEtxCtOQSzkt6vIz/6ebiz/GnGiPJWq5kCkpSH3G023kvdCT
0ZMh5LhVH+GCQBlfIRRWY85w1AYrGmcM7v9y2Eq8oIZvjOMIVLEh6X+ce9KXCqR1r6DptmDgUAIX
+Fv1rBd5kx/+luuaew+Yg/EybLGaQpHIs6QqG0AqHqzC6dIss2+Ww5PH85wh7NmgekbNJXu7WmJi
SSrIdce27T1VkcQGbQc6zsSVpHJEI3OuoRF9vKXB2CDjnRWaJB/lpYYDyCL05C5JyLMJ/UyKJPXC
A6kODJfUtrPxQMFoS4bbWqpmPH0mU9+eoEzpk//MnWyRCLy58rVVYgcgZrRe8xZirHknlj+5PiCG
27Q0fpqHs93E/niYT23hjhdr2G6IqZ7tTtz6+C+7fS6c/tI0wmiS0eOW5A7W27aGH2PN3872/HSy
7i6cG9chs4RbpOcpdwirU3kHhZQyM6o6ZxjNRCLqwqw5PSX3CwUb0/Ps5d8ORuTbeoCwbRY/MFKB
4M0fnv6JcNTnA/8IVOR5VLc/xf/GQrQK12J7VhvTg9963V3Bqw/Ckd6VBeV+FXgNITu6B0wBo45P
dLNeui2nyY16OC2OcvG2n9yI/usZ8Fm5siBI3tZZZN3w6GKeIUrUyhFcvAP6vPXX0hz2hw6spE4m
tvJm6GJ9eEVHgp7/qx35TCsbwlgOoV/kIB/wVljiHsm5RzasQ5EGsnuXD1yGTv0/uXY8lep1j7Hp
kGcQl9Y0yB0+Eb7bP1SF+aF/PPxF/gYG/AdTcJI5DvxdxAVu9cV2ry9NcBrVY8VmCiOEsSGnOCBK
WwT3cE0cyFTsIubivOi8VH7ptNKAca2MjD/nbNRE0f66WxORt9Pum0T/Hljpyp5lp9dY+lM0qKd1
WVbkXyOT235vHdjrCHwNwJ4XfoEb0vutHN2Axwp1L6NeTh+kpARneFBJsUKWvplqkZH1fzbgBhwM
VH6ernKrK39emjcCLEps0mP8bwfi0NHb35hBeuKcmvL5+hImKCkpWZgFeW7f+JzggmWObcWLLAYX
Zuf14+tzI1YdNxviJtwl8KiV9MSYnU+LV/fSABKi0yhRzLmiOiXUDcQsn0ucu6GXVyOz8X948pkA
tJl5pgmmqXkck/J+VoSlj0DURTvKDaCLDwi0HCSHQh4m8zYQo7Zkl7mLs1zCdIDcVzyfnAs3E+3o
ivA8+BDyUhf5FcoUFX1euT0sJf6KEhda1HssXoO2+2Er/AHrwkWeUWUX8u2xgfyF3g0r9SKS0g3k
XuRc83yAMHOn68pdmjQ4hn0r1RsN8Y68BlkuWo5jdctcc6kJEG+eRBT//c3C6cguloxjdprbIWK7
bgjMj2f4CZ6mNrcpPSUcFKZovVtVwHTzEQ/AQgtvn0XYQ6cOIK6pfBFc6I97sa93jFewpHEhVqGN
+hnsPPFyVCBgip2AOYDymqdG4E/S0s73PBqb50jRlqtHk0MgHOPIQkqBnam9ONlIZIX54RFawUA/
2PkLi+rdEjzaB9vrtCqLbCClmHdNJkISziYVA9XjmB7gzGHmmCb2DJGdtY7aw7n2MT1GFmJDv/aq
lm2HM481QaSbNHNe8GdJKx961w7uZQz5mX1uWPbMbR6ui9/2w6chN9E+MTs/TvjB5L38EkN/6z9U
cwF+N0E/ATX8M+ZqiTT0m5ORkJlwNeEOenD2ar7L98/isExgJGXBHDoUkR9SU3AsWqDkdtS4lf9c
rolBb0qh/4FlvSPjS/oiZwJ6sYbaMmRwnSh/9gHyH02oYcNv4CHpHV6LiNtiq9FIRPq74/+e1yUX
hZuC7b228JTrIXjNd8j+L5bI02UFstIY5Oi1pPLGxkFJgauWifQJWcPhFkl+zLBbkvAlZ3vf3z/N
eUUtNmz5co5V+VNoQnZQjN64kLuPKelb2FaC23iq+rpb8jdxrrQJua2QMUH3FDbQrmg0IyolpkiW
3QNwwThnOgTLZ1ABMkked198EgZiTmQsDNaH8aXLrKK2hfC7VIOqYx4G+bagCthlz0r5hHpZ7J87
qxtJFUKjB7xHUA3/uDU1vfIufOKpF7GTs6Zf8bE1cyxSIdJuvYctgP3vtuhVyX125HxpWalrIwdl
BFfDsgM47f/vQVfFjki0lSd+LNgP7X2bR1eW3CKUZZHDYmjkvYUco/3k5ExUTI/iL4iy3bQi053t
PqEkoIQsi8KYn2eP+R8pkmvL4pQy00kHVybbycmeYrRD3y6yDam6GTtUzPYgw9CgEplbnfily3jP
dXqAh6OQ8ePIBfFY4mVIKxB4Rg3nLkYLc4vRcR1b+1pUd8jwJ95yBfKub1qHjhQo0DDxj13Lat+R
lFlD6enL5txZvx6cGuDSbnF4DwaHO25KYLZ3sbbvS5U8ei3EQAym53Hbe92E9WIxfLVzKfLTVp4S
Xa+1DQny9tOOFzz4vSqvRSOoR04sXQ8AHjN4wq7nv6//p2Z3tpNs5KeKXtzWKxU1mKa7+Y3lhUiN
H1PiHVkP+B0XGO67hQUdfkhfC5KYXljDDA78IxvSCHMYLRHY3aqtSAB04Clr1fKwgdq+SRykTNrL
eKUHaZTXZAY1LEoKoXGAYAQr1MqiiSmqRSIOR/Aknm8xqYsxEZkI4qiDtP8yVOMsqy9/xiTrIUlU
U5ZQXQ1pylzFYBsppjntxSjYAsI3oq3WQaCl+NT69AmW924dZuAetcd9GKuyMrvgX9WuG+dGdIpe
OeGaQHjfhTTDv9GjcyH++arrroU6twqojR5LACib4sejUqQhBqmMVrQ5ukkBQEwx6cPgydDXke4G
LzktJ0s4hYZS5Q8RLO2W/9P8sd3SuEQ0qsqhoowH6fZ1P18UQghRchIUtoK9wP3wpZtrQHRKTx+z
uL5TALf4MU4cyGMm1vggReLJGZnAB8jRb9h3AevrXvxeN2gHFtuNsUXRcwEHs7kwsmWtzmbDsW1I
aA2PibuQRX1q//URz6NrV3IcgITbfVp4oP+CAH6HWbXW+UJ4yoQPp4jRFjv2yjZ1LHpbofr0dobP
YbSPEG+9nH2tEhHdd2qYOPbMhbUO++5M+sAwWnhzbhw5AyAlgWkLs+olSj5hWYRU/4klN57u1QTZ
F33Pn8paI2VnNapRfziyVvsB4ggc6y8p/4iRwsszavSBsFNGEe92k0zlg6J9mNHlxVDDRiN5QGKg
ylBoEILgjC/AZm4k/tBVBXzsSvuIiF/Etg/WXrw7yOHkpIyaxcHkzZDT3ufWCJa/m/B9hRVJ/qE0
VTZLrwC/t+Vfvy0LE5dLBCzWu/EcU9T+ULINbEYTqzSCkM6CY1mtt0qZ2clklu6IqWjpDZx4eqV3
Ed0wy2TlW7aBuNWi2awnPZ6dJtbXQFEyD31KoImkeUgTMs6pJeBbtX0zUjgPW+D6ObYpT46ELSHz
YNR6dKKrIzHsCg2hvhKwhDTkw0636DNjJsDy7NOl/fq754+kGEBPjWtxZ8UETYZ2SKvSA7+AsCkI
pcBynVynivDk6xdlvAWiGAmOkdb2gCaqPCAaJetcUe83G5kRR9ETJwKREkFmFDRhDK6FuM6NQngy
0BO1cjbSsPF0rRUCZEPwL1cCKbZxejHp9T6z1TvgvprCGUeGLaXgVIieVQI2x1k1LsiMuqTnz0/5
hXBdUiTRUVyNa/CZQoKFbYtR2J0uzZd/8lxh7JiRYvhkABeiqEF+JeJw3WGaG1ZizlqMjB69V2T7
yJ0RFhlDm/ydtZoYTxfGCWUz6AQoynlDUM1elFbvYfR9rK0kw1//LaYVx/97rrFJVcuwVSAWQlE/
QkZ32dHa0lUtb+ujGWJDi2GdOsVWzSy8bPeAKqFwEhJ7dtAjUyFoqBXEk8qKfhvRw4CgOEeB0XYQ
m1+CGrFoJgWQV2V/wQtlSVyTKQtK59N003uQhIKRRLsyEnaW45ACoD3RrhvNTLBgb2nQ5G7v06do
0aJ30D0mpBP6FJDNfB83VpBsm8SQNmJakqeAttLB1LHj1CUvK6ZdsPo8qLGCqoDRXV98SNd2I8xX
TJlXX6QH2IdRIHw5oEz5MvpJ41rxA8dJ3WvwxI3xidifEdolNvy78KRaftLttBEJz20OGLwAX649
a+RBHAGMndolovQ2XBzetjZd1LRE9MHNZ/wIr7y4qxSv06evd/DY1rIE+WUN9p/4AI9WaW7hc4k6
KMJZ+njmE6zsuBbH25t0eJzml1nim4H2itQlWSvbtVxOz5WTueNiYYGh1SGS8rwH0UBnChZ7Qvoi
RS9Z5yP0Kmo3o9LVnvVgvd+XmhkR9eKGTYO4jsaEswA9HX+wXpOhgC6jdsUPOyLfuQmlmg2o5US4
N77u08PCO1CPBH2rHtMarnaFaClw2AqyQvosT13fCWN4HmrRikTur+mxGHsbSJZHVSiZYpJcXDNc
1BwRsUSGLhW4ghxsJxOZeNIVwazvKYPaL2ktRXII26rCAU7swMFKnUYlWr4wOfrg5qpos3/knDL9
foW7kcDe5LzriqugtLFnEoK5dfHPb3SOKIk5zfzODidytIkuoxDQ+jOnMuYsH8pVZd/pDRWUy8CT
W4I7eTlY5HJLQg3Q2I7f7KlLvOvHk66XHx7KtGIQNIu+F6r6YtvCBlHRWXa6ClaD08Yn+sY7JGFd
hT+V59s+E7PWhBIW2UPIY2pRjKkrUnNG321fr6Gqhp+60tKa3SJ3PLt00KJe9kBuheNboiXEwvG2
hpBNkP/pGc0qn0qf5CdCTqjxGP5DSYiWFwVg1UPgA6tN6ToICFiKyR7rXW8QWdt5YaWgPqUiEprH
COob4acSOsHt27WQO+amXMqhnd5Fyk913MacmAPYbJKiwFkSS9McsUhSVRWj0NFKdyTMGMTzWog2
TS0Slz7dF+xA6lY8oM3CTkxgKPpNPvgTMS8CkhIm+azNEgf+RBqstKmPnLYn/nfqH+Qqnl8GZjtt
JOAW5YoOSXI44fGrEKEE+PW4gGCO+cUKOcU9m0tYODmqcCZKPEpHuuDKOU4JzOpCK74+8kY3u1oT
bJtFuNmtEEhASnVBbWLa53xsERr3YJSaL2WmSbk4M/9kU0aPNDPDCL908ILRW1a70fPoO5ilzVYT
/qaOaoOmNMw6U19Ho+hOM0a/hxZY1Wwp/FePBf8qYazUKZJNPpAMZn6Q2ppZA5YU73m20xq+i2z0
fls1jEIDEmg+feG4Xl7DezJmELxlyp0/uNt6UpcVP0aptgyI+8UB3LXv2qQv+WVgZ8pywe82MfUc
FCdB7B58jxbzRWeA/riYW6jkHqDxwi+66k9XgiEG6bP7eDjLukYl8mZuuOGuJ/vAx8MwEzCQEw08
ktMf0JSpsFj7MGorMkZh29PYhjKgzDFtPSC57xirt4AWbzj/WdNL6iUyh8zW9TY+ug6/4qh+I/ii
Q6l0vJR2n18d+ujI2tTDygRvufTr8iD55Ik2gc+s2bzySPNMFxJPiHQ/PFmLnQhkAV6hu1nbzcnw
+xdPdxGIfBH0/CCGNFSP/m3UXADq6mvnbrTshyJnks+SZ7bTaA+VcY+2MaQYz177EK6UgdAerAKy
zzYhFcu1tNv3eBsaWhwnRtOVq0ZHTexc5ebKfIcRwsJ/YzeaU/oNAPaj/jx6M2pI2LqQfo7vGUgn
TDyvGUFChXhGqd2gQszgW6vrKjBRYy+v07oGN51rwawRyg8sS3ZLg2Am+JZPzT/HXj6Yuwr0r5dI
D30IrWe+JmqLmzuo+VyKu3XnFjkLBX3++dZmyT94LGzDCv9skzm6wC8foVikgtuBa+x7pFVLqszx
HSixU8PN3fkoGgP3YXeaFOglOINFRJhFMiaD9NjrnIns2Dk99Hpzql5z3aGC5YJ40nt3s8o3g5Zw
XrO6nRvJ/TV90KHC/79o2dKLbCDYkcn/LhPEjZkAaaz24dTgDZYtw8YHgG132S4VM+td0fTBmmZB
gAAfLafM/Ps3A1JgYJ24X2DlLo2vlNkU0JjNLqA5O0b+jswIDiX4Q4uZ9KGkI+TlkLX+AGGTNrI/
p261ncBJGMLV975MqFkiSwX65E7C8t+PeT+pVBuUI6t+BnccNdxI9VM+chWi0IqzM457uPkz+9HC
W7uZuNJH++t3WgFO+nBzRpng4xiVlsE7x9SvqojJArWfz+C6it4FAnhUUsnPbbT8WRuNX23SAXck
QQk+5KR/epTdyvUB7o8wHPUpJFerQrP5p+1nCDiW89a3416/7RQjIxA6NTcSDuyNDJ9HmPprMdwa
My97hB38uOOxJIeZGHD/Mtmm2jUqlyPL1ADcNnwSc0PVJdi1EhNLCB1tKtZFNE3H4cdRzv1lBXEM
wh7qcF9gPstarIaGAfsm3BK8GSWYuM6JFal4vwz3LaerfdA6ejG+TtnY8HLnBnLqdl/NhJOOwqSa
ZZ3xVKEP42VvNRTTvhY1xSfinKz8CZ4prGSl8XIbe6r3/U8iyuQJVPd7J5pr4pBmIqgoUtf8sgxJ
CdEgK6ehYcrTR3o/r3enkr1ooULBdpSICDXMol3GrbjW2WgJM1t5QzH5Xd50a7M2SVYz5JF27CtK
V1O+Lro0VjNL1BxFMCkp3ttW9hV9flDI8RInuBtFLE9h8dKa3n/Nd3BNMicizHIZguuBu2QOgxB4
zCKNkn8I41AY1bqs/Uo4BvK4R0c02MM5Wpv94bBU6+4TB8RL1hIp/Kw8Dn9H6rEo2BMixhUIKipb
PF/x2K7N2In/PqWhpoc/n4KGli7Qh8b41Ci91TV6Pm0xwCOl2nQ3DWqCMK2LAOohAfBIffmpKzYZ
H3VRSyi8TY+NLamyr2jkLzw6ZC+wK082WTuolz7rpeQRzDzlBil2LspjNdhFq3Ka36ZQ/2sH8vjh
iolzkvORQMDJ9Z/4HSCJpCnHfkadQGZXokzy8qKHo57WNGa/8+whJQpiIx1/KDO+4QrOQI2ywJ3d
HrXwSPxiH3FvbwxkUumUHQTRqNM4YqqVDXNeOzmm1wHMmuZm1iX47FCWJHfvKag98iecVxkyPaU5
hlWf+UxBsGGOMdj9hYtGbkwcHcJdr+PbWjRb/IIylLISrFR5lMg9ED5551SRQO3Qw4OIgs2OAzTF
lnn/XG+iDNIF3RvtsA7rc8ENUKIlFeOS082XUzSL/xGOz/kJ02rEPPi/58OOUWTG0YSZdj3KRj5D
81QZnziQ00mBsxtnZHBCVTfkuNNvZ7IitXAHPL7WF0zztoC2Kr8PIVcqFJW2FddK19sFIPWppila
B7XBl1anehVNa9DZ0I10Tq0YbYlq9aHuSll7MhIkDPL73pfj6FU/fwDw45DWV/Keph0Yq6/IKMn1
R+lzNjYAYTjuRGGZuy2s3pkrmLsolOfeV7Aw7jG87MA5Ja5IWX29s/Ijwysw+4tQLL2xvshvNgIN
ZdMCEfvkAhLAxbwObF7gK4tIDSw71fcuBVcs9Pm3EpRJS4lYPYEE9cmij6GxGfKv+2zvJrX8z008
hUv3BETInH9qDBfj5Q/qYH5YB00vS7btUrNtE+Pii5SJG97QEEeRY3p+RKolAJIW45A90ioJOZIr
Lczp0Ht4L2bw3kUOyLMA8Cg80vhVo7hw9OHHFWHKP7u/Tp7yi514nSHpciNklKprBiyodgq8BOE8
uXVvFJNlZFj2rFW88/uYPAv+aBDL26atKCcHNIKDjC8puA+duGxnPYA4NryN6Etcn/49caO4Bjke
2kcfZoeshHsegJZ416UgJvg3WaPmw3tQWOtg8jx89LUDLs2bITar6f6B7fa9ROYo+KXPeL7Sk/1V
SJk/lDUYusvf2BLB3ykt3x2mi0mIUnflp+vmZfO0v4851K533pDT0XRxIZnhKqwhKaGAP9jPpOwy
K5VDzoYsg3fnzBemxNuNDHSRX1p7KsRAvMc/jsCjdAHlnO+dsK0jjtB66QYc7qW3ykCGvucby86M
+d4c3hzl/psP+VCdanScVBD54TvM1Jhxow7T0wSncWDfttv5d3t23EebmbO1IpBEN4jqtilrIAc0
lNNYvRXPZsxf9VLN2I/0bGLGw/9Os2mEEzATRkYzwhUcMSk96z2IvXjTplXpbwESrRDhJETPacdD
8+MP+aY5TR7K+VcTCvZA7uSVjKN/DZXABfA1Ddjbd9N1H7wO9iTcat3kjzqHCqz2cLsX/4ft0cLG
izxJLkpbAKotq7RYPBzBDcwjDcZ3yxdAZSO32seoq2AYNhU+V8nAyUpauhBCVCcnkBYG6M2wwzMV
nAw4eCK2UdvyHW0SHqlKLtJD8ayUxdEVIgu/LVprwKkQP1JRwRUgAT+rtR2p3MFyWwGeFh/Xpc/L
699epKfWJrZU+31XkfEirFi4ybZjfZUytUG4xSL1K7/F4EZVhfqGds0A39u0MOCtRXnuuiX/4vEh
1fFzZh6eMLEfytFJZk3A6LlVqMLzJhhUDySAXOVJF/aFpOkdvTXKrIZJwZ1e83PBtIEYM9rye0RJ
mPzl974R69h7knPz1nesknlh959h/4aSiCNqzFhu1nZfF3gEa0tz1sjN/5BLq/cgE18yLbf2EvlK
2IyAJSQz/1rt8BkRxaUo4fp9GV3cNvkm6bTBV8S+OhjytNfc9Ydf0hHPkL5QPubqirtk1NMeiuLk
k3h5DXZA46fERu9uhGHcyVDoTzNN3JclMElkL06AGMGAXgAy06GhNs1waiAeLe66FVYHZvRZppbU
Lba7m12bNnCklLBV/CdFgfJ4z6bFkTzfY/x0oyG1N9nHOlx01HtqibSxfTyouITXTYdvNCo4luol
00lZJhctpvGZUd14J/iOzjNMLjsURTSFWEOemLuBguDIPKLs0hvgmMCBv71qN4c/0wsOz5/pcKlg
ykvS6lHICCehWl1P+ykLr7D5mXxk2VEGdHB+sB++yPO9q0f0naKXqMs4O+Q0L95MSe7/T+gDlJx4
H3s47kSfxDfp60t8zhanvchpnvqTd3R07Iraa/JaGHYGqs+Sa3Hlem0sDKjd1XZU5rBItCwFYDeD
q6GiptcQ2P8FMEt9r7TlKmfu7UDS9GbkFocsbFAWVlNuROXa8+nOP/CTN5OrIyZc/OaRUEGehO34
csMa6BYLk8lnSOqNDQy5BPf3Q1P4s/QS57K7QkCV/54W3Xi5aG6WxPyK7mn8kTYe/tg8hsv5p+c8
WCxqOLCfL+8E4pGIY3MMtTiXddTWSCH1LUWZ6FoGF7WaLU3E+NKTsQVHzfYfY7+l9AW+gYv4wZ0n
qxlyvoDDPsk1NZQvixSlbBhvZpJSm++LTgGboIpPUFTHWn6iEM0Kzrf03uNCw2o58fxNJtf9FEa1
Yeqcr4vUxzq2yRBcB9K3ajcyk4odOyWlJKGA9drIZY9mYTmIystafUvC2d+/gxPuFidFQaPQdNAV
tZETSklP9jvs+kt7QUSqZypxGmJfQvfNqDo2JmQxggQGqL4MaeehOZNeyP0vdC1hmOViAyDxGpYh
8eZHZTzqllDWCcMhSfkS55TpH6xEKzy/cOxxf2hjEJqVPLkbiZzFbCUexUoQ93nBwSpOY2FU6a0A
XMDR0PEqymSsBQ+7w2jW+DTFaprQXVC1TA9jd+SVT74ak295cATPe3EijNPCXA9frcd2fCsH1Vjw
6ndrt8u4aNa3KQ9vdYnzMbLr1M2tdyBOUCo+yEB3O/VhVioco1FPtod42Sy23dD7v30oIWsKt3/T
UStUOpiYPiiOZztwyg04DpXw2NkOX5NeP09yA2XBJUC1Lde7Aae19AUc2J3SAwku1NtPaR0ULx+/
R/mjiXJry15FET2Q8C8ami48aDDaoe1n7ypy6JioiwrA34BvyPYzlVWnj99ul/a5u9iDFWsVDCZR
AMuuDAKhOCFrtF7ba3tKzFuwF+LALoxdCj0bPLumqWGawJmOTWWAuEQCcUuuo8BKUOB5++md6Lfw
K9t33Fx750FO8Oofy/z3nW0kzAvBeWGmKEbCj1b0kMQn2yFeFQUZrl/2Pomx+FCp3NMYLjcQZHqG
Bu1P4UxC32YZUbzuWyL2mx567sKcXwU2n8U6FnK9RKLo/CqVOU1xKM11oilbToqX3CvTl3xGV1A0
7PHR/Y1icQvHpPNF/A0RIeV8ymM9f5BGwWS2Y78Au1pYDXVldVpZiAdC6kl7kpfZjGz85oVQKc5e
DEzrIwLuSitVYuorLqIiu37RCycVUeOx4VsamuD/R5tfXBkEjFI6LGUrVdAVNbrHGlZaCcCOR5sd
n/hOi9bG10GSs/XJId/191YPSfaj+eyFgPhWMFWOit6iVJi5LjBSFhFsUd1QJ/XyfJJOTXeJToNL
wR0AP0/UqxQwGh6+BkG3kmjDbs5bSf5bWpXbKASCYufAPFdpD82yQhEUkBSeYmFl5tuiRCOfGF8D
SXfCxVCYicsKP4c0JmB+q0ayr8m9PNsSAsy0wflLGeN+R3Mb+xE75oLWwOQ4DVs09CUXjcNlM6pA
+9kFqJXi+aJKE3akaY4sU5vnMW/5El8N3H2xW08Jn9kyB6VJlO2DLR3DjdaedLSxtbcfs8TRqD+S
OqbNEp5ujYPu7PJUR31gWEmJHJtTdl8c868b9R0gHK9itS8RU6KssDwTZQSxgx1nVD5+0o4OFQok
IL1CV/9ICWhdr6pmv9nvu4jKtrSjnp/DZ3j+CQcalWM5Rmsegy8Hu/nDER5qiiy0322TczTB3z8f
PxScvCwgNYQRMDTUhe1DB6en91V0OLI0c4te3MyZ6FdFkD4IhIY/EBPKxH9zIbI9Ws60VUYTa12A
xZBKuYwTXFiDlzMBETwj4rRrKJsRAFMzibhR+p1N+Kdzpg/eZPvEUgMTyx+MFx3lYgDFZMgOPhsR
X49Fsi9HT7g1PqACSqyAzp6iMdYJtyoRnRwNbLQT/9aPy1MChiFfn8cB3l7/krgqEqMQVWwvZ5HN
aRpIAURujoruXpq8WfUdUSLlGgPScjMr6BENlGYhQg4sQHDT7f5BwIMBslbAqz7MFMjaawM0WlvK
T1TjZqdT/dZbJcFwOGKtcaBhryYAiipaJbvghcVLKCyTBJ49jbdCnL18Mv/scdCeYKsm0foXeu0C
bgkzIyd8AtGdNVBbMhULoNLMbfrhTUHk/Dwdhgoz6fvAS71SngogrAe5EGQlKOk7Ycx65k9e7UBJ
VwK34yu0DJc6uGa/IgAVkScKF5wRMnWN9dlUe0R8DarxA2gV/C/pkb+0/x26f7eC4wuQB76P2/ym
6mqCURdmH9VRyrrGvrPVhB5T2NpbjCsIerS4acfNzFs1LMg/SSnRBIOe3+U0cjVreznDTDpn32zD
+AppjwfvnqtH2wJn4Tq4sd4c+F6P7YFWwxqRcn+ok2WBrVIb9+S8FMh5AFUuLHyhCI1qHTG2oNbk
9nvMCBr7vx5ilUE/sJckfrZu+mXK1zl9MGFXt8hVW4FznR6aqJ3kxBOo+kWJHLvi0E4xVvd//l/P
yiRtqzxFyNBPt/QJH4njKA88CQfTcV2bB54Mn5WJcoysy0EnC671uFhheKxm8DF8KX2feRFo8Kdx
2Fc/vliOKwsFpnJJ0yDdq3AE1Oc37LRIFQKn/IswS5ftlikou8qXBnKuGP2WZ5TbH66Ou7dsmH2v
xsGsQEdt9u+ogPJd9+FoawCnqj7etSt10zzGLil8kIfqmVrJswjWWLM4cMdMOGql/1LicYEQIsyM
VJdb2+dTq2u+1Pt1t1Fwy+v6hmr5P80CvXl3M6fWuLPAPSV5RZcHhrfH4lnZLebW+T7jk4CZWmh3
g9xI2w/TJXmlpr2G3gnTKZmxumhlvcl/s3EzTN7MtjV0QOeQepnf7+Ey3CwHShCAaqUUeLGVQpI3
xv96R1DO9gp9rnSOcsLqgE3zNogrme4uqO/zC5VnMoOXWHJ2JfYtsS1/7Pz+N3F3E6VCflEL4O2r
B5ynNjIhuwvyh0I4iNr7QygGWO5XRevKMHmFIe75s2ap/QEXBGbanZn5LkzmRkNPua2ncKcT9dGW
Vee1H2aGDK0TqHmyWh2RFyi8MqJPNLfNzFVnVV5m6Uk+VD1JP4gC5eTMlJOE0J9JBr1+bY9nvxOr
ZNIy9/0KD5rGsyQL1DRuUqJ+ho/gkbp1YyeuSq7DR7KI8VJlU+5MpoPOfKw8ogK5+8VlgCHx+1HB
VCnO1E5V8QEDMDlSug4zcWLhoQ0KIoM2zwR7ca6L/USy1nGaR6ZAbqkdibmOif2c8eWCijsnqIjL
zrb4/R+Zvmt0dTsMaWZY2bStOKcUm21Ao92wY9yfuSPFJmeXS546YAEsOQLwwI/mCW2b+dvSK37D
wTvgsQ6HnBu2ZywP5cofFHoZKaggwpckua4jYwYBGJmxPxKRmMgrpL4NWuqxtYSDs4KmjioWLzuA
J8ZDp93lUkbCWeJNlDfuGr+/s4oCMGQSxb/c2WCZcHLQ2m5siMY93wIcbGgmlMNI1wcJZWfx4Ggk
00h5WgbtSypLwvcPaNAxB350reiSuXrgcBiDZ0/hRmbDjCyOW96hviCSAJaDiuein3wwl57ShEu1
1cV3dU+k5OAZ+kreLH6yUcT0fXeR4tP1MubZnL4S3VvZqnsCB6hbc/h4gtt9jy+dbkFPp0+tk7AC
N422PMa9+ntMTa3mKgv7iBhDB0Z10khDdysH2yVHrZH5bV8qZ0E5c6s0orAzEV4TlOj/v1oKfe2O
0xUiw9e36ADzo+u5n5ttcw0EhMGVZWcQhzdFQT9SYiTHRcfKuM0SZYppoT9+jQ5Pkfosc9h8N3Ba
alUfhbdAMF3/fO+d0zEAPvrE359lKu2X+Herl70cvYVayIc0BcSySo1bDEnIbAWcwW9Uw3o+Xpbq
LtoR8x75JNvDQ/FKUP+b8mqDNrdaD3wuwyFAJ/61Y7qWeulWzUMNPVwUdfWZQNIUrkGaSDf59izd
EMHhQl23zVMtdavB7Tm7K45EO8d/eunvib43TtqUwWJlWmZhaoRUJzAAyGdPj85ID7Cbhj0fVOq1
nqvMQ+0T2qBpOVVWZ7XZ4ikB4nqUHmWeuhAdIL0yCYWfe8OhdX5R8eYwbvljn3KsFh0JFHp94fhK
NxLUD3E1VhRX0qw+3+Ljzn4qFtcPJWjEMqteF/zahx4/OSe21opmzvyyyLGiVcix6B4g6fWGtzJK
DNoKoxiriEYAMECopcsYpbbOkCjcTshIG6MtGAr8IqHh1Mm2Za9JAMs98PLi+dV1CNWyhbATRPxo
PabukPNgrXuc3quECsldAr2IY7+cbCzfREzcH3RQBS77EZR4HHuawoMpryD18kG9zt0aeteS6OM/
5NvCwnl3ts5LYo6CfFtHYV2CVsmqqoovInZAgvoJR19P929UAH5iAp0y3FHUQvJR0TwIVxSkchpk
shjRuCtfg1/NvFdx3fgmSWAht6bjOjsJ3zBHPskug4PVyOtSIe1p8MNk2mBQKaNeEvoNdnDd6RWk
rYGg5JkWeG7IOkopqcW9a8eeW6h7MhEd1BUug3UtJU6XRaKW9w3PJ0DXEwXot1qhm+O5e/mqek0F
qHoNe3pPadye7sXKF2R68g9WQiaZtQ/6VaXIppZ2TDw/Z10q/obQf8SiR91atAp6rLWn0l40Zb+E
gIwxdvI3lUp2gQe+l47jzHzhcRViLue1sZFd+6m+nbLVv+UcUXZf9mb4Wl0UEh9tH49TgSa+XIY/
1Vxo79dOZxgdxxJbIqFSxXA17xrxt+gGPSkuVcxvLNaUX9JUvh1RVTKGalYqd5ja5/nEV3Z9WZLP
mYwo+1YDWIkRnW0iUEWwwtu4rT2DV3kXBOyU9fX6aAYjxao17+2oCTuIYNZqGr4JunliaXNoEuxb
EZcfIZvFrQNqvdgUi8/JUJqXTwgauRA2XU7w3UoJR0R3Hc9LbjGz0ems5zzjEltYlMQFYQJ2An0R
B4e9keNDsBGD/r4bxxBzeFnb6ZjjcFcYBBp6+jgdoHkynwju9ivFkUPZOT88Pc9t6WtpqndtroIV
1uthaW58MjCfI2X7M8Nhnptko6R1ZVnqlgukh2tB/GVBBcGedckPFLRwCxY90F8IOmJfjp+p9Vo0
QoxAad3HN3q2X0XB/Kw8j1lCO9T1VhvEU+0I7RndehD5IHonJqt2Cw/RAJZMgj9VH/2of1MSceNc
DUs/Br2h3oEetrPp4EH3PbV6jeIcn+gAq6Jl1fWr+TE/wU1RgJOTCFuvnSm71fqzTiES/6H09QOv
or7co/m8FYY8hedDazf2Tcc9V0xVJb4XBqRsxINedXA43Fmrx6HgS0FAZ+b5XM8IDLAgG/haWmxz
xjN9ESzxwjyuNxX9lJgdLUx3OT9kX1WFmP2fRFjkKmtlKp1Oy3M3oV/A1Uy2MWnVtIBijYho1NVX
Pd9+C8dcfLjlFJhFoGffbw3ixJW8ZB5h0YpH5UMcOxF243O5DmRpgkrJAB6jXvlQYgV/nHDtx7F8
kglKbxzzJEiga05zk+iK+mMyUICNZWOLG1cecfXJ5M3DKz8mc1bY5wcIDOXs7mdbLgSKwn8kucUr
Sya1+5lF/YYo3sdfxm6ICGktmNmq5v8G2bg6NOZyVvyP6DVBeEBZVUOyBb0IJdog65cZsOsK2gwI
KoYmpYz2lsZJL3k59M63D8HaU3l2Ebw2JElFEZnz4Bq7TI9azdEyfPdkd67N0OpjzvbarVvAl1Ke
2j9hF4mH9qLBWxAPWbpVmkk06BYGSQjPQ61ErT53/KlZTKikC9KPRT+8AMtQWuI1rozZV+ZdyJt/
clS7Q+Nn7SrDP9WliV4o+v22Nu0glKaIE4a57K/YojCvFi3zX0JyB2kAIGfM3csya2I3JCquInrB
Pw5q1T4Nba8GiDbxf06e7Bb/dbAqP3Q2TEvDrRZU1Fqf/kxXF4+y4e5X8HRqy5/z+NhZ8f6YABeY
tM7IiTXpgjnT/8ucU8yBeKptHzPdlKKetO851TvO/vNQcHv4pbO96CubwfPuRPEVt5RODGPflxQz
c+LHKVriCaX5skogQm8BEOdiVzuhle2YxuuCIwPw4T5r30GSevhYWXrl3xTUHY0JNUL9MhD2iNdI
oA4k15yWMnAQEg5MIjCxYF39zpQzSMp46N/lYZdQF+EGGMVU/teLyOpBmSwpySiNkWmYaIbwovb3
7br/xAe7LBlL73XGSVhf0x5yPbbl8xVlQLJovmMGq6rA1Gt0/sIGwDYnj6ijl+D2IQbHupvSx7Ta
EubYpjgRkNU9amjQ3LG52Gaxg7+PHNY9/taEAv3DKTpsvCyoBOz/WNTq71JVc4HxZZaCgvvtbKGL
ZjIZaoCwszjoTxMVoc0pkLdYu2Z8ZEdMjWrbB8NJrIhhbSZCShx9DK4zGKNR57CI73z8cUk3ERik
bO1SU8KFHc/QoFjwNDfeW5ibzVEbrt8MOC094BEyFZ8yjZ24cuskPfBBim8n47V3aL6fqfcqRcWA
ZX16G2zag5kpIjsbgGxkJhRRC86NtPn8xZg33XQeB3u+/tf1g9Oj22CrNKWgEDnCuBLMz1TnQliS
/+H7CmAPG/gIUb7Z1d/wQb62R7RoEAoa/tqVWqREgsYIcp+iazXG7goYpmhYvGFPe4YMRDYYgt79
YCAwqgrLyekK/01j/a3t+sJGqad8Jkw+sq3BP7RNqTxdO5120Mjyrylc+Y9936empJJGHkyntHSf
GKh6JMmRYGCk658O+vDd/V/9gBynO2tKH1FvLPIvwLX0/bDsKsKwbW6H5eKmGv9LfLO5QgGhhwkK
79UNfLuuubmDeQtu7qaHRhwo4FzewNcfUX4yUemyQGPgHRE+7nq00Wa6icGr6Ze5EsP36bniAy3d
ng/VwSy8TiZgXcIZ4u7png+ex9iwV1CKw0dPEEBgqBRYgTS9UlRq9xuccsiy5YtM+yy/8YGXzGNL
zh172DT9+ecVpYWqAE4D1X+3euR9a7oAF3KrlRTsLCAb0HjB3bpAn8UkkshbQsfcOT2TaKzw6QG1
PzRkj5IGhSwin/ltrZOWR+XzYXdOpDM5xr5zT83/oOZYZiG+BEeBQxZaOKGVaU4s6Ar8WbhyM2zH
bWwMYbVEfua20tjvXRCN3Ocdlzhfc0+NSimaSf0PRgUOKDOj/DGp9RorsHTNMFPgMcttb/MM/cv5
vq5qcgtLpFQgM7u+i9lirqjEL7nz9q+WugljgUyNfkhLXXuUjPZeRL7/WKLuevpd17OYshl+2+TH
tnCy8bwL7nh9lNHugKMDzgD8FpSLUigXPTpeN+3c+hdzXWEMbCaGq9zExec7fCw4tkIUK4b3okKQ
/8gflm7vsHhQV3k/UaeOPY4L1f1iWOjkcUFS2kx9xBLoMAWdL9+VrbFMecmORS0WZhGsKpJCJtRx
RvzRDMmxuJo9sEa3SVFpJA3s/2AYdv6pnjyzYXZsi6kaWdulicBqHjf1TjPMhCkAmAInHgn25TuG
1YnsozkHGIf3TRlb4wtOvZCBrki5NNr5R8YSsF6qIdkIvJ34Pr2eFK7oeaFeqQ27YKZMnul3OyT/
eR1Q2v9FiwhFbSADyg2bUPTxmWB2xeGTjvTo5mRsWkIuBR5+jC/Wen9ZASxiHZeumxYGVUtkdg44
WREPq5A6zNmnY7mttfATFytnYvoOACnjLwoSoad5Lo1jQ0k7/0yKxalzxaFerzFLHmGYXjBturpi
ButykWhjB/tyIF4jbjIcCu8o7BvhwvvRAEjPqH37wjgBh7DuAJdGVmcCxEZwMf4vlZ9dgWedDFHn
bEtEM7fiSKUAchVZjwdbpZqlouroYwCX9gOiHRINbwXJO+X4zELOWbx0xfdTk446i0wyZOQH2ssc
I2lNtixxelPm0CDSK0/GL6YaXe/bSDiufDEgTmv2tNab6KKBM0PfC71CcagDqM1Ac1JGk7qXB/iw
qH93aelYhaKB2oCDyYabRUJhIFj5u49P/5sH3ewd5hXvN21iT2ZbUfyLqecc/dKgCczD3hXoE2DB
nfLvIHxh3WRwXgnQqELLm/jQrxywQT8ea/ZI/0MyE9dv1OdlQxtjmgAwAbxH7pzsixB8xvVZFUc4
jjJ6CIDLQWRa8Se+08DwFX9l7HtS98YdTbYeoEqxYwGP/TFGI9H+IVIKuYqYNYlc+p2yqRVA+Mim
GM3/4ft8+jSE2Dxv38we0F656slpijIIXubOdRrBqsFMu3oEG5fr/HpmmHLuJv0rKjj84xicawsv
2l4lw2gNoZeu5nRxELkjpheOwKN2KhPneH218Q4p6QTOTBjdq7JfAuQeNeu8JOmbfOpdQDetJ1oj
TQPalcjr3XH0QUXaDEFxE4WTjsSX5Pvu2Kuak3CwnzLBeZTaTcMt5wsldLoJPwU4jN0Y9FI672fA
WFbBQ5MQrxlCps/dCWWwF+K+eG+xPdg47twSlizfyXIdqplxgUlYG/UeBMJ7aGwBPgFGsCFcbjpu
4muIBOxh3/mW8qhOLn35LIaM0XKY4wUIItcjmAEkxRNYuxGuLd87a4drJiPgxxJPK7t+NPl1MYYO
K7qfjCLjWraIqwDmMGLsN2wP+p0Wd/JjpGMCZjzqThc507wcMPuyS18YXSRwXn2tYSZAyWDq6p8n
l90wNC4f1H4KuhWBt0KYVPK0PRrZtZGCp2w97+ZZ843qyow+J7AhO/vV0hCnwot6imxodDS5Zvfd
HOKUR9YNF/DF9ieUxF3fhB45peUjqWYCs/2xSsy0ajhp/4/kyCgKkBPqaF7X5WPt+dBRhc9/475f
lrOxrqYolePVF1v1ffDS11GoU7DLu2Rj5lc/sisB+58beCP6m887WNQ84oOq/r7ZKHESh/HRoMTx
Z8Jjox5Imh9Xge7G91gqziVwg4Be+x8845YyEmEOXUOFeRHcHAPE23XyXBUhoBn1EcpXkar3vVRQ
Xcd4RZB7RXN7eFDyuudz8gwu7qjJXefJ1ScGPb7ok8I2nXFhj7xxWmGDDAi0d991QdnWCmFTNa9Z
VMzSpg1YrUy8C65AUduxFIoXP5Re79DOnjPN6XNzSBI0TrhjK3EGCWZw9OBplld7PrkmD3/CzJE/
M5G4jJHQLIeP8H2bgfbaee6ko1Frt78RSg+yYEY6B0OkpNlzIFqHLiK7cfBcLLLibvng5me1jCca
0NOM2/wUxznpQKOa3jmOZEDN3eLqqkum61Xkyes2fd2BVAChkdCZndvYXSZNEFdC5Qny/463zruK
xCd0dPVOdkdQ5Q0tm2t6tpIXTeZhneSfoWW24xfRO7uReql8xTDNXGsc0u8Wgpz6j/VIVEKPalIX
gKXXlLiVxdKk5q4NwoLCIVaAMtYls2un0UMNasy5b+fGuU+1zQfnzYTvdIQisDN+fRyL0caUKbOX
PN1vT5Q+jrS5+DRlisUwbbegi9KTjmF69POeAlB//YOKaRB4wwlUTCt6Vldv0qO6woMqXpTLkp9R
5EeXFBJvmKpC423V8l9Ehonh0aOiy/tjByFgjFx8YFTrCm2Ooc1ksrdd8gwgbBqlNpzWCpHCE2qk
yHEDEkbpqLMuhfHDV46RQQ6HtWEFMxdHNrz8hWGQwJmf4gjwanY/B6YgRKVTvnR9ebfGu/ckFJ1A
wsvOH+NZiTQ68KpOaj+1m95mUO/t9h5bzImckBcE7D10+PqSW1g8WmYmm4XnI57tE5ZR/LqZROUN
G3G9t28tYRFBEhSp6w8qqiVyOHFO1lMXUKjBEt6NaKqPRqnDMvV/QtREe5CY6HFqqRwS1Yf/brCL
0dFiERxgxXrm3uvE15PLqIMwk2dY56A2zEhVT77oBw2OQQTnpW7HDKTCuYFM0dttJw7JSyRWkZUE
2d2aiLOu8CMNi575x0Zjv9PHtrjgff/FGNAU3GirgWzL47rGi7Xe1VSKJye8h54uBKEQSCWflaUD
/ZhGAFvux0/SA9IKJeMdPOl9hKoNYejl3x5cfDbMqEOlGE5+9INHZ0m9zuAfz2jY5ZBw1u8qDtSw
mwY9jOQdRfRPIOy5ZXMB2cp/02pJaxUchufz0cEng+aWBddtc5hPzhR4g74pDlzJGXq2gR5nwhmf
NQZo5pk9SPZVsIaIyEQ/ldwfJrsZy9wWJyeKPQCNbxDTgw+NYiey+laPS7bV5CvL3jJ/admNK3lD
4k8IIbYTLmztEPR5Rkd4w8Wj3tRQYNaiiMioxJYTV7uBKTgj7zyTysm7t9uSnVldVGZHeXaYcf6+
N++9p29hALDFPmErXWwKZqHYwDnlhRTaTIIus3hgJGswZoK3KjY7QMv8Y/iCDJy9E1vvOEXOiKye
Jh38CnCn3aSPeTTO3pON6lVfV4V7H2m0iGrbVAnAz+4OJfApL3lveKm+Ej3Q725Dl9G9A+8ufVGJ
4yRMjDHkdbse+drWY2m3wALM+dcApFdkzFl4sBFoJv8yaP5XtUyQKVI+vysThnDW7vSZMuiXbn4k
UXfLG/TCWbByVEkWotfxAB2I8HMcouGXMWxU2PxAVtLpyn9EtzQKwpa+wFiI36cL+fowUGPEr3Mp
alg54enTNepgrpBGeiLEnDRPxe/W1g5K0tyXJ5wy/faFkS1Bn06JG8z1w8AvamIUFDGm2Cb+CxY4
TthkrwdyUqui2byBUyTKh5/NhbfL8PqHGbX2P1djuWjmbovya9XlTbiOdJlJZskG/Ti3D8BtaH75
v1Vr9hlnGVyFul+bq+/KE9CugAuOQuDZNW77BkwS2TSGkEOS2MuNPDwfdRzjxy//E95rARjYRwaB
a2/SjuqXS+gUNuYE34d6vkaRHCwjvm8cwTMYKPsHGYZB4IYeuFeZoS33FxTTDBP170w6yBdIgyme
QCukhZC4AKcfl2uPyneFt8FPbBER+ds5IFKT2/bak7KvWzqlnkw9fjz811AKg8wcNeJRho3VmGnR
wDD7mjdgixurryESp4dkE7z3ma6WQ5jjrpu2rvJkSgC4qHEDX+LynlTlziI7YYglk0GkGtSI6f1X
j++RqQ4wuAn8w7rP/U1fWvVZacn1PAqF7uaTSOjUF0JUGlQhrb9UksyRWO9csFuQhjqoL0B7qm0Z
hVsacUbMtxgTjBELmtEfngaKnmzkOtkIEvbTQrEh9X2C9+KCsw2NIlGpxdRDKcpwC84Eu9plUmNk
xoNi04BS36DL0HDfzEwMYSMfjKeshUQmu4DOKZHhQ4CJ48W/hdpWWu/Kvo7AJ4c0fUBKYubzosUH
skitBqrU69Smhm6P9osbCq1qqLCedOalxcI5/S0gBE0Zuj9x8GtS4nVXMJ2h1mXUAjVoVkrCIY6K
Vh6V2O+SRyLDbidzYtZkg/98rsdTwTUgUouOozZvmExw2NtRMoA/FQC/e+jYoCFYxC9/y0gQmUQL
ft4VEiAyzVRTPppX/BfAIU8V3iAS5Zl64W9bL9uJMYAnAR+BcUESnCAVRWfLaOB/GpZlIGEHIC7G
ZuLkgo3ycLza5m2DAdfcWaVgHugprnhifl1k9NwygMx2QzTTcsyKO4BWjDiEBQYAf+G8MM+VSR61
KqLAtKBTyNF0j8PV3eFzSvHbFw71WZoueqhPqe1tHLAeFD4cKtTgqURWgmegPxDyBwFTtBsr/H7O
iBCXVm+/SE9GYSg1Z+sQWPq85mKDq7rlPgxzNGwSBUwbu7mzt8ResBIAbRGxJ5AYkZ1WE7TMRH+n
asfX2WXn+nk6q1oeh9onj8gjiytd8bARM7XV/fUt5+W3UhRfXJCldEIepcflOcHzo1ZqISFDOIUA
ZAWO7uIVxRszF7S+gVsBycVcib90iFYxCtXtMPHJES5a2w6V3n3tJHfF7ac4Vi/8o9dGRY/FJbXb
/cesxIeUc2pXnQYVUkOkvm7SzVVMa/ev+MjP8ElIqSwNgVEekNyjffWGv1Fxt96w4uX/RNot0ZCZ
IE1/VD+GOIzilWYszJ6mzSctK21AofEFmmlMPEcA89ziyFCoUxA38xezvDXoO6wdVUHVAG7CwZWK
Mj0bHq3YrO1J3bA7GGm3lVs/O6DRzQFw5B7W3HijoJ4uSVHWjGKjCmPjw+hL+E/7r/gZP8odOzAG
xajOf12VbUQfgYn1MnmQiBfwodIa+G+0Ca4MyoCP7Ifzd60dhpYgdiBTrArQ0u1cGWiQK7DFk2ik
+eCAyNHGHhYedq8+5VD/tWZEcA0T8zZlilYpls7DKWoMpNQifhlTTBGDiz4DtditQ1jiHJrvyqeY
SE/YnzbgbTQhXf10lNpC0YbxSvOi7iiodQTEyfS0J76T37TveTLV4eoxatBWQ2dbZaqnjDia9bpc
Cu5fHnFvvKS98wDQJqi81Wd2tSVdaAkW5P1OjYL9lxoxmvR0JcvQDFDruSNAKFjiqTwbFoq6A3CU
v6137JkzyL2p/6In//qJMMxdXcsJpBJgwiu/wi+wu/MTT73edfn1/bOrz4Gx56E/rOtHykLjeXzz
WvC7mi20Z2a/NDBP4jq3ZJltBqKko4BoOO9LPtbED+n2nExeBtoUzbqO9zCWYPNuh8bF2qNI7Wcr
Cq3+qJMV/r9nM9cslAJO+AHG9F5HZPN5bqCPyrNhTkYJyk0OIhn44PO/0hZzQVfiSNTc24vcUSNZ
MlPCKa4GXtf+b4zomH1Wh12exXtJJnc8GGI0Xlbm6wTbOq82hsVe7Byp2WKvXu/xGyecj+bgztl3
Erc79aPT7WNiQaIAt3XZBBKXn7y6tkaQwnvxbtQwbwGBtTro0X7bLdUl9obsDA0YXtOlLCPAbOzb
YW7dSzUcTfXwv7gPLKU+GdT/swXiZdvhB6AX4nac4P4xxfH08W/YX1CuNzdF7bZWLXpq7Dtv4KSq
yHjBAGNZsjdEy9O8AJ/l+im03Ytn+Ch36n6e/4KOlJx3oCo6iDEHEJlA6p/7kSeogWLVN9VKcr2N
smqEtK6V1boSkbpX9Pb+mQRJ4t3DKTtzI1QjtoxTqc63lMyBrn1HglCw8eI4CkBxCGjngEzFOG5Y
WXxDV4wI6NufPXE6etjBrwLLW7DnFZ3JuuiMp9oylprNX0bKMbFHlKz3ebtWG77duA4LNSFVrSCW
U3MLr+KhQjGcD9RMl3+dvU/ix5cgoqnfPa3asmn/dOHkiX8Yc1dOw5LOCaZkCYT8kseMh8MiFvJ5
nsVCZwiUC/HcbPk5eNHB/2Uw6gSXFLiu1GKmVUjRhWkUwLE3hCozRkCX5iUwUxAV8v3iO4QVXtY/
78+zMErqWujhLm5PwijA7rS1drJMEH+S5IxqNBi+rVNgmvI3id9QwAZHfMmnq2uILxOuyPuPnDv5
my5rlL2g6/j5K9uDzd87U5Zgm6q6FS8KJLA+PczU9ZP0mu2th/yKZkwz1BlBIo2qM/5yGA6s59eD
oB7QfBChC5a3XU3eqxCjmEuX5ZJH2vx8XQf8puYybxxirgjXp37rO0/Bx5PKFVJOLGsfxebg62eT
zycxQ1hskj886Yf/TOZ323+z63JH9rpiX1lDDc809XnuUTMKfB8FihUZt4g74U+p7p+PEw6yn2/T
U+POGRp/1zDcyn0htjmCsQ27ijdPT45W9RG3DUgffXx2g+IN/vO6alPCiO5W4uPwSvqNY0pEYolD
BguNlo99LU9dq050/qzyXombOrlZkamNpDJuqEhTf2INzy7zutmooa6K1lHMWPdwhs3Ipw8ILicO
eQmMaxv7Xpi4L5uUGQSpYITostixlXXhWE+/cS0U6KK0YOgys1SvfgPWx71Qhdsf7zjnuf6PNOxO
aomH68Q58MbWMeE7IhPpIJWNNNguSg+At/iH9EsVsocu8G+SRJc5XGkAfY0bXyk3tyyg4Kgpuw4K
lMDJEkXTjihb7ARFnRfR/LzXIjUC+4sCX2ZbXoPSnH+NV2KYwtCrWWQrbRbZHhXbxL5M3S+4BEOJ
If6IRW9pNSi4s6m8n9jaXUf17u8gYEyPSFbE8bsHYFBbQvm8ynJfemhW3A8MdIy2/TdGk2Ehe0bq
nGoMzbBkVyW4UuADgkHYRdfB8T5uGu9ZPpyJVYYxeXt8EtSa1m1XXgYaSOS37EeN6yUpDUX1IRgA
YBPpt1fCEAp6fGud6QbbxZgUYULJOXQx7cwODIlMHen26O94NSwUBsvMd+Lj0QEE6Wq8w3f7Cn1n
Q3Sbq2pZJYYCe9IaqxKBW2SpTweQ04ZXI/AwB1fkqKuvIopEeiogQV4h23m3TU28VVc8X/N1SPbQ
ry3E6ND2sxv6Ygwjzjx9hJJti4NwXCqkuxs7H4EtXAommcpiB/nzFiRAwkoACBhH61hpNxY+zC4m
QK8qheXKjtAzY1JReBC+m17FE5ae7ITdDDqk25+nB2d3uDX52ObJNfFSCDe0B49YpVWYlNOw23sC
/rDzCNFrRbk2eePmt6XtZKB5MaVnMEi8gKJ9q0kNUQu6io1tZyNkRDZDn+xS1JpLMOvEDJ9J4zC+
LbevaS2jKpAU5ca+0O2yMHV8sHiqTrmvTnd7sy14+GLu4uJG92ZaVNCorMRFXWGubGrJEea+4IwA
IDlxIEgJReneXkHGiNZ4PZJEFkq8amiaKdWiuVkmuPEPQI8JGJD6zQhPIV26YhFhDECM+sn0YnGE
iCF/U8feajwwZjd+X4vPLAkj2VdY9EAaYlpTHe2WysvJcHCGU83vLXEZMBsWNQre7CRcViGIqZRP
A42hfwdm6ATZdPUg+ReZXxBeO7m0YXas//+t4VxQ+PeeCHwqzXOx2vdYsOjJvlCIiF0PuJacoOO1
BpuSgdl5dGRio/ST+m7B/jni7r0zr5VQK5aK7LmYTTVp4eD3NkhU3lHqHKsFPJyiKMobCJ0t5+CO
WWnE+S5Jkj447E5rlzuYk9UPd/aDrWHtkMIL9z3CnrrCRH2XtRZr/INcFySJfsnQBR4Vcl9cUTJA
Rnrd+sK0r7aJVLp0uxLBvFAs5WJEc2Echxd7xrVcisiT41E0J2N/u4up+BahtS4z+J66a3rzWTiB
sDNwVzaz6LF4wM7qQsJgIMgE/7liDOr9Z7ccPmEg0lThfIv/AXSb/veMs7PxKkLFXqdHG55CRDvc
++VX7VvGv+sDFBUyfxRT4QKWVpzNlRIy6yupgvX/hqjzFW6ev0QnQFf4dCcwFPAX5llDPszADlCV
ikFdn01iAiGs4bux6xZ0AGnquPxEphjJfVSw0ztvue0pLT/ggfVhBq19XYvKVZGuHIAzTKW+4VjG
UVnyCSXo1NvgtD2TXk/PgvVEMo7cMf8EaRV3sTSZOGv4M2OsipgIUqtxLKDsrFaTAlATowO1gxfv
sM4jS24Zvc6+2hF52DkVMU2UOikS1Bgx8sKj71ciRiz3lycBbxVA8rWgC+sulnE5sTVUYI+khpvu
9co18EJyda6aAj/hdeWXz+Rce7r64HwvySux5xdSJofOyhLyIcBfue4KJi9rKCrDYUWSqeAakiBS
zrmiuZekiPQfWhadP5LEKmBYv2aoQz45F5SaOnKoNvvnTG2j4fcB4KJfETtobtA04ybqkpnuvXXL
4UlnKOkby2wLRS/GKCt67Ax8TWyOAwMkUuFRBY8ZbckWDIYVWkCvQ1WeMG8zVLsxfghITePa1oNT
yhpjA+tj0jzspC04eIqsWajvhuYHjUTWmXjHbK36i33O8LAtyiXjRkuNe6uhHpO+m+C11P1aa+2T
VsKPmuysLt45T5Nx6lzVqu8+DJTDokPjrsuem6yLIPT37a7gB4jEE3D2rxbxK77uZePf29Kzboyd
mGFiMMXr3ubvRPtRW9ycvbneqAWVQD4Ti/eq/cu/1GMKRIoLRWBbbg8FSPynJ0JgQPUBCXLSCCv1
MFC7Nid9ku9pAFfgDrbg0R0UckOG7UEMumyVzVYgtObQp7D47VhTmw0Aix2+pb/a6wWPKVjNv6jA
5TwO2sjqKUeCLo3Wcwb1wkaQh4AT6WqvMpfSBb2e/PGqMyzI/or+9Tzp9reAW0l0KYrWeCNfXweu
/Ao5+ojgaWl2+0ODr200muuKsUXEy0RSdrRdSobbE21QttntpLi1Qvpg7nKTrBVQ+tnYOD6NMaV5
2ahbc+9xKJ3hYY8spDklhz9ZWuantuP2a5qkemEB7DYZq/WNZrnntKoR10nSuXVEEqcUgdSrdm05
edb3u9+DiZ5Z6IT6gFDaI2Clgu1dnVxDExBYSU6rzWfqP1vS5wwtLzJojFU8vwuQZuAP9cqR6iAU
KzJwZLpjtbwEwQJIVRTiuGDKhNxCNs2kHxhRb2fhPHIXwHbxHSCCDxnL5UuZum9UhJOgpvXWSJWd
R1WYSBgYlWQRoYX9SrYa7Fz3XflMt29WSG6QAYWBNn27GiavGDcp4CjQ4knozR7y5keaj0kPgp3s
W3V9PoqpQg+53MeWZkuHY2SLjyzuh8MMAJEYqvAom5FsKM/s8OksPPmwqaEfJEQdOL7eBONkz/at
q1BN74D2+OTqyzc5lBe4L9rvctOdqSWEj3GgcZTmHOJfXNP5IC7Yz9x1b0YWxIU3SJO8K+LY+Xnx
PlcZAWgTSF0KNKJI3m28jn1kAqEcJOBal4W1vPB3k4frkUBKjZw6ikWQeRPjicMtV/KMptGfFZWN
QwwVGB8lT4Nhds8bGyowmNnUAA7IAaUlxAIYZuhIw2TDvQTlYVe89beePu+/dWHcZvTvN+GTSGXo
ZZHfTOWx9IQ1kXvbPHeOlllDf7qZfrq8qgPsWZnh5cFMLlKil1yAyrOzl3Ckf3ZvCimyLdWG/FxL
e5H3gbZ+Ux7vnAmFbk6LhyDuogmo5T9nuIunXWlnxuTjsaUnvduLoh8dKMixlQ4wNbnnMS6K0r8W
Ld8T661Znz9t4t67m9NH9hyyW4Y7w3qFegIlgj5Sz36Ejqt8qt7csNNUPMY2rrYv9qrNOQrf/iSR
0H780agaJI9/UKZnOe7bJz/aBVbJb89w2kSOtcRE2BsGW4qtBUYm0S+xOYgcCl9mS/sclrx7qVFu
qZgjr9ims23RUZkIdkV5qTe3WGCQ7D5U2heYi0LI17q91HDSkVe+K00mJgZl3T4ZiSkYFyk71R2d
hBiysIu0oYFBYqm5tTRIbIajhmHb28/RoBEUHW8nK+CkCi65MjpqHBeI7fLV/rgmukIpjJ3xIcJZ
6fsDsK9UF138zgUDGAbtx+/3tBZMtnLGlu2Ulot6YSGE2JHxyuQqiYXzeckljinUf++3C7twArL2
8ncSb0Y3TN35O6iT5JEZctlw4PZi4wa0VPXKwsQiBQw8huRnsAwxMaaTu4T1aNzCP01o74E6ey2R
ZNz4EKJLt35eRWPEGP/Kg1P0dQY3+VGcX8Vz/jaYflEbljz7xw9L8GY3f6QM54gEDIIcQFM5c6FZ
aiLGGkz2BP8+JHboo86mt2Xvbt18ngDdXsvJl3D72KHRq95QTy26fyM4JXgaNSWzfNC4DLpbvgp+
qqgpWR2vbzIEpPMWlX+2mnl56ciT58aPfmam2QlFf0KeSAeLiLzxrJm2Jc241O3ItzE/UPnRMreN
xJ/4Xj4llrjj1BsCqN8DnHr73Wr0sLWoWUwpCPaytwbIWXA3by88vW0Qi6VgKo4KaD9QhMpUSJBS
dc1ZhUWWOtxDyUJRD7KvlUfpw1c8RIUdknGhbRpa/WtAlZEnfUtfeb8ofcBRnbTpmCv5/xqNuUPF
yaAO0PWRGwghanwD5cIS+2W2VSEEQAde32pG6REXbE0gzKfvwhVENsxNPYVOgolEKjigkEPT7nb7
ieX6/QjKFHpOXsN5htn7rNUUI8RDYR44kSI2tyRm1tj2gqC3yEy2un7V17risZsZO+gMZ4f+UYDb
4ZjkYRlpIrFuRV1Wj2vxYMm5bZoBjxh3heqCon2yvPoHN07z7JjqcuGIYuWDw7yRLiFtBkwy/3ET
P/bFrKPUP9FJdes3GOjcQiLSI2WOT2wXVIfZU1Hmmv8d/cnDh9khZH3GtZc6LwqUqfb7TgeEDVH/
Yc4ZBCjKvh9vipI3T7nV5MsuR8N8bM2tVfHo0A6FnWCX66gTA2C9apDd5zFK7Av4i8qV5N7N5OXY
0oYTNd9nV2UcEI//Ev997vLPBR0Jygz07Z0JpIRuhNXEjXjgCcEcghF+dpWhoImYcKsZbgC6+gAc
n75MvY+9HO7AlZyUBKawPpx+DiyeeS9To4nuCke1/kcdX/fCphHqW7aqHiUZRgEHSsp81cB32nVM
LA872fHWyAAQcOCxqD0Lm9IvkMBtyP3HWmjAzIzZGzH8U9h73HEpt7ZTBCSF0+faJjj6bXvPaPj0
On5SZP36ZPz/Kg33easeoRc3enxQpz+q1t+ZSLjgEWu1z7Zd/aft8fiVru8mehQp5ApRkP4bOrdU
ig1Y6nm4jVw2QBT4kPyCWTYNTTHvhSVBym9jSDJ6h2T1Y4yZCUtgTWV6LtOovtn9aqkIiLtQZl99
CH4X1yTY3wGJZMRO1hXalpImXXAhlBW48xmqD24pBJeyaleRhXb786Ql1V3e6TJ5jm7RoxJz2hTO
lfSKLrCfyBeadPAkr9vGoKy5BgjiGB9BQjeKTYwjN0GFkxN/skNCQLIhydcMjTkdTvO/dbFUbU1z
Y88rqI7Fhu6PL1OF1sUYlJPqHd/T5untx0TmjCX4HpKuwflNWlfiXIVjdUe7pyqxLI0bYw6HQOyX
PmVnUkcfOwZLgQWwf1PP+OkESZWr8LRIEpKvAsi5HgCjkKw0Qjt3ck+Yx42A7je8f0/7+69XU6n3
/RVOPlVfjRXD8V/GPkPHmYOnNhxU0q4y39DUfpaljsWE1WqlHUzqcKrGSsq2F1hju6u9zLMvBmY9
6X/QLGFoA3wKsP6/e4OCuzzQDz8eKsGMftVPrJsBcHCR1kcn4ePx7Zl8TrAvUSMjx+uwOeG+bLQr
IJUdflfBxDRYNUe5CjIIN7uVXUzK+4nQqM2XK1jLx+ozfdWAdMQK/YKxhWBifo5uH362t2NRW6Y+
HMvhW3M6MdvQI5PfIZlDTRxcTEEywXuXid1oy9Z3+37rZB9Q3pU/GeJEPqRPZR3zU76C4fLaBP05
QvZ1pPvFlLXj5CN8hEW19AotXeKGY3RunE3FPE/pzbwooEAoWkK0vPX9IVj22knSO9BSSRfMG7/o
5dPv6jAEyAHcVGz/KrEn8ykVZxf5IoeoZjxJye7jAyrf2ImDBAk7r0EGPF8eZAbLR/FXxL/Dsuuu
kSWlVDjINaAL8IP7j0d+ryuRaOj6qenMkDcV/85bu1/QEwgnbl8JmFByEFmJ7k09vpBfebRzEQoL
WPu1sExfvWDAkVuFaMOFiPl9glle64ZK6sHWVpRLETG+UExwyzB2LATUozXoZRgRz6J5mDzhtKKT
1UCvgffwjzPJg/Y08NmsBhSiyblDpzpIuy73ncRTLvZ7C69sknhWbdbwDjUlPY3Io4FG8XcxTM2W
Cb8+M9snuoGvNhL3Oxwcl4ShHwbSjzVnUMw6ZcRUoZTPnNpHy8yaOIpauPwelAyWLmBTBQoaZhgU
nFG6DNtUzoZ+4BgK6r4dMovRUcAL+QCMiTtxopFxqOxGk5mY9/cBZns1Ougze6Bz/kjPzDlyr+QD
sxJbdRp1dd/T7+Dyux3cdm+3xHTAC4CUkDQOCm+6dncCgKGA30ve0NleS6uil7KrFtFnJ9O86R/8
GvqWkIhVPkCHw7G9ohbvaoPluI3ZvoDryj9flng9kAnmpRS3Z7pHa/BenhkeqXsPxooQ0Y12Pi5y
6fEKiOOSKzwhAgqd82+YGW9wzxABD/RObbI1u2uBcg7FnmVinqvb5tkSBYTogD+8UKpk+pDhfD4E
N9nD2OfEIGvmtWCK+SrclotEiSanMDYb/qpF3e8CTLh8oNSDRpqgonY6qj98qfxt/6cbWVBezVxy
GqPVrli5jtDgzZjpdVOmzzJ67m6jf3OlCGvTKN04MdR0OGEId3+qy5TCNLdIt/iWAfX33YBI0MfP
PGyI0CGkb1vDFey9VdFtZMP3nzRUPCTjO4OvBVJkm98zwXV5juJEBBBqCz9h4MxFi1ZJqp/Lzzbd
Hu1nRkZoojcJlzjTr9XVQAOROQV8uu76mWvN5WMUI7WNgqAN6AFxNf0+eN6NSDu92xN2rboOK5qy
9HOSvIo+oN9EvIS4P4Ka8fKKHdwIRxidUh12D80soUx10ZYOWffBGETSBdM/IqKfYYCCA9O01tAf
a5THGou2eqEvWEddD6hxCTwuE8oFly+/1lyZfIwRgXErxvoiE9ERZDCN507pI7C5cJRw5rZlEI+J
OECi0rW+5KA8s8jANfmXFfTvJl6g+2HlE9pL7AzWSGYW9pBtmx7D70OBzjrJERDKgdaqS44vndRw
916e+Tt76w5vq5x/cpB84XAfJVMTBf4ER56ywEGtjBvDRHYMBMiJ/+8CC011i1Us2VRZ2aRZG/Ca
QNrx7bkhVStGI8zSvTZF0xP2WoPV67Q8kPxexOkMOULZ+O5qdE4tLBwaQXFxnasInmYOJApfGR31
cnYwsiyRnaNiQ5RYhcqCp65sY0CYTqgHlN85rjk3q4iNE8eyH+ZKTH1K+uwLQUR22JoxT/zC3B8W
nr+D17jExwjY18WTJvfAqtNeI8LcbKcFpBGtCQbuqs5WhgF5sMlwu4aPRb9lJHssYNusuascomBY
JfWkIYppAjFKCCpXvywgoKA6VrROwmxTzRRu5L+9GLqSr7a4G0Cdfr/QXe4tZfdA5BLBPRlwNpkv
jQeAzoPMG6HCbqqmLLCZqlRuEPOirma2TuNuq+SK6sPoDKmaLG/cAeV0eSJUWgJy3oZlFSxuuEoI
uT/HSwIqw0+w+JXJT7e+n/ekoNCAepWzdd3TmGdrnL1pOM8bO/qzvqXZGbfvlrcyB2TE+ZZtStYd
J1Dg2T6FzMTa0rodAQgURtI0cttejbluracUiQdZ2gLjAYs5SodOig/lu/+FFZYQrQj76ZhTAN52
nH4cw2WKKW8DsxHe49BbkF3HuyMT2FSQeUOXmRg3Hli9N35IQ0ff1FR72JvqCl6/m8JXQubFIHzG
Vcy3sYjkQ9gSerMEP3rMzTjDWhCMn24k3KXO3HIwIAiccaGYNzo258rYXlnuQN5QxFXLtEu1KkAH
aq4VRhwMzJKU+Et2eFdTW6AkMeN44NhGWM3oJR3kO3YOjdl3POYpRk2Kc2SGZ9084Um9fde7qr6b
ny7CVaUFDao+IdWwpJu/VLHgzzlmZyxYp6HUGzJiDnHT0qN5AvugJ5iyNyUBAKi3KkMbmkjBBZnc
i29uTubQ5cORYtUSPrVfAoES/PwVYxHvB5KLZ49xvllvORtCDCJYB50EvdgNtVKpxb8hQuxWHUnu
/rspKvWvdF1TDJvSh7EFOwAmoSfoNImkUjEYF42ezyh/+7Ldr4SjpYfDvLnWfIuy1yXWIyhZqcFD
n1TgxCJ3lKK8KEILCLyR+a/juw1xszhrn/7sIyUJPMrDPglHAmauqwOw4YRI4Tqn9hU2otwwfdDX
qD3bQ49cBXACVs6Da0ixCrcTISF4fE0NB8KaEQ1Cd7u/I/dpi0ckvrW3i80lZcr1gSANkczpfUGb
yfdyBHkf2gqMeF0W+v4wS5EmTFIMaNM30vh0oyx+inuEkVUFb3edHEESoZPSzQ5nzDvLTDJ2uLkG
QpsenQABLnj3/jUFKRKjFynGas1n0R6bxz3Taj91DOnxeL9RzWWUE39WgM46zTMvXnIJNuuvxYa3
VEusjdXIjp5MNPxLYrHF+FEaesUsIukeQCfIqidMnR2k4cOAPy/T7aMDL5MP88RR0qt02rdBOYwI
91lq5AWN/FIyamEIroDppISIlu9dJyNaLMQtdTxTNEsaRq1N3Li2Yod9BNwnebkoFePiH7mrfg88
N+2lcxdZfHXmEveZA9HMg0BReNn45oYlE2kN5+pFWbnBdjd5uJyX/zHCnu13u0WfKiLbGlLeHy4G
0CaBA0HuIqYnMz3XbwUFlPkmfek+hX9lCyRv7cbj4bPPKagaOoaot/7W9nsqjCi4eIVM0NQ1RI+U
wWykXyCfwIxy5xfOSLp/FiUjIaeSswIy9J2rZIUZ6Je2lBLiItInKhB/WzBu+UKOdSurpyVOx0Ga
ND1BHcJLm39iHH0Uj6BnHE4CWLyqYtqiTibnk1AfJI+ZfFWOnoDSboJrDDONRjp5eyvr5mMDkXVl
RUo1jAHF1RRn/eVXA/hUKoL2UjweYivvBJcZ7J3GGZ7Ju7UTUISc6GueqNQbUisc7omSu7Uv+VSp
ImsPmOM/oFq7ox3u3b7mfranKeUtRAAxXYmOcymMsCtIktnqtJSaBbAsxMpo2YcHfMYGZuwa2KzH
OPRMofMGxKn5CQUwwqW+qxXnjoRECLqnjEl3MjdH6VC7Q+D/um5VvN7zV1cLBIqXFhool96RGxB2
qIMlb8NNGnWzwGEPPZPHeysXLAYDQ9rPNu7I2qGP+o3X/43Yf4z4N+VYZjZ9ON1tUwtEuFoXdxI7
ZnT6jwkheNViA8lLnoiNElbJfkiu1XpfC2H+85L7EAGiNv8g1Qdu7mJxFPrmGGLAmwn48xoA+j1X
oYVsvDbo1g6sWxYikrPtqSh5BcEeHXRANb3iEoyBrrNbMXEwXsQb3GbPW4s33aaH5CK+inx3t8xF
K8iC/HTUMwtUV0QQf6KiHKv9g+C2keGpJtLE+l1ku6WlstPkWLw79UY/BZIjt61W378pLjKd92dh
smdo++fzvs3XVV7xdDW6XBeeQQIEfDn65dhUswkIyqCDEIhk5vTDlkmoJ6XgSPZFpxjfWGp9VKUq
Pkrjjlsj/Wg7YB5dcgb0NFQtieHRG65na9YW1YI9u+3x1rTqfqhVb/Xl2w3+ms27cd8dUwCq9lZX
q12OL1JUlK0UB6jvMDnKnlcKTZORqkB8rRrodbdSP4yR/d53H3N3BKBvWerkaklYDbFw566hP+CM
r+4Bkn7w8LkxstYrizZMYOcx5LiDdpOB9ZN25BOnkuJstOsvge8xlU9WWZKFiWMChNnvOKHWRoIO
+/8Tw37jEi0JIm+IKJko9ldLYYCvdxqFdLIsMNv1JCT2XofNn/6R/ui9UYwVF+eGMA39ZVO84JbL
vRkowpPjMQvPni5CuvuFeiWsmZm+niA+xqgALJBckE+rwfOVXoSPS0+YACP4wH3u39IcUuUM6Rwd
901moXm0oKpkT7DBSNf4LkLSoQBlKXhNEvL3Dt0metDwEbKISEOkxGoiTX1YsQQUt7keXmpq/+jE
HkAM/MHUtOTNCZOZi8EDj2c0pjElUTGNPIm+eZ7YHyenKAvUqtcWVPBrgO0XSNGGmC8wK/p/uYai
5xHEGjabjg7JeWVud3UwqTuyEnpiJBEXZml7+SUW0nftR+f9+HJbqpEmqEfEs7piq5BDecGyGkoK
6L8lZPp6QBqP+l3HvCmSERrxmxCrID4en0Ul5vviLtohEBEpWl49dqEzbdd5/dFPTk1ZfiNjk7Lb
1+EyOSOQuZ4v+1zKbLWLb4EYYethlHuNk48NbzYGOpirEYydhvOmc8zDI12LVqRrX9csoFHHJroB
7rOKWeFfcO3vYeqIDaoTZlZy/tvwUB2VxSnslvkf6kCrE/FeevZeKssi4K2SRJPF6/cxM/ROcIng
f80abDQ6oW2nuMPi4YpmkPLhK8w7K1Sp4ZaXPa1hfVk1o3xuywKeFg0uNUx9PtH7u5JpJ5X1wh8m
IoQHGfFx/g4+Zh+0z7qFbxoIEvbusEFTGTePqH0fszGb3GDaQzi45W9lt4g46sd14tkp9PSGtdCa
r0/5sko+DNWaYukSC9jzRAhoNOsCDnQ0ZnDZm5wYLOJrGVeE1wj0mKkGLN3k6tagMJjsQP37fk7z
MCUExL2xDqJNUo+9/PK3aBu1ZWCS5UXsAtWMvO2Qf8+gHGMS2tJEZlrUUDTjgXpt1mfHc4/abUvN
ZxzC48irgnX6Vdbjxp0eTsOtzHMRMDwl9UBjOcBU5lpTqTCgkEiux3vCIDBvzK+lUK+mXBBn7nY6
pIjiuiaXSBo2jbDdQJA/FzpMsjYpuAA7hKrtj6OfvRSYmmQBTUOWCoJSlqxdx1PWnKMf0UKPkREJ
dMbQJTb+j6UPf/elTqZxTAcczVrQAq01qpp2OlY093ZAdVtwQfMeECJ70gYkxiDKqGJnstGCpNeA
cTrBzJYzq+x6ru5PEAk1A7zpcvBJhABO894V/fgLsEjUQ2KNIiA79c+ZFaK5anCke+WvbjSXxySz
3Q1RnV3yU1qm8eWrxtQQBx7u+8rz2n+6m1/RAl1JMRpm5ITSxr0oYcSKw0DNR9f4mafGE5Iwxnqc
Wr3+lOft+1MWCvFTYDPEcnpgkXD8h0hbovfgAJ6Pj2KjbahqQSNqIBDHyyeMjZmmiFxRVYxt+zqO
BOzV4pOR8uItPqlADCi43y/mDMdHqblRzrVnZ9YN3py51PE2rM54AOiiRF9BOcG4gcGHuHq9E01K
EAv8/vbXmUZWUNjSF20OdzFuZpLTKaTzF/jAiQzzxreJOvkyVoqpGpJEX4LbekTN6+nJiv0lTyOd
RrYYPgy4zbuqWCCkkCfKa1sks1Pmj9JuR8Qs+0ljilPqLkS2H0DMbZJDolo+oRZqORQBlhtDgcdT
Gct6SuvXNSZIPzy4/DYoOFWwqrQKKJbSyiFGMFhMhxij7XuyRF0vT1USvPAoH21uTHFvH2Ja9QFT
N4cWtBqrGPqVemILZCgNB3jN+GE33ktpoqF8TYZAYwjNANFJfBlok2VUIleWWh/rbmqHYoxim31l
buMcbhf7DpPkEpMS77ENamiEiV/fA+Bf0PBVL5euvI2I71BuUz57OaGb8pA/f0dOhde2gbAaTNSP
L4nFRqbQATf9SFWgoRE541i8pEQrBBIElc7Ewe1+XUKfn4751NM1IGmtn1TJkNeFmNVzAq4FV+r/
RH+2k4mdPdY0GsOrPr56GBQa/vucTviGF0nSPCCfdWH4o9j/WK4R+TSHRTwAG9VCTMPlyttGIEQI
nARVqGWTgc+RakFjJ1DOBVmwT3AIdHShXDN25Vq5ZWxLrnotSlS3MutwnYqTQOXyYxI4CggdgxkT
H6ESki2CkfedsgkuZ5C5118e6hDOYWYigbN7Ji8kLLOoWAqdaO5I5ghYMrlJanmMxDZRjZ9YQU64
6GbGiOvMzen3l+X7OZ37DCjNWnrFIcFTI+/UgIm1Hy76/JE90rCMtKgjv+kQzir64SeRW0HvZbMd
Q273izf/sc/GXFpubU3S6369GEDeVlhlfTDt8vCya2dW+IygTEyNV6EZDXdBHB87GHTFq6DK0lwo
9H+GH+F8aMrHw0gfBvsX4kZi2NkzZo8RiDF29zKk1D2HY8F+/fd9DexhqLxxOZ3XwEGZSmwRssWx
pYH1EI3liHt73Dv9sNzC9vr8b6i8Bd0zk1T7EeQzx07vvm9JcTzhxCPL9M/JC1xtV4yf6IW6f95Q
Fdp9Q3nMw+C2zixM77N8tBSsc9Y48SYSoML2JzfCTQ5qy4A+EV1ch17UyN5YzmdKv4uq6QHNm4JY
sRVYDL4B+kjFLmu4lqxffRuBX4nOw5ay4ihuemfeJ872C/2dgq6tJiQvuyw8Fqw3KrgNYRbe1tqH
4x6JWoirue+f+2SAD4ECIjwGzuMNAKoEwjUDEqBMlLX7QE/TG79U0E9wKh4WT5oW6O3E0XF3Ujl3
nef3p3D5bTK4Ru1wks2+rxYFxOd3Qfjbhx7ZoQXZlBlWnZ10OgE1k1h1GqS8bt73S7gecZnyaTfb
fLzqf5Dy9ErN1lo0mL3n6huIukYYgYJmvtvFDNs3AtH8L8AGwuttxNZ0zSEbtBfaQb8qFn1LXjOH
IH5DoxVsHYLbaQEz2R6KdvsAWr3n5GcpdJpVGEMQRBMfUJr6cnH4l18oFVhexIgNKzXpNFDMPLos
lmIdSAh8RhXd8jR5vjhnErBGyCCvsr4g8V41Tkwlg1lnUc2LVfZ9auWkcD9pzx19F4CC/YS6KQ0+
2h8dScmXcpWxrAfh8/y+N/k7LfKBQUtMDxUISxpLk6EM/F00JFR3qrhRPlx/QcQ9B3HKNEKZQKVJ
pYZKzmvwQ0ciZOtKKYpBulfdU5xvmKJxQWNvP5bIj99puK61Wb87idhDiYacjK8XSzctg6L0NAp3
8Yno0CFoMQwhxiJGIr7q4rpGpUblkVOreIRMa0h7fih5uh3ybGqg765/ybjNFotvvsGO3WaQVbK2
F7nGBdo5fnZetWSFzbUnkk8YnpcdS5gxRQPFSDvq7hMb5hgB5XQraurO88x6Sd+AXhn062NtQ5fA
S+CDh+Hs9/XGpHRmvDimfGVDwaKplKnTdhiz/61tp6T2h7U0N8JVXswd1B/UMEcz277HWCBbCn7f
hSeN1hKLwcd9EogoPfzRhQfgeBHm0Pl5YBLQQqPpPU67gMnL7V8hwHQJdCCZMAj3Ay+XpFd4sTpu
kYqXx5XpCveNCwl6FwP6sqyLdzNrDB+FK56asLJPjb4IkZClJQcFPFvrj4jHwFWF1emgbnhlcLW+
B6TNeN8KSor82GI1kHB2WpkuWVzjpbdC93AyVxpvyvMAlQfIH/v0tzy9IZ3OSskKDkC6uQRm0riy
mIqwZMa9dv9ziFiwcvOHqQtZyRiJ1gB/5ic79pc/v5O969vWBRbJLOfckTDc4rBdYmu/tnt4ePPd
uKiSRvf5FTlCcWylcCa5aRov5ih29Q7csFd1v9SVSAvv7fKezqjXUcD3YD1vruBf9xzPjysk8Iur
m5iYpK/KrRIz3G0K0cuVC81IFLBPOs+xKSdOUSnvciL2s9IhhXpulkYe2VC56wY/2JJT5facxCB3
v96ow4ME+jHepeJLjyodu+tsdyhQKszU7sTr5RGAMxZd07isjvlim04JX0ne8TJlZQSe3YtwTFV/
6WNVm+R6J3EkabyxPF3S7naDuGTGcRCBuDD7qEVqotj7uk1qbdHmopZQVCMzwu6oL4kpPHQCgM8W
0xGm5voa2UDOoSKllvljX9hUw18KXOTkiUkdadFAbGeXCjyqBxsAkKGA8gZ/s16nDpYx0y4JE3N3
aBNEyg8ZF3e8+VSq8kR+JQ+V79Ct7hsGPuaS0eCpxDj65W5RZrVxcBzKP5t9OzDm2DarLtO1uiGC
m1whP6WZd6eHSlz29MTZrZUsKPBa5d7YUdsgHs10vL8Mucy3WhiOxYq3FI6SRDnyfSQrKNEyDvni
PNL7JihzNuLNqQwrycyWU0x9/jzwLTayev29Yaz6uiJyaY4RAOPlnE8fDY2baVmjC/K+Vr5f2wpN
7JXIVmo5A5eHVcVp1BcVNbaIjrajtu5saOQSaHzHq+g8xHZpwf4rV9I79Hn2AqNYTWLpZZQgOvWm
QXHS85CpX4DKIAK5Sr1KQ68frWt6COCRGKCWmBjQbfexiEyuErNrNMQdnshEsWRuPKOMYdiqpw2e
NWlksq/xl/Bgn6M1bN4Q2he/xcj5goJ8m8s8wN2Iy/UmP/P/Baq3P4Lsi3WOiK2DtFM8eMI39Bd8
wubIWlZYMou9pbFBW+RCYCq06xWsVLbb1cMzJqt78lwrOKjPCDgaIczAxZGmqSuRyyDzBbKof0y0
BZz/OU8Omak/qesFNCtbk+iVfFKPcpmjbliVnIN/lkYzcQ12bxRil4ddR2HD/qqAaRBEQIcMZcoA
yY16L6XvXcfGcVeG43OXAws05Q+iW1U0lAj+ih1k7qnNIcOgnaJlCZSbqipxMCDQGEx1WQbcwFQu
+kgzLUpfjl2wKcfEy4QDm3eq9moREtPLcSLrbE8UWqVjGf0KB7uWUS19FwDqvF+ZG0bD/YP0EqPi
3NktL37LKM9ytrBE58TWqHp1gpyR49W7FwSAp1nenmxIq4nMj5w1EdzgndAeQM5PyedMMdG3zW5S
AzBoDajJ76R7w4TGbgP6IDZUGlZgfnKv8FD3azajLtNMBUsIQbe2GyDBJH5Guf8hOUBtgoLf4QeJ
RrHi77FQsJk+M458MSJwEAoS1n7EHoQE4Hwuh83HByiS7w3WZ3VDNRTMWDrUV5Tj7BXb3x+Vyu0a
K0/uWHU0IzxOGA/oSsu52n0iFlyUGz6GIziiojtpBp0TGYRcT8WktSKQ/Zcrw4St5pSkWXae6oiJ
64wgp1To1FjgHcitalOjdfXznsXQi9JV/zSyKH5Y4RcXrfMJF8OGWqROP8i38+UqjlU1cCk9LNSc
VjWjo8iKhkXa3nUbrPFSDam0gxeeTtwLiNhKcQg1FFzdCA2mx95AJ6bDc3+fSlZFFqmbPUdAhi4D
VPwW+5XX4vaGTjaclkclOIKknK4lGXem+EP8IpgDMHgRN9jK+V3oxtCkZ1AGcz8NsNO0tXOXGdsh
vZ5SpYyGAJ2QDpSe+S44gEbqJJ0MmS9o6B0b58YyGiKs9kTYdtiW5zWWk0/bkletIuhbImGZjkIw
jQlXc4pBNB+fAD59i5FuteyOWN8vgYf6Qt4Fjuc+rdsDSNW5CD/M3pguEI+gvuMCwPO9FH7CMjAv
ZTv2j+gbwpoFht3CdK4vo4EzJqSoychVAoz9/iFjJTqU72pyssiFjxhfV97xFS36PjacS60qm19v
PcxLFWW8ERHLAfD29jtumCBIRGoew0cN0BUfmjaQ14OCz63GGwT8nLYuMBeu1p1zIguzOpn2WHo/
9epYVFBnWBc/w7wBGz3rNXS5O9rzUDTl5bzuTeeA+8R4jgoO8CfSgz7GZR345nPsI9m3cqYJQZtE
1SmlUckbw1XOJ5KVcl56KPjYvE0IL79c4ZLsDgpZ4srrT+OBm9wibJKx9siYhDhH7Ob43u1Tn3fh
hJ13gmgYcWJHFSkKfH9mBF6iQ74vkHeMsvEKDXbW+se0aPvF0In0mmuTfl7eX7TIzd0EslWcOxh1
KMPM5aPe9AgmMEcgpxtqO3CmDeNw6i2fouJTrlBKMti0xoQw0ohjEyhuo+iyJP7C0CeisCd/kul1
GvUu4KJJiKWsGQE96xbJ8ulAEQk5EMej75wMxtk74DUdM1uH2gFdJcWh2CPdpIbWOEicHVQ88PCz
2qEXvj9xZtXSXC7h4AJW2Ex0VCbpYS1/zfc3kucUpumJJTROWAHgZeKKEcKjYnuJzQ+kTAr+uoff
v6PJzOxelmouI72b7UgcVQHbXv92XfuHQmZPXHVAMZ2cF7aSj2mHct/gAkfoCNEDbApAzcDBMmwL
grmZ8KpcJvVLaA3Cp6oxiV95GO/L0RPdcMO8xQOJ7u0tytwnKvqk7ZFnMkkZHFRY4R9AYXBgjEI6
IHc3WQUz7dU+eI/2apl63OcVNfiR1rKV7DQh7/4EZ+C7oSoRA73bpOwt9lRA43/D6cw89IaVaDbQ
FN2KvaKH/wcapf+jI3i1N1Yz8z2Px4WzqS94hzkFUKVma7/FrcG/Z7K8bqjeAzeS9UI/30hzM1jK
O+O+s0R+4ZT1ORo0vZGVYUKUWhZ6IaMHmde8lqEDU9NF5hE9EGkZNkOf90Pb+tpS85WAycZXCgxI
AaiQ/tJy4mZUMbQCYv1jKTqzyfIOFWPlmMh/k/xsGAvhJctQbJeds7NVaUzRj7cYWT0HyfpkUdFW
G8KSk0ntS2okGWf8MYCP1ICSRXu1AjItOzUouUDa2MCcQru4TREm386zOY43d5XAbdzD8idncgbe
mgQHEgRJhhKhz3AqklU5uoRhvJHEnwU2/uRZxOYlFHduHl17hk7roWtl0RM+Ir7fTyNEpzCeaTwX
iUzt8aa5mEcnCL84HJaxwyvPLZbe7T8UeSnZElz7z38s4LBj2lZvKPacQi0Hd5dsBxO+bCoGIu5U
laF8bY9jfqJDIMbDUfG3a41VbRl33wLGjkItQdpU330W6w2zhYDggXKdH9SAAKXYP3Y9Z0yTEcNh
fcg8GcoC9MCrHLCyW0JBAUpSmO6FnrZoJKlLJCFCOLMPAG0czEH1c6V6p8lp6ODNDOSWlEeZJdSK
HF4SNoYaekDBQ8js7z7vt55f2XE1oZrdVrMs7vJuCbMNC+GW20MkmtyVq5l0yKZoz8V5J7GoULZm
BDwvI2IU9B3X+kQW+ECmgDnRq0yh7NTlDrPo5oLWjVXj2iimYYTtPMc506YqWrOMxcWyxLA/hkpy
rNw+8fhjgUgn0dP6Bz21fYLnKyaYsMFuxPiLVX135YOi7gsJQU5OZwmbIDKrDHHi9XJQquVPIZAr
15vB1QnfW4x4vtoyK+cjUncFxTUzF9vqWwtDV56h7WLzJfrmdAKxJAdMCocOjfcbkx0YZXkguu/a
AnasUP3CAvCszB4aUFwJIpapQ84pqDsrpMHF5UKCZIGsK4KdmAgJh2O0p3MAY5z84yuptq+VLjD4
GIIQ7QBWNJcy+4ZZlPqnvGO/sEmf0+3GZACoetYlqJzXvi4kS3Ht4PUp0ae0lIMTcWIkig4XjNaR
hX2QW9OstV+rwMkE+p/H9O5F/83T4vg4R3WPfMQ+xRWnG//pS51fO7cnOFmihgXE6jHh7a1D0EIL
GxbDpSPAZvd1boeJSzA4vF8yCyAC+qib2KCON8JLM1Z0HRk5s5CWDizmyuVOahl3ctoeyTcqaHwL
yDA83ilzEErfrFkXxmiatYz7vE70Ru1FV24NXFpTE8zZZFxFkyg2Uw1q5nd/u2Wz8dE5izxLFrOH
Q2g82Ko8bAQ0rdPHPd6R9sFKCE8ebr9c2uM62rIdq/Sar5jjT29O64Zv86RhkNkEJA/j3pv5ZV/v
wI1L/PKX+BcVLVaOJYfHDCn6PNJ73UMYIFueyfsAm0MyRWZOwfCuz3I+J6SoXY8/b9AildRH2qol
3gi36wuIJ7Zl66+zpTNKGOIg2pAZDFsQISO0BLarE6slphakvwXvTMpVqk8eGnFRkX7BrlnAGt6X
FcS+uWxIcbmS4y/Y128tTjvWEXiA1zYPkcpEVA8yvCXygfonsc/ro+w5TR8vJ1XYUAlkclTCIeAY
07D3DWIG+LLYcGHLmo0P2gXqkkJOp1IOTPcpZuXoq26cZ/1NNoq9E0ghSHdmvFZ4j+dvZ+19CfA3
nohYa81LX1b48qjuw5HGXFkaFnPdR3JT4gKsFtVQMFq5QeXfaOF5ostA3BBh/++Zq0jn0gqwMsUn
M4s75nlsj9Jv0JK+BxrUYzQQ0feHljGVhHVbgQewbrfAgr4tZV3MH9mtF6josZyG6thA6nIKiXY6
LN0t7bRz7EQhxelxu2pj0YXojaqlrHl90VVdR5p4vTwD14gR6xONrME8AlEh/ng1e36oAuMoGxtk
BNQmKeyf9Wc6WhCWRClRC3K10JBA7UXxOq/eaFY7XWL3Glw6kCduL2Psuhzwu4wjUJWe+HdTmbn/
JUcti0o5bJ3SOJ306aKxuv9vwVUP5vAjVN3acRVQT/HF1VtwET8n0vZQbAg0GR0QKXMXxINZ+Qnf
pGtOV0pA2Q8q0q9tBY07jwH7znau8CptMzdnWpT4f2b8+C/VqLIDLmlIpJR+e44QDgBikemBNKoA
UHAE8G94ntn2L83XhuIbcFLjpATLoRYpM079GWc3OUtzVCmeuajg5nKoE9q6rBnVmHHutRyhxdna
W1ZvHJgnA9So2JaSCnfUwqd53iM9XwxDV/bsO3haErpTui59AjUtDRL8dfB95hBBSDBVcK3wx8HB
ajZ2RBgmHwT2SLz96R4+4MMtBGc0z/6U7jHGsHmJTrZRtymJJ0doLRtNZ9m1a889py+6cFb7DAOu
iCAUa9JwQ9SC9KCJtUbO5rc8PIVKTvZAwyyWVDQdwjkE56hwvwIXOQX58PeWaWa9R7RT/6MB5/St
U33wjNWJOsC5/NkILbvOt0Fuzq+j3C5N3kedTmMdL2yEyLK6HJtkw3+O49PrcDfFbdd6D3Yg0847
/u/szwWvFxVaYbohmCpm6kFiimv1iFB99eTQETqWMG4LansoFY9G1fwDkT4MIPe2hxTT5uckGubN
dx2EoAEW/VMkVMMyLaQSqnJHu0DrCJ+ZCx0ijdJto8+lRgOgpIA9OXgnuAXRi+hpY5SM5NQhBtnl
/mGBUXimFVv44yeychmSROiTzzVVWmXGwRaJvz3JzLslQdZHvaw6raConugzsjEH92/OcUlCk/C4
Y5+bWKC3rB7fEwcRghDtx0d2YlbRI+CnH2opnfPJ4WNbNuBS2p0+yuVhvPAqpSN5neHkn6z0rZ3/
Q30JTWbDFCxQ669bgMYZ2HsR7WEezPB1t54G0Gyp50OL6Pj0O3ZcU+nER0jtOfqz7sT2yScy2aoe
sEFWzaSNj7ly9GRBvabARbe0SpXqdc8L4ZlP7U6EdcUQD0fKnyrQ1AJrbG7tLjsyUuWMqJAeuhds
CZ4vwnV/LhhCf5Y9qMeM+sEI6S/M0IrUARcyQXPxyeb/W+FfVRsTT30TUmpAcZBdB8/rr2Ha8O8Z
tk4JJ19s8DUqAMW378PT6haHd/uydQZAlx0Fzf2YZV3afzmU3jzCymKKT1KH5TdCpJsETzmD1JO7
5uDyPYeCsKfboAqsW7cf+igZVJ2nxPmRBfwNFh9WNoQzB35R8CU7lWosmDxi6C+eqgnpek57G5t1
9HJ/wl3lRtDw2558ZD3yGqT70FqOttAGfT2uK0PJo9w/gTWwFHLFS0eMZcXh53/2uzk/SpYiUDMD
G0OnWWqFyXo4T08B2KCRuJDRb5f7Jqpu4arOv+fyq+7qkbx/OZlDpA0nm+nWGwfpz5VIAHTqLS/7
1tGHz8kdolG1H0CSgyRONjkOh2mlmaddBKCuB9N1hvN/neyiP+L0EUePye73UT6YRu0c5eVWdtvM
zBXGlT6MrVChkHZeUMt4w5s4maL9eZEpao2dN+JDBDl4mNx6doboh781J25fWkoB4011HxVopmE9
xHI/cM41FjVdzRA+SwX8xaCGapjKvm7HuwFydnjuMSuX5ptE5mwdAuUOatEOF1Cn6annr7Sox70G
UFJc+J7wqES+JLQPG3ByYmg8QoSLl7gb/RCjNRuahmImx09XBJG3mT/J5gVdC5MCiR5gHAatCOQm
fytcRGSnkbrKtkjGxcxcP6RDjuYIWQ2tS/ZPbzo8m+VSeR9ZhFomq/0QzOD7RFmH9s15CLkyRqyA
zAPelauwURzKl1RLBVIUSS6WiSKiCtnKqcGBEhFX/PrWzl5omBnnzNcAjCDQd39ZVpwNISYa84zT
+dVnyN55mPO8ncHh0HietsM63rQDjxlqjv1+3E52mJNy9smQvUFzgHMsxv2SKMGLSjY9nIadYsS3
19PUt+zUeZDgmr5mX2vk/6HrDgTziJQ/GmuaYJoqLVJo/npnlpsh6NLiQ3ddGT8ALC09NTt64mQy
oVGUzr3q8WGX4GARS+3oLkxOS1IPQ0v6tIwLIckQHduyTOrmSVkC3Q2RXoAz3G7L+yDxK7hF0hK1
GpfBOc/bhiITlPzlonojKtqXURDIWWBq4uBwh22UGKCw8e+eJ1Oz5ZR7dXY4Iy8w56CNETjnYoW0
tbTUnRhKCCaLs8KHCIzJBKccJXb/K3NsuimIiv6WhVVYzKr+P4x60ZeTPkuCYqQxGYIywTPDbga5
qskk4xn+nFw1PAyHqklchFbWHjhA0amojZWIXdWOOP0a20mxOmejKhjW+c3ZS6sRK58//c/et3ph
NPO6i5Uq5Xp4iBs+rgER/iHAuqkQUUqczSrLl+PS53kBRJxqAvUiUMcFp9Ettj8CEMcTYPY4QHRF
k4JfqPlTp+3vSNYQVm1jvKY3SGanACulOCWUHBIhkjNFTPgBNLjBq9xrVKjFmASjvKPr6Y3kGRIT
qtjB8jBBATqvFcXybQQfhfKoj2W6tB7rPQNdXF9kSrIathTOedBTEcaik0qaYZ7/E6ps7XfQsNMc
m4bE4CQn0OrOe5hPaxoXq/NZoIItxA66hOgGR2SULfKxsYY18N+JJ3g76BPUSyKdQYNZHo5ekZlq
Uop0dUZrrPV+X1FeLkaP93ExqDWlfAI1cyv9/hpyVXSKDKarZuj2L15KH1FBl/BtWClPhXRCmsY8
t/yNWpAP3AtuTsF6IGeVgtwvOaIi2MwSuKPy+aYd7QJZbkdn/6dHF6yvYUekSdLgPenOb1LnTxLM
mmRu5tootZkCTsTUKM7JlfRDzjBQF/n2y0cHmcEbCKITWPlu8z87fVs95KYa9c2xVTWGNxnHo96l
ic/YPeWBOVoeV+k09KOqIfrdoUMZ/mk3dxpFZiHtnOO5li1pl72s+HGkY97LaXWDS/W4R3g+TbwO
C9teIZIWdhN0TRYoDLbBue/3EUvCV7AmfeV1AkIbHdhJw8ElfeFYpfGoVchwIB02ncwwoy1QzKuH
o914wB8UNr1/dsrm6TnUlrOXJQSYmFMo4tsgu8RBkxRdRUNpTbhpM+tY9BNaS5sEocEKnRVnHd0/
aU7Zji346oHsM1uYILsaMsPE46hp/ldUD6eNCRbNCapn76G/6+1I8x2bpWvNjVWhNw3uV4ufTpe8
BiepOVARhQRh65v+PTw3ove/cntgQerAPSqIms2SWzpXIMRYViA13WYMDj5XMXJ1R0rimOP5pe+h
WLuMwfy0XzrYspAIEGUxLOSl5dFOjXkaxWgMyKC/xCoH1inAFkNx+8hdnMJbI7b9BI62TLMdyxPS
qTK1+1AgtNxSt+PR6fGKLiBeEJuJyuMl7WYUMm85bOcvY0r9mblbGnt+ag97l6ZDMzZQQ+a2oAeB
rQx91pzO27/8tX1GfFIN2nxHpePqCL0fLhf3IiOmFv45fRCCLgCcQr3zY7NZcAFZQVnP29AeLa6q
nUNphkXj3DnNIVo4+/WP7cJK75U4+fMQ8oHLaTL9Qqt7pv0K8Gj5Vo+2blaTco8ermtlX9Z/EEi1
fuY0QsrqJZKGpBEX+Zw7aC2MKHpoAurbEQmyJPr3IW+SpfjYa117l48Ennyam2Uo8wsG1xKc7bTu
0+Wwn1yj5TKH3Rs9gg4XA90i2R7SzrQb7IAMwqTtXrUYQHDjc+FP+p94a+ZksnWZbFs8UkK8jIRE
EBSa0ilzOuKYxVjq/tyA7c4WmqD/qXdKauuQEXj4ney+SLVW62TojA1OuCVuel2EPOjXM6FgMRdP
5OzvXnFkoJGgERFdsakCFXIYai/uUCSF+zz9G+MboMfZxuvx7JCUFc1kElqiw5n+lMEgHlAcnkvQ
RGseAdGT1awpRSpHQ7Diw6bLb1AA4WlHZPNi/hnkStLSKKKw5JmKNTSMhNOuJp7o4g8CkLmHKJsd
8WGmltGOjdqkoC7Z5ZahQ72k/r9xu5MSbP589t2nnBExdP6E/JUBO8ClvJY0ykYzjVZ7Jm2vlxTh
OtyesiTlQWJC8kg9kc76Yp2KJN9YIsnjN5NCB4QlyYu20qC//zVMM9dKa4lxQzT+uMcp8NSzMYkt
kzOAvhdUIfeBqvGvgIVHuX1PP9kvR8S/p1KVMy5VwPFpfHjSUMd+j9HpZizt/LOmiWPcoHioXPWc
qt+eZQiKJxYeKyobshrH088lydtiqkluPvbEe7K3Mi6OL91uQKvTOFdO3o6hVCNMimXAPKUEhvhf
7ljD7xcsY1SPo5Fs5E8Z4bUGldp693eYi54awcmZNaLE8wy94UbEP7aMY6/w6BAy/tXN2e3IGZhV
lmCx/d6I2qL3p/i3j4zY48vL/eE6az/IAHhOSzJ77RuZGCG3Ac/m8x0Db/pqpdy8zJAecI+zExIS
n+W3Jzgg5vtIeiaQdzlJ7Rj8kTn0rZ5elLheljh+Q0Oo5XfUDz/vh9bNiza9ZYvMZHwfngU+1eCk
Ifve/MedHtDjczBqVb3tQlEQTs+3nUZC2HzKjFh8oD2h5/e4vKK6KQL/314j2/12cgP/qczS/1yP
HfwLEuZwVIwgD/P6H1rB+jxxfuj7w+J/Rb9slHbbJA1ro8fbzzq0atDLlpf/Y6MVEZusibYNG0Ip
0NYWJMF1/ge6JeoRQC4sx+Qr2JC1R4NoBOWe5B5G46pefN8FvHhVCczSxredTRmlyO92WxyuIfm8
2obRm1BxBmRlWdM+GpGqR4zQkzGoj281IYVDKln0dBmdN2QWr78EIhXFd5Z7m1G3yOPnz4TNZAuv
kNHM51cQBMc0dRtav63flUl/YjOn/3G8t1rX6SmWZpU7UdPvQKDufOcyM2a6oJ50gw1VRIJinOTh
b0TGd4B1TVPzReXPGTljKcgxles8EnAxVR95H4hKXnVByZWW0K71rFU8u+SxYZmD6JN4ygPryO/w
EvD63a9rHPLsr49QLBTXVgeLJyW549NO7bvcpyyAZb+V7LKYNqUrCpe9so+MiZxFBkgB84fsWnsf
/SaVxv6rxV1/uexFoyshyjxYr2BMDHV4XsAV7B0Pfm56LEPnBZlWiomurMBkeutA4ek8BLoF3Ib9
l2Nj7qWkNHDRH+p+7IgDhME7Y7bh1AkQ781b95yhnWUHcLtxFRo25RXrCJyUfIhY0hJyCMuco6sL
WH1KSpMgCosTo+GOUK1q/JxjWLnxLoVQ1EfZcvBWuHhbJF46yr/gNwMPY8KcV3TguKj9aI33XFhU
5UpAv1dZ8yoWgke5rojPOMxTeWxSntBx7vDhv986+HrnVvN9mFJsGA42haDBKf64A+i+wnZqEK4Z
J8ZcPpjjxnOApFeEdpLS7yADlYkwk3a21fauuqK1u+UMTXglKhJjHKmC9twneY256J0/tDbq0Aa5
xucB14K9ZngTvaVr0ZHuQcsfkFfRTITCdJYLNe+qno0TkO9fCPa+pYuDa2zupwDD0tWXSQflGFbG
1FQ4DnKPNVmXwH3GMKOvIdGqVb6JyMChTOInFBOjDwwanPOB0BD4g8bFd03MiOaQpu3QOMuTkzH+
runqfCCageo4jGpjSRNvJ98wIQODnkPmxOzkFFZs4BzIWFyuuvxaasK/uUIjrlt6vKfXQcQHgHd2
2cqVrG32nVm3kK4WUqugGDA3VTko97vNvr6plcYIVK2U8PCrXZosSKPfEyq8yWecy6M24HXnzc4K
q4Cv/HXmraqc6VGV7857InXU7psjbQBDwEEW9rmB9DP02XJ6B0CZRU8HuR7J08ircrY9Lq4axyPS
IBovdhIbzPtNXfO70U6+TepuiVnwpbbiMqWRk6f80tnVddW9Zzathw5NQyq3Pojh5GRq81GsDnHL
/JV3M9OkiZlfAZPQe6Yx/CXeMYDVDNp5Iq/U1PTH41PKgOW8t4kEFuLvviznntQc9SwiLTk1MuV1
puKeCShXavPrTRSzvldS5vrCf7ZYnRKUl/G1EDljrzGBOtiJJddDSATdKFuWtL9H3Wc3pLaGUi7s
mfPWZsEKv8+0qkdwGIc/dzD6XXF7FwdIBk9PVKXvVtAeVxndv/AkX/D1zhDu5kX/6TeqHwNF/Dtq
mM40ARtKwbGYjZWjR3xqqB1lVJe0VMKAnG00EVHuneN6oi742xdNKL6NOGkCtwfPN1x6nx4KPBEV
jqcPE8mnNGUO5v/JEOt2hvQ2JHr9b4HdPTmKOhudIwXeBzvuvzQyCvzm3MdVmIZ+h3EIm7CUK6H9
XmvKh6W9SF9SlZKsPhA3WTwu1zqZJjWFrFXsCjcfrD4HU8fFna7shYXjOlgW6K4agnhZsbmVQzTF
4jWrLjJC+Ww4gyna1GfIwLSdOmLJzlquOEVTEJUaTGG31SGtidwSKZtwuX6q789D+g8CG7rRapYG
lf731d8TZABPmFCGaqrSB0gLKiaB58NwMIxeLmUgJs3zRS4v7Pa2hA+uJTDyEC55nnmctoFXgKtf
AqZ/rf6oztc2Ggwf0I3ISyitSUM0N73pI/IJKB9VForQ0sP6+eqCmMqmG07TERmShwEtW7GlxgMr
xTiV2PoHOHMjgh1d1RmCKFxlJfkpbSY0IHHB/ZPDRPfgQZpj200xoBQa5FSB6XlIJutHfMzi53/c
+ArQYGqWgHcAOhvUs7TEcFAjnH0ZFenlVLL7G1FP6JRgrgwt6fjeTR6jwDx0yrNQ+KoP34Wka+5l
T3fgXF6Gr31N8jpBaTrhet+JapRvP/qT4FRffb0xc7yPHC3EWkglQFR/WHx8qghO2KTejuLH21wh
aDw5n9CGrehuC0qsZ4aws4jaLu9H72sOna8ij/UQwBozMj621iqvtJvZ2IDwXT6hY9nF621iSK+G
eqaVK5AMzEI+YpgzZGTmGveK4/7WyffUkYlFRyzoEgaopDbzXy9soEjt9Kku5b2+ZnkbMdzxJfdC
vbzkBL/+AkZrtPRH+eT1dT0poJTUKiJ9vIgy+q24u1yoHvGfZs+78dwiukPfLXQsa8xXC0hH0e9g
rAR9mXHIpkoD7ohxHaYnrIe+CY2jnXb1KNFhbBNR178CIozp1sRHd82qbSFdq2Jx5CEiOdsp2b2T
Rkhm/JQvK7LCtkkJqT6Rd/XkIjnnPFfKS2qcA4DUIWzJPtxFLhg6ZRXDwWbV0mFKPYE1skaNVtTF
RigxHgyX9D4p/tkLPkxhEpd3XaveKEgkFpyYPpx/pazKUXN3AZdDcXUD1jKXV84Tl1bZjeUgTSdT
KspZt3EbUPhGUb/eGyZ9LILCSOZrEzkn4zobr75c9tgzzsEqu1jw/NmeBBQ6P+A6yxXDyO5Foym0
Z2LDwgX26zzBhF3QC75BZ92qBFDnIHMKRn91iv+r38pJ7l7n+VUKNo63H8j0r+bUP42SJkq/UVDj
Q8X6zp2p5OwhoPj5zzAUoee3VNIASo0a2NvudaT7sUrwHUVahfUfPfurnlHLMZ8s0RMLr7P3uLMB
n5bja5prs0ujhsmwppa6remZZg/itPhjC/9AoRA8sqNaDjEQm/brX08ER2Pa+6lFUgDj6208Of1X
fLk+Lbxb9/WcxkGilCNJW0hByT6G8k1Uwj+PnIv0Yt9NiUPVhG1FTSFPSFH/s0ATIYYYjXrErqVU
2T3dThar/+y3ZWCPR0Q9Z1ZjR5C1I+5WUB+QgC7o+GOJMCDWXKrwF8A9NG2cFjuwzwmGbmPrK3fY
BwKZdHAg915657iraGQyGew2720uMxTDXyWhAA430qJTMYUVHUyrhMGJ1AlHVrD0c2lsek+ipnU3
76egaa8JSpX3KYqSGqqSUQt2dRP4gm/+4zEFYgDTayoW6D5rkR2njut8IP6onTjy//x4MSaafWve
AQev4cX0jCY5NJ3C+cUon/UHXh8v0VUxIMhgYPRSrP1lGnGAoxC428BwTHm0YvVENYuFEcYDbg+0
t8LhvRXisZltMG8xibRwq4Yqntzmsmp6zEZGCxyi4Y+sRzqZ1MRlmvakOkkSa/INCSWaHtEbpRng
/3Tuh8yGBjx98nAvCaQ+DehZ3q9BTgVEmeqX3ZOJivgcpWRWQSDveg0xpKrEB0pdoSgIq9ZPa3+4
rI3JqI8MaaQATPmiVT9VWApYJWzNUhpChIVz9inGBJft0zE1sG2kqA0EQZWg+7iAkiKhJxQsYFOo
TSocIRVlZSsgCJ+AsXzjYdMaqIwuKTaGY3r7EU2TkTICdzcYgqZiPLpMYGhoX6ly/sM3VGIjl2zG
ql0NvplrvEwixWVtS5gkP+4fWNraeOW0Cz3krY7d6G2Wl5Ybz547KE6wRFRPCZ5hn1YwckmLLNSQ
eeCoR9W66kYY+DSBUIu+b2QQJGNN4/p7BFVjQLnxI3Aeg/we2b7ElRoyMc7chExTDBQLV4Tds5yC
UCloImnocncIRyinyeuhI7XAYTZIejjJT1RcsXrhc8yxAtx2pGQ8ohqXOMxgPjfN3Tcd5KuVtiaO
P7gH8koSxeoMijoJowmIdeQ1ksZ0lUpzNpBEfW9DNn6B5P0aj9GlcdoDXlHojisssfrXWA+64fkc
O7APpKLqK/1MK7dPS5RfkLCQRvYF2VZ5cCt7P+057zvYii6yS83MYP+18gPCvaH9OnnHyvhEtJe1
jXdoMP5EulSBSoRVnTrWkwgUjRMzJgbKTC/A574dRKg0JlqeQMxhZnyzQDRS/YgLBH14Bg3ykFTt
QH1o3auLRue631A2j1wX0WiKPr3fRum3+B67zD1UQT8X/1KcvULbOgpkfwMzOvj6lg00OuSioZRj
N3EWfXA2I6lkF+FjLn49J0JjNJ3K4i1PcjTuC1SwnBZ/cPAmwjRgpYdXbmJ6DECH7mwzDIDIXxLM
t72dXe8RWrP7IvqlAUKGGqtczsj+FdHHhy7EQv1hMU+2Vw7FKCAPUQur5U63I6ynJcPDyvK+orY8
YYCBymmTP9cSH3YmvyIhWYa59whXbpFTLYHltrwFleZELx1x9nAhxMYio1/wa/Va45G1qPrQYW63
17v3vZYUoWpBv00Yp3Zomv10Pi7en11Ku9L2yFF2Mb9hbO5S97R5NnqdZJXQ7GvJqf7KOWSj0S1F
EswR57e38/WQjWc2QcHZ4Hk8XhuY+7NX1AbT86TG7Q+8MYMzilk962f6fjfWExGkoRa/GXeGUsqO
toxOg8NrAYL4NjtedM1w6yX74pwbgZb+jQzTkSsxYoHw370ccPwraTl/DFgozvrwe6E51fSfsHGu
0U239us4S9cvSKJZniR85w7/JTbn7bJt3upD9hVOjnOKK0CaC343C9vrZbqf2wXGedDZIYOe/KEt
sidOMB5YiUORY1hRckvzODeaqP2boe1TYbItTXad0rXLtgZ4iEUBt/fbWttQmZ3rr6gucP0f0s4/
vcr8gVHQ3Yhe421rnOjJNDfU8MK4lC/k8ZlDK7W+XyQhATMOEW+wZpgPODC3WDlmtNTLnedbGWqc
5jZXCDNYLwQhWiVWGx1JkBSqap63GCSDS5lgPE+Anq52vL8lVxX/IRlMAZhOTEVCF2vpQ3ecZy+G
7T2GQzfxH8IIqgaUJ3Fvmn3uSdVgfC9yrdAV3Ca/kl2RlGR2PVY6CWvTU1V4UYuOlieQIKcC5Zuy
uU9+0LTHIFMtnjrv1EarKidfYRVivfeCqlH/Bcnqhyn+eTIvWPZgbhIcvNu1KMWBqlBizJV49bWs
lanNhcf1dZOwcP5864xKRu/PXx2nO13l2PUH3Xo/9VW9m3i6c132u21fHLHCRKmQV1n+PsFUq2hT
7DBrLtccp5ZRPSQrvp3AEumbc4Gwd/g9XdgfejuUDjPEVKS9ZO1sq++OG5X1CaouJLuUzLmozCFx
gCHOuWXndmn9+bntPKXdkuPYBQUiIqoDf/O8CGgWyhblTNZDrDiiKH/mdVUBOUPFbjxyP5cI4YdB
LlQTgQG8fyz0WvfIIt9biSPfHeFY/DpWz+zCNQFwMLKgoDA0vpPwST1bLjtjJ1Dla/9Dt1GNAzT6
q2EC6xCgf/sbeUwdpK6M7mNTrKEXuyNkrI/L3Y66tlCvsG5kYVBrhhL5AfZ0qVVWXZCJ1V1Ycgi3
w5ydrkEV+vt48KUcWujFgMPcTYLX4Z6CMIr3sLFExzXo9nW7r16aUBVDVveN5d2W82eODMn7DphC
e22TdLUu5dBcTiD2CaTeTRcZbqIV+EUWB4zLj2xSP7KxLIyZXmsO+udbtzhVGvdLOQFUZfNrHl7J
iS8BGXpLrLkn+DedviDzpklny7lLzXejFfwTbH2RX1+mbqp1MRHRo6761VIXjrJQOISsqBqUxYNF
aEbXe4ilpzFl0E05IM/TbJ8lUiftufqmC+zNNDn/ePlqu8uNdeC+IXVI7Z+YP6WBicHe3JLPxZNG
rMQzKYNfPJJMV8TjHLHiLVeMt9Te4vDuOj1zl64dAdHXiQ8YwjxAFRM3ulp/H1I6wYiztaNnU/um
RHZKP6YDkJh+eh85hZdldJvNV/XnAzlvu+WSv6xUuG+e7l+Kr20vZMxeREVxt/lhPjAkdDuIxlcg
EIKwmv/tnM+xhyti4xaQ6kehJQfsxkBfjTHHAYbtRBrpGHth/uD9iKnlNFrMOlDrhHKHvXRWS0VC
5CYzB1U5R5OSzpNz2o9Vr1GheeTVC/O87/BUFJ7FU3d+roTdZ/So8ayZApEYUWTR2FQ0o4MMrX3H
BJjJ4L2ICwm+4YMRoVSZz8Yni64mCTjGut4GA4c18Q+or6hb74Oaez7vU74cGRUHpdl3pvuP7A2u
dGmjh2enCkfv9FUWVrXTvYbPmDtPbqdH0HQ292YalT2SS7DlNw4AANjbYBxn47ls+wD64wqFEtyA
SddGA7P4PAMPAGbZsK4EIhlLWGc8deJfmRHto2IuDq5XYK6MrUoVGxC/LpTZ1VflHdoeGp64/wn7
GtIq7vOwo+abfI+RnNKgalAcpu66MFlXYZ6CafcPC7qofDY6r2JD+RWcJGgNvICmbZbyos9MyB1J
8dsUL1mcOPoVjpCGjhEa9TVaBnh8SZo0PJab1y2mHj/o7Z0nxnHn1vGusa48EieGm7M5hIT3HWY6
Mo3Maetf6/pWR3swpdyrezi8qNBFQszbP+6sO/YtS6PVpIIe3p1fBA8PqmxwlHs/MsPKODH+PK47
uVe41KF1Xc9h/+RqeQjiG4RqQ7tcvJzR3XaMfcbvlbkxFHoyIZdw244+hIa1gkEz+iX1WbGMdRhJ
KCer07kEFoF8ZHmncfEGNztHAHkToxB7qTsE2N8M8AEEdm+f+NsJgLqep+bVTs85vrPOqyrfD1Fr
NR/oH6EjeuGbbCEVBb3Kg4ZF0+BLZ6PAG9seWmWLlriOP5CnH0q9WB7txMgX1nV3pr93nH7MeV/k
P/wsvniAfsLonzwEIWZhJ4wKTNCXyj1nBjrgT4Clwoj1kDQzuBbREsT90Ao3ADW3fcs2Xl2xIS6y
kjZKJEmvoudjX91WCXwlW+/9TTOwT0DyJJoaZogglncLmXPClgf7NXKaoBZLiQ9ZuLdddVklSSOv
GmvxJnq5Qlnkq1B2km2jVFKk90boa73s5vn4VADbsa61s+WE97duCCI0YSW/JDq6VrIhcHZ2ILiN
smC4tdMEn0YBYRy56PvD5/eBn9ron2mbo6fVQRzTajFy836TcrnnraOC0y+BF8tY5k5VDQPvb5lJ
rvCQpbXZ2nIgltT0c8giJhAjZgSjOK9PQs/xJFlkmzwlyru9A7Rd9sFFYwFcL6amWGvuMrWkj557
Ma17yYB+UK4yiV6kOWOfn6SnxHejLqyZe/aIH/5KoWM9EeFjnWuekQ5PMzCQm4oavH3nJ7Vm7KIu
2/7s3USwLSCOMFTlTA1Z1yoqWB9y3T9dky0nISzbzLGGj5TN6Yt9q9cuOO/DVXUDNHlRpRiiT7mW
jb0ZLovD72dL6HHEFUhjq+8vqG+5uxy33AT5hKfZdfxk/fqFPKcWVkGGPFjN7JMGhUoe9WbzNLL4
uPRE8swLhmuEH2ikG8pJhFDo0ZhJV0aJYRxTpHDQmc+Te/Z2CB3L+lMumuI4Awjqtk6vDJ93r6R2
UPOaZwRw11yc+C6ASyd9kpmJUMghLHVsYNZeack4QDGPnLDAmh+FPetmyamL9uo7WCQ6/kU+/UG2
i1HE2NuZWR06uOWqWtWCCP4rchMy8T2NwmBU1XR2hmx/ygODf/jOGsjT4ugrg4tj7Ub/UbiMZokH
NIBuvFZmggiTwF0n4cSfP/FhL8bzC84RS8e32wr7F6j4S6rxQYpxc8LZrbMXZqS6FniCPb7FRhK8
hmCOGJeutpiiQIQf0tcJENzgf9HrWExQijNs21oBTkj99hVmfgKs0MwmYTQFvQ4DAfnhAVJe4/Lc
5BNkyTHtjPPOzLs6LiP4PKsmwczKypzkprTQMEmVSdpjge2w3MoUccVyDEjg7ho0rashJciE9R1z
8DZVo24NIScVlH484fBT2PWUK8VfNSHCgnFQcuMKmMYiCjWB68R809tDmK7qSfkE81R2HW88PLj5
G3/3nepVyG4QxIhDxakrGC7xgYHsX+kQwlySeG15AAHOqGNqr4AgmKZPFfcYkKWt83xwZTxKb/j5
nB/JgMDGrER+oglm4lmbxGWu7b30+0JObf4sRITQdWkMSkvTk78G6iV+9v+LSsBre+iuNyNt1NrP
zh0nKccGrcdHoRU9aii/qK7RThGyDTWr9Uz+S17QBbLKGaYN6SHrdGXsrAw4QpBgN6CkXVd+RVmc
ITpCllwG91QJDcvixBDdN8TpamJH4ZvR/v68Ti2uUwMIGBkfejGFLbdR24W7Q0nTn2iOI0QKu0PQ
5IYBwsrm20O43WtrEoKks5QSLOX66BkH8kMJQ9eCSjigzKgqaAQ4N6zuhMZhWG5PENOOo130Qi55
SY+UZEMbtcQPfpD0tYUpnULaZbtEMHNVud0Vy/7TakNyjJwROmscXQdYUj7B0mqpkFTQDlRtUFU9
Is/PTmrsaOT1O0/Gigt9LIqQWE+FF5WS0+856izBJW6Vfek0DS4tTPuYDTON7lQwVtKn12OWTYIB
ZjkpAItyK5a1H55uig+smqKm6sxy6x5XxqMEUEgTTP+Br4XlzB2m5XDXwg64ticKdCbFKobslsQj
F4Gl8Aw6+dU32w6ZN0jO/aYCz+E8z32T0oFYniVUyQg6CjDN0LrhF0hKIaPLlxWdvIYqmcWmPhQC
ttLkYGTrBz/5dIhDgkHcuihLAI3ft6zF5ZVOl+7xUaobZ7sIISt8B2oXpYmMpdOPLIT1eYJPOoIZ
bqCd4PJHfWJnS7+Y3pz4j9/eRGpFuEDMkPZWybMHUkztlCJVtH9ioleB0XmQOfZgTY0UXWN/MEhB
pywkIgaeteoxU16bMEQz2+GTcVTs2UdOGDW/r2xiFBE8UAZbamuxPNwSB4gMJdy5zgSiLId15Xmj
ziD7MBHzukKxRl4Bcp1iTf9PRYcRR6A3eEB37ts8D8zJ9pDCOc+neSBXAsT+g9+2+2y9EcDRPCsP
MPO16MndtUc9dkFU9zPH3tVxPBQk9MBLR+5Y65wb5oOsDQHAiZvT0X4FnK/VM9hpz6mZIKgmBQ74
BXPUboiMyV63INELkLZg8c4lmBosKo5i/u2JeLMYp1zwp887G+qTMbwSnrYi/FRil2FaHGGhl8gc
Z36/p7avnzYBvxbdWvR4aaAnajYHwbA2bzRWiKOUhiibamXakz+7Uc2fooJdTaw9y8iKbLO/8xSr
lNUUSoRTORz3xjxtyWJN7u6h6oyjuZLkRmPVS6w960uU1u5yub7eV8XcfcVOQ+LWnL/EUZDcveMh
6iEnj39va7OWBQunQ6u4Hh7taNxwoQijtwMbcrSIi92aI/fLucNf7envENtFZlgisah/SaL5jf0A
vhERJnV40BPAvw5nRQULAv9YoW1/XTwUMiFJzAq6scOLiw4ugkAIvISCi2Nh13FSufjHQfY48kpH
+95Sm7pvje259czmETrEcN5D4jMIG88CJDaVOry01XyNXa15+cPMZ5uDQGKUWjpoEJpdNVi8BXXf
6qEI7d1437KiQ/WDZxGKIVdgyNoVaeQmnzOdJBLF15F79cWI2poaedd3jzCQarmyqzs5wO7IbOYy
2Q3Nz7HO8tm2wPc2Y4z/dLl0TLAr/N6jIfGLfISaeqRMb14P43Z+/W7HhdFE8jHUiUvijf5hUuWq
trQpeJLTp2/DR65BEYR1CfccgRTTECiHTb8MXDirs/344G08npOtPywLXgrqLUP8Ldd9AFxjHIrj
Ih1W+xzHsoqEh8zy3dCyE3MJflT0T+wg7K/Y941dLB2MjF/qnro5hcItXlubsYFT8Sz+djsvk2W9
Kaj3LX/cv60ihYpiGTz4xsp2dkXTfUx1MPesB19GVvz6pJIVKpiN8Kq8GI2ylYGQxkK58sW2mv95
JVM7ENpJdI4B6daW+LDpdI4WUOs+QEWsgT4BsvD3XrGqv+nI9sFTwhJhjFsLTqItQq01ZeV1jwDZ
Vg860ojfVNO8MYvU5P5e9O5dM5TZlkujDq5gx3POyd/F2tXlY/7wIYlhRs+WzUCqF/jKR60zz/B0
k3foqjSvQ0BYfP4e0KdY2dlk75X4o01QyFGkbQcfYDAAyjJnsifQc8YyDEkEdHB3TIrdyI/fYgea
RlZSlRBxEbxe2JY+5mHSAVsi5zeHWVvQWTHFkKYGmpItuzTdh4o96afZFFH8s7jzIkL0aKOVTkgg
94Tlx/6oZVqdHPtZkt766ILp40OYY/AqUdWWFS1LVA/FFunB5cfDp86Du/8b/O4SR4eAfuKggf4O
XPeD6a/nssKoGImZrtuwjFdZUxmm/0saqdyiW600VvFrmgfx2XrqxnrhCPGtk007EVVHEsfQu2RP
/gaC/CjUh/DRtf365VllOdJpXr42t1+sdJBHzU1PXOeDFIjWw1xJ8M+h1Gg+LyGJKX8rdOhT3Ont
qcjW/cwJ0G60W7LVKXJt8YkFNVE0UlMEcZyAWVKsSAYzRcTqgH7x7HiVlHY2BVqlBm2cuIqyfjkj
lpxGe0RHeDfdEMChKqLtLw2GbDy+dpcOJywUkvJNS5g6TygACS17tZ7GfqZg9E4E07msxv5nnEd8
u7Qd8NeHJ2j18tVpRwZ1anL3wAm/GeTe88y1efZqhJPMa57F60kj3N3WKpy031Re/hApBUfafh0K
XiO6mBzujXuQS9OOmGYOMjj6gAbQ6JRrs4kylk3sB54SlqdGSCXHf38ls8kPHrVqHcKEw5Bo0zyl
gQanvMNcjP3DiKHqVNFGPSzzlqCUkCRjQt7ajJqDcLkV0o/3W1BTnWxtKhU23Gi23Yf+L3Uw5HLT
jCAgdLtUziijB1iir7YuI/1MqNzINL6IHMFe0uiSRc5HCJvANwidU+piX1X04DUc1J1zVp0++VTw
ggK8S6yjkwukI+HD1yg2GMbNBkeHG+BfEds/Gz86rCWYIEWPvUT9DdKYFhHXC0hV3VfLxdX+iGIw
5mcde/XH5XIXJ+4kax3DOnWtSTChD6HqeqPS6zElrl8GroHOa3dFXST5XVlXgYjEAv+TbmBfslkN
5XgHUwH6X8AKE0FJGz2Rxt+PUeqaHIbx9qdhKca0m0l97oqu5aTZ/UGUfU5n2jhVAuxD2ZpTDhRn
xSLqnKWGS7/ny2Sb1135QNw+f9Pl3YoVw/35GGvGjVw45elTtVu503F/A8swI/cokDA+no7Ynpae
OVb26kbpYLOvdXkoe0LDwwcUYqlvGI30qff4yCkduGtn36w5dOI/bTKbaJFgqDrEJq7Vjw7RmqcK
nkd+aTckXcxY/Gt7SxjETsMjUWoLcQgc2RKeP0QYlUkpDyx5T1zm26gpAxJkmVcqTptMr+H4zxif
V8BgPlAJImoKxkRRH4m8ddBGmerH//SMj+h2yrpZwrK9jAZogpqi7OdTf+vnjtfafpW3FLaewzLv
GnSS7uu+BaiymPbOu86qZCGGg79YnJSeZc0dpedabGgdXJrWIFb85XN71BCqvyc5yAJuO8OL13YN
iZQoi1xFblFUhzN0nywKvbHcLL4uluXjgLl/gmTVfOeLCE5uuUcz5of3UUMZNOEqn8TXCa0n61fQ
wz20mHQIegYE29TpHQW3FCkg+IW68upzpS2Kp7Z4+DyL6HKaWMugM2DcPTxQKaLHOWc4Zl0D7ruc
ExOhNC9obyI5hR74+U3PR86QhYZmClBtnkWYFEjd3oJJjTAf25/WTKxNn6KJK+fq5OuwoJri3yUn
TLr7OmEMR32miuwRnm121Q4cWwD4BbW1i8/ZOrKyp8GUkHimm1MNAauXSlNAeb0qxqcFTl3B76l7
G9Cnmhx6E02sR024rxHB8XzsWcdMDsnuvo4NzdlN31kXuyX1AAV5G5HTCYlD/l3OtqtBeAvv6jxd
zmOgjbyM2IG+gZG9n5BJIQ2r+yCHK6EfwZVy7Oufsb30usdnU30U/EyPZn/ik673UBMvcf/w2ZA4
yYCQjW062sF9PmNTu2vU2qVX7BBbDBi3LbFdt/7uIarqF/f5zFoblYGy7pNzHaWXAcDxsPgDNrKI
21AUGzHXIVXIVUHBuBk9VeG+4bQvIlzqSttgGllLVpnM9130qx/A3t3iCIRnu5pY7N2f6CWUtAVR
xFYxdz54/HkMKYt7qEbzCyQAPH2i3R4HKwPVDMMI0HdEaukswV+XULBl+K2dF3Cn0IzIhc0sS7Y8
CfO9l5+UZSQXCjGs2BlZ89q8qiZT+GdohpbCk4oKepaa2qif3whTDRhmgNvzfG+VsojzWe5zgaNt
HCepPPOWM2CELPhMAitDBpv/mfWDlY7023fCw7B4og7pxpSJmXQY7tFVXkiktzlgfdZGjjC8n3kM
1QQ76ROg+7ZIeHyE21/557PprHf+VqJy/bPROmeION/zQF3FGsDQc5wtlWSWqOsFW10K1YPMyDDB
wZZXxbJJe+j5FjZAygknq5pGpWQCfDruIIk/TA+KTYX8Ru/Aa4L/exgQUSrocWaa5NRMjG1w/Qw5
q+wEZjh8zv21QFmZ/SUO2PtcfU69+qPW6pStJJWHOJoQs65TQ2BdCfUdrg73tlk/Qmaqxlo/Zfze
DTBvDn1UKJZwvyuE5oBhDj5uCziB8mdywUxL1NyphGe+w8aNSJEI301Z7fR4eqBbJUVhDE31lCVh
q9iy2phtuPoQw1wK6/dDL7AjyfRjNcCxGGGJXULTtTzjE4ZMkiKX+2t8Wg700tdUtf/VWEgQZsa/
njRMaCKXEeIDer+05jLr9gtvKWk8oNrXuwB0FUf8KKBfD4NPhUOy9DU9BcsV8Ajg5Ri78WYQJ+yi
2a+SIRd9L9QA9urOnammFKpAEqgGOu03NLdayrgNJWK5c4fd+8/WUKA+ZE6BCQxrwBvDoGspzRFz
br1oEgh4rbc83SLQdET+6uT+LnSKYa+C5FbClluBKCNd+IvQOi8XydnWotSleEJsuGOlkCaYrdGU
Fjh+U9dgX9wPq5zOCNZsi0/mINbUzgK9k8X0jfEArEcE+3+KR071dhKMs0Zpsa5SpZnej6YBZkMR
oj32wlxfYzhFwA/59SY/8loHZWr9qy8vk2WK/Lk+zF7mNv8s9w74J/gseo0PQi8+ufa/Padp9Fxs
35TRSnSmPvOva9USgavfOqXGE4hTaWVXeEMhn47sp/SA8IuOdeEqkVYw6LE4DLAHGVCyvLj71RXI
EN/GuoD4C/2HizeHvQZaAiStbXhRjXIUUmQ3Xv+H4Ma7Y9Ze6I9qhLQrsH9KslLgXXS8Br3/EURb
qi1holFjSn+ORWS4IGgHVhHOzBIhrg7RKDeoFotAJtOmUhn44ih3fty2O7abTKO8S5xTrv12O4iZ
LmS4KsPDq2gJjqapLnbcINMoQwQO9XhiHqp59abZMdhONWEMQ7Zg5rS1AKPRAnY1QXWrgQxjhDIH
On2BUwDcZQ6WEbT94k5Tvo6hWvwRLAf8o6Mn0QRIvxbJmDL/9R4tXXcrSzqVlA0E7FFLp091fiTX
gXxLDGK9A0MEIUatC+ygdAK8Rist3Hbh2m39RzK54b1aVvZK8dl7PdrliRHyz024dnQY2Gy4yVm/
pWd8GX93dmzVMphI2C9lKaz4bh0C8kTpZgZUbwTYQWKTidF0NYDlDhd7I6bae4uvcl9yJN0WnnGF
kC+Dzloj6bm0R862kfn0WGxxJbYl264YF0wxSU4jTH6GnmmKqfhL2m2axUw8AcPq/xl6rPhjd8YG
RwA+oo5r5jK6rTF3vxyD6nhnJure8cENUF9bSNRGpVhlHer96eiQvBGi4Xzipabw06IT4HNYG1NI
JVyp9nk2zctwOfLGFSGuYkm6iMUzlRpvc26CcxPOXHiTCvn1OKk2yM4AL2mmkvoib8dxfTyosFr8
fDJwD3JRq+RdLmOddA5H2AaQhK9BSAraKkMybyvAfv+KK7x59FImcBhZXbKWx/K1cauNTQlZiqc4
3LlgCLFEMNdLoGIsPUYg32z1/TmWfU5VMYhyPSahBHi64vGJEaAhIlHFjhQ/WqAuGh5O6M7p23Ar
ZP49l571S1JykpTq8yczsCS7aDl1fOlGlfYG1eVVlFnDmeRp7x18Naztudao46BuDqxGRYjAO3wN
hT3IOAFN/x3FKJYKmjMZ+a5IZqp6T+bGMnxHs6tewuSoRG09SxdNhOKQgaZUNk3NoHxsUEbeRzno
9rY+iXpFJ23OYQjYQ7RB5UjdHXe76Bsv5Wp8PckvzFe8w1QCLuZoDRuYS14pIKSKfx1H8DSmzSt6
O2abcwJI844Ep0t+z/SXl7LM+V1s+LXJYEHfrYe9nuSt3PnXmJPszzVpZCcDLpbxoJ78op7aRR2t
kcrvYaARJVqSCIqMFZtrYapR52mkF6kV/WK+qBg1hhGsBfUS4O/H0X4ruqUwecF29guPzvyLAtSQ
7gXmUhPz6kWTkelOD9t7lw8iTH5SxbxaY/sFzl+9Hdft2mBNVTBeH1sasYNCNIph9CbmNJRqy8xr
+Bcqm8FEgfp8xjoyYjUKUIr8WQW/IcyNBAMmw+nWpBU7FmkefWOh2Pj9xAS5p7/5cxq+OI29mirW
AnY8XBOw9YskLfQK/ld7fUTyjd3Y4im9/+jhxCvZJfqms+KWyX7aKJSrEw4BGOcMSt5w8quH/Rpn
/frHcjb6wPERMSp4HKa93+sU/+ss7dfaYy5m2uSUGCvPn/z9UOuAN8oml5kyuGUPQlM+znAWQNuO
p6qEx649u3r32uqdG1R7h3EJbT9gXQhG18g4YXPbv1NrW0Crqr2HVZPVu1yNIkS8f+eRfJtcFZUw
QLYhDUoWgVY1GWIJpwpY9sO53SVQ2CnDDhkBAY6bvACdAVs61Dciv2AxjtPnGFQQOMkyjX3vtTqH
bxVW1vWTQj0IaaUarMDsWAnb6Cy51LsNLlFwMWx69x6EKF/iy3ACQbd+CqjVXFh/WODVwScgTzJT
RmRd+UAm+9r8DEh1Bz2MgxBeUE0ztaxwUm7WgmyDVTTxpGVzt0spIX96GtNYI8tgJcechBrYh0hN
aPsx+m/lI8/H1DY9vR2uStwFHTw/msdNHHjjXhYZyQn+c57E2b8uGS+cd9aVFKroyGBKNRrxeg2V
hJvJ3zaHnk5UFfY/Q8zbm4ZGnP1wcSomHcswepevbiPxSAzfpKvF5Krmz7q1Kn3VupRGN5ifuWRq
TYFaBYPaE4LDgyNpsPyzR+zWFkNUtcg2Ad8sIB1VRVZ/uyTc00RU8F1xrO9NQfRa9bBxSeWqan43
/UHAMyKwV2DFtohufj2wGgwvsVWfCn0/7IuiDyc58fgyker3YAB/snZQm0u2ru0lHWfJh5iKgDhw
NcquH7wERjKnvqP39IEm8mtfkmiH4se1vM1PeyEsFWT5zhO2xrhglzcWbJYx0yK3yb3aUBUjGfKD
8I0qQRh6sVVUuHpQ/+6KWrRiKJzSHxjGImpV9VY6/7M1QWjT01lZ61xHAbZDNJbWjO6CvartM2gm
HKoFHuW66jmSw95EUxaXAnK/6BuA9vbqW8TJpnDhr3ymhVDU4DKGtRDgGz0TWI6XbHWybPm2nt7E
AFkA6+h+g2GK0mDC99fcCPjAFHCytbbsPEH63/JK1N9yCaC30cAMsMzl4Bx6xlWKQJmYenDvF287
0wbWyCNQXVs6qCIxqx+FStXZ45vYBkJRF1PRXjd1FciYGZ2jaDbNLHdlZZGPirdHbobEesKNOUbu
ZwVyv8PIfwqYdCUa+jsWcQvCjs4JMYVjiW/AJw9Qpq+MUQtIMD25Fvp1CEuW9FX/JB6GcTWN9Wrw
MO3Hgzume9C3ib3SQWnLT9oEUZ5nk5jQib4bbtAu3159GLOgpgg0GsAOK/jUM2XUNz7iEyxfa8x8
20K9RMDC4fnYiNsJfSelXmSuXvQ2qcL+vMDXQtIvUrulW5GkkF6wd6EY8UMI9csiMnLDMKR1WeeH
FJuiXw1M2xLk3/nj2FNphKNgjjZ5mvD2XVqijpmWPbbkBcLUDDRqHioF8cXQzMO7xwZJw1q7Iomc
JtjAglh16Sxw1nKTtDKMnfxbvNvCIjqHvhOujgxvHEzHcbbT7/dt2Zhq9YXwtpIp0fiTxanS4h8N
YxSOMSd25nnnpzLDJ57CP1DhFXVFQ4ArfqC/q08zXZNeSBZqPIOlHrbUTyAghqeIe07M/eKa4DLy
lVy13bGgJKZPayTWqxKQT0+2QCF2mxp80WkTDP/d6NgMEH+IcCuldKtqvZvW1ANS3m0l21xeZM/z
mOgTrRGkU9btXKRZBqtBceA5jAIVWQUGOhgyQ2pINQ6FZvMJ3z5BAjd0leRu7ufn2KYU/1JFyPSB
L2nbkBpKmDavgVhhZZfvjFsO+EsHS2A2hVByRPQ6ovQi9ka6HphQYO2tQ4/pcwCzhNydoV0/CAl/
7baMWR66uhH5PykYzjLKXBzbaOWtQ63XSpolEwgpf+P5UuXJFFlYEBA6NkJYnTBYbP/4mpOXYzGc
56dmpmoEOLkbBUtBoNpOYs2EDcMAzmApp8ma5zDB0OXXjQiGL1W2Af0FLE+WR5rzQUV7Cv0WuPLZ
WTil9FqbHwfolKtjSLxGWzoSeX0mku3R9blmlFXd6Lec46YPwbvKzECSpn1hzgM5Qn+V1F9cohl/
D33cz0B3v9TfbOCbEuVbUaZnHbuFm89JWRLhilrHFCRkZMAsREPP7ThvOnCgsleGpTwowXFoQF+p
RkqlqmeXCk1W2WiwIarVRKvloRRTyR1Q8FDff3M4j+NxG/EkzIX+FYuYjNnwZtyOw69HY8Mdeheu
0VLVZyGvGhYERLkvi8Ow3rD/IMBsyYH7BQbbMo/3jxp026aXtmU2yvsxanc1sFLdh48RUWhwXsFz
4fBSXQ3S9cxJbEarpUV0AZrIg8bcc/3opOiBdlFT3hEivK1I7NgQLeelOf0CcX5kEo/o8Bym+Qhi
JsNAhcbKo4T631XmKucM4viogesb0IKoda/ATHBNUcY5tZkC5JA8sSk89Mtts+2Le9OEUeF6guqz
XizgyUP9czUO8ff7gXieZaaBR6XyVIgQucy6DMqlHhQ+quYCuohUqeHrwBa/o5duF/a5Dg1nxtb6
+TTAPY+jZJLMVdnJJoy76HENuH+PrC8GgSVt8uBJKZdnvcle6KuIsP9g6sgKmeFIbSD9YSaCuUeu
f4t0yoxGyV/HmelUhyn3S4Sz77AmfYQsoYhnLSpZdA6aG1z5Vp1Z71CimJvbvaXtKu6BHrCm1QOC
yjYQxlMUqwwERTMOnBCIMXDKzKcdXcS642T5QuVMeovBGpdIuUbpenSQLf0soolJDpVTx6oELHiW
R2HzVPR94FyHoJd9MNKIC4XYh4XTtDpRYu4MM+racvBZmfAM2dviy7F24WlVL2CFitSQDAp5mMH0
oqPXvYTx80Tp0hz40cY9GHTxhFqLpERAi7hL3rQpnXy+rUPcLGrrCmJS87xoOO1ptVBGgYwW/f4n
5/J9zXAuEexl+aFu+xbyJKQ4CLgdZgIkFhOvsAX1ojRAONSqcALGc3yjN3XNWedo1EtbdUD1Qw2E
vPMLgvGPaTvQOENKJeVYpUbU/lEE0YqVv120gJNI3rndJWNEuInhYQzW7WVeB3GyQDPLYyCEx4wo
SrLG0USzSNd0A7dlSM7zQyOTpcx8Ib3+tiSyxNntXc9Si3H/WFI9DDmsZpV5RsTsfGtAGKqangpT
N1hQxTAR17eaX6sAKMvEUGzbMwiN+gcDB2e23XSsTfo2hExUjI8stdChuK92rBxXKM8/cJRkUDqs
Q8vddWP5g4MKsK2yu0C3gnlXCVCLjP8tNzx5+1QXqEa02K7gq3K49asqLNhUzYImdMvlGfMhN/Jh
txJRIE33qWzHKeU/glS9DgJD+gglisaqlIMLcN4G6OtZ/vzeXQNiHVFWS1lJ9FmwvEeYTexliQyr
YvH4X63sSjG57WHmcNRnsPMx5U2r4ZRK/WAuvC+GemwqcqknWTKLF8mgjG2uvZF57wE8FxZ2MjsY
j16LVK+eeD/y4oZZaJW8tIvghU2GmbEDESJ7rRSgJnOrQ1EQDj8h3w+pK9Z293RrFCitVgCgfFry
y916QSlNDlmxPzmTFZ9DhVmWzhuRxansJfBEIpdHxw8b73mLpLFOYYIQB7aLcrO3hAdUZCAcxJvr
TdfZzClV4s17+6CQZse6rdnl6mnbDAY/d6zjv8cpGQcf313GcMrESOPboKLiSwU/2cUxUx+y+kcj
5rO/REjJFfwNqkr7jdYKddiG7de4T2yiP+PwRHDc1UDsaq36LqbG9F3gFBT91kEaDbURzgMpxgFL
l2+jsTIxeKKM8Ah6zxJ8EvzVKQLvOA/fkmKti9UQClzMw01a1TtTULqWceP0MmIn2I/bcbDy+hoQ
1/54ctfG434+7dtDKfl6o3ni/nyQA7E9fB6uXa9NwVOdudJFWRqZiMfqzzhMIKkQy9kcblkCGLlm
iBbH9tsAMxJrZTxCIfD8//k3PnEkwiPVBbZpKdDMz+6zcreo3yzPF1ONkkDPv4r3UkFecDwj47VN
QA82GSWw9d7pE3lyIrdSGfAqWMnJ7qm6n4gxbg7TKgZiRCgRtafNEAwRJ0wHtOXgHyv6YLIWGF6g
tnkHsVrJibokSm0VmsZAIINCOenstlcU8tHXJtxex4QUY7xME1/74ED4jID20KsS4246mE41IN5p
v0tfqaMPORFhO9OtaJsnyfarP3GUtm9JS/ReJQ2CH7na7iRpYaj+LblC7zGoCvYpPkfoShEIE70T
K6ecpP3E/7aIq5pAzcsSMXR4vCcjpJ7qzW+XcBEhU7ciZxRjSD9XMmOIvokZ9xYv68yCUi9TWv8h
b2UI77/dkG4H+DSqNt+thm64kpna1KBpUetFlhA+6aWx4cqgJvZ/gAbXBn1lAYPhXdy6VieQKNkt
qNt6MbST+VyqwaLubH3fDluEN0mQxcipA5Zpanr8DCx7bHKlo9gFXuc3eNq5KUnUpmTL87co5GOP
8wakZrWo24QtMRt8/Ymjd/ztR/u39+qBJRRTAH/FkWzSMTyBRGLBK0o7gGmogXtjT4Hz3zuPSN6x
y42JuaWXHWEc/3F+KE8NKGdES67v1MO3c90P2pufNZ+jhJ5BeCzEH6589+RTzzl1UUojn+tchjTM
xxlcNQnhyYUZma2hB8ZgPFLEdeSkn+B4ixXX9QoHn7Bh6ubuMKRRrIlhm+vx6byU85IMLzThVLjE
dLo538HMyyN0RjoxBms3oAkPqVrIePmAiYbfM3KyYCHz0I1Wqm78qq1G6TKTUF+KF8MAglyCbCvw
mV06Uc23mYklHebea5xaF6vLgsfH2T3hRtCtVQivczL2aX8VAIHvfqdsTb5w6BKTz0AZc7sjD7gy
8/TP64vNrNNlMWNsjX3CPZO3DQJVzQvIsBSuy1XO2F+nV2T+R207VGcWWBB3WorOAY3rFNDl1D99
URMslPbS/A0mmdHkZ4GPIxbHWZ9SodzlgyRnJXnG06ii6HaXUPt/AblUAFnVp+QSEl2qZBWxp6u/
bqVEkPl0brTnUVzDzVfH5S6UsrIGvhlX/kYocibKC14je9IPgmR4mqfQGM2Qxvs1CMmSb73kaQ0p
eCq+52E1zWo/efCeIDBp2BZ5xCH6keq9xIHZ04l4rl+4zcg8ddp33cGo3MNg/f61iVnVhCl6OuYV
S/t+291dJFSpb5vMYpZK2bCoGq+14vzoLtbN+4mfP9oY8wM+tvaEF34n6OE90zkWzzpqPF4JYJwc
u2XIu0gUTdIsVMV8RTXBZ0t49/FrghYKZ7lv/sbdgABDFlkzLbAJPheCMbwooQARao3NSfnkL1Cb
atliGjjV7Ix6zlKZbkHffCyfzc+SedXarfIzfQZyv9wfXNb8W16icXEx1LvcYqblj87nv7euhNgT
svZ9mzDRo3jGGfwSv5P8LFSPHGl4H991B0FbfN1loWE8hW/CVff4l1XWa2eQdvHD/2C14Ect/s0a
6mO+P4kNs9w8cZcUJGF3xPsz7XUvPCaKZqF0StXUrEMLxPLV+f8NWs0rT8VPtHRbxMsqsGBQ1tqt
hN1DG7/0DXJh64CwHzwxdhTTuf5ieD2+LhjvuMRNQHpzHN7TI/MtIwlsU3xGWmLZGpOUjB0xfRQR
pRsconRSICqGaEUKkcDiX/+AaOFOnlqIywLfC/qHiSsUDwHytozVbzvFbkeGXNdMrJogvsS41M27
7pu5hly1azY6PRHscdJN7Ea3lDFT9STH7swjee+lGTxiXIlppIYsy68fDhkmhwGTn/52a970o+w7
HkhM2ZyxjzCJCCaSo2kL4vBztZYNyHnVjGbEHgVtruVYIIKElhVhGNkUWyiY3MDO1bKk0Zkd/gnS
w/m0xND4TtlQb+MfoWHgZJk7e6hwRgsXB21+RxJjXMeNxHo31x2zIOruD7zzLMX5IvvKGPI+FSOW
Y8tI/hHRnwAkM7mln4/Hf6bu1QozXwKQ8QOUPVcmk2aq1Zyl16qfQ5Uo22yzOcCWJn9ZyBt9i/+r
DZjInFKuh3R80ndb4WYhce+YezYvV4l4RVZkgUJjpuDJsYs3dOGbItyvnYJBDNNpSUo/bCFsiijf
+0bS+OMlQVVl89+7s2ZAI4epQf+e319bbe/s1m1PtqyTsAbOHSyqt1TMEc4tzPAywu6xL4LiQo1J
imZKRe1TVnlIzuaYoFeZMVGGX+Ot3u4Vv8r5Ju6ds/TWFu3gxJGXiydMi3dFCoFZ863DSOpKjFXr
N1Wryl0Jc8fVykC8i6AclWxoEu5N1jEQY+eXmJZL+7V3dKmPXf1JnMHZcMtxX76Fis5oVu4Hp9v9
jpn6n9kZvBTosQVFMeFDsOXLcIyGJh9K95c3ZnTJO8tW+ST+SaCgJtRJPN22bvvueE35l1q8KHWv
kl/oTaTuwnwgnxKJ4fAaarrKzroUIv27665VAWgKHC5r+t7hW2IieOzilUVT0cXmfo3P5U8lgomg
xkcXAuaLwc7FIqMElVZuzqmRw+DpEaYm9UhoHO3o47JlAqgPWzER1dwYXx2TJvvzbaI7qvTLm8U3
kLO2YIq1mmjoIYzTZZenFrRC+kHameokBo/GMscSQ1c+0Gc1F+i1fRG626pEIVUtMiGgjRX/YoJV
fI1ab5y7v+bIgytpLcrExNHAlv8XY/nNZji5omIYM2ZGs9aG7OPxNczQf/m5KOQnasSxb0bq3t9g
4sq9pV4askzRn0pk3n0TsbW6xU63PDlC/gjKwbw+lzSq5Ek00yN3k30c3O1/T1ZJNSEwvnakqkci
M0F+6i7MvG5VUzIDWHGMajmV4YE/kGSBgUZuFXwZOrUm6vw+lYr48vsjC9yqPzlBsLyzCWh6Mwyd
W4us25p1DxyZqVJrJ6TNpkhkxC+Qi9tS9Eg9/T5c8vbmBpUfvyd3aLFeV5AFrIoKpQwKb4AjarlK
zc0OkFM8S5VVfs+ajHp00xQ1BEpW+O0FyWYOa1AtknIMaADCg9yN00rBb4lGXw9BHkz4xdK34GDo
hnZ+xMqWzXgpoufQmVKewDzVqNcd3s+PcuO0lL65yRfwPjI9+BBQ5sG3rR7m3sYB/QTM8WmAZaIg
ZvjAvKVxfZT0tWSqlSCWCb45T/XpFS3zbQ9ZAj/PYCBAOkqiDi/EA/IgkJz1xzsRUtu1DvIMab8W
Ix+zlftSFdV5Z4gwgP41K0GZAgT9LPaQF4fdNkItAXuKftOgZBxVK6ZrnJpNefn8Pz8Inw4/clBJ
/xQ7PzotISdangKFMnVZ66O/nMnZrsL9cOZYmvSDGDtNhaVePa/gAeQGOhMTK9sGW24yxI4zg+qm
aVOG/se7b7cGq/EpFrBBHSnylAVjVSUH6RIVpyJWnm2c8yKxHkblBfUaB+N+JCfIHUAC9CYcZ17u
kfWgpxGeMtBDT9lgnpugeYL2/NnkJ/YaC6UKUEQhRGIt+0jkBItMXas8A8DXxs1lGdzkBkK/+ZJs
YgRN49Zm7wEMXyEBemoebFz+dBzibHW9U1q7CiyjZM19mWw0+BGBkY1heeXQ+PKarnQmksYFb0Xm
VRqgyle8UohaP0QHV5fIOLQ77X+pQOAD2uDllfaAJe2VhyY/zOevGuDg1cYYd+bYpDpAamQbob/V
iHNe2qGkfGUVaczUsba/h6Pf9SSxo7jDe0/9wKgpRZ+k2saiiX2WrJOTQOHqqd77nFO5dxO6pSEb
jE1p5FI2ZtB4MCP8gETDuElBvLA/EYFhDJBbHkhnHDQa55vHr4+9qqOcK7AeUXK5ZpiBDOka6Vfz
qWYuDltaJzl43j4RsqU7wtWXelvAEdqZGtgFRSLegeSXUTp/dBX2y7todEaWAidQ6cqSVPDXWVQ8
2D0V8s5rybgXQKngum9DGSEzInw/xqc9IgeDbQakNGEA9sI2aCAzhOoo/8qqMolafaqpklOtD/f1
zsTg5tC8bQDdsIi7mqHjcPoE8rv/NsL1Cf1QpTo0lEyv67oG/h/Obq5Ox+5JT8BM50XN3ZwpdkIN
GX57JvqVMw0uN3jiqVV8QDJWuxAHVJJeu+TUKasQrFchrkDJpRw/GS48zyVxb5da9sJfQzrARXrA
Aebr1+T048jvi23iNE0wKHOyuoPWuX+jDIK/AWNavR7sMowQRciciFnfath6gK3CPh0+8cZu5xCY
OE7al0jOYpCqYy6pJl/fBn0eMVFeNTrs6dfw37nSi1rabD9O00DKmjQNdd5B/J01VPug60dEHQ5s
85S1A9nf80JljyWKB0/BXBLz6cyY5MH+KOgt7WLasge9b2q/3usX6EztA+pRvgJBdU2S3jJ5FMdL
aZ5hpfPo4WwSRU2Q53vnKYaZ6PVyRkSAnqotjrU1+o5/RytOGNzTlVZqNV3VLyp1t1hXBU9U80Yb
/HPrzigvKTcH1NRvJX6kwZkoU/018yODYj1NerwfRa+aX7XvHM4KQfSXHZJEInqk8WdP/neDJQEc
Sy731edPmB9BjhZA/xz/eexCQ25aJdBsrc4uY/4sCvcbu/d7smshfzhq95NVTCiSG66dM9C0l0Dl
klYTGIzXFJQDlT2TVpuOPGMOykO7mCmaDeP9+rX8cvAf0TjdRvC6xd8vhwwkkY7eD0apOfjrLS7c
T5BWELoRpmWBeQoTrDkqhPp/EB4FjKja+WHiAi75+3lcSX7x7s56eO6fkqr1pw9SESTRfJk2jHpQ
3M0u/jJQlQOdmYkmlM1Dx6Kq3zz1McJKG+7InMgUYk4OwxNXfRntxPOiiEckpph0Sg3Z5cO97hTo
PH0YMKZVyiuBts3bn0dF9Hn8NzSn8spCSut0oVRA2iDJTQuKFlkdg4OsO+77DMVmnthEb63YLrym
LbDfD744jq9SOR94OEa7IDm+LKqgbIBH7/JgZttKi7yw6yaA5vdWv03fNWrdwruiuEk3KKKvMUxz
b20bmxN+6PUQup+UE1mJcj+Mlli+O3FOkHbnzgiyHgXavZPbmmcnYwMXneMD/4O2NfbiWfTLk9jk
iYGDpPOGu0fQj7kz9AJ0zSgBuZS3SCfehUVmYXUwY4e27LqDVX6oyqs8h/Pvk+40K/YWCkFKn+Rh
81FTrtlyjfYQk8ev91xD5+w3tTdfnb0y/N7YeZW0gfGN6RSlSWHuKi/WjZEas2wMXLkylAzebNjB
RoIJMlZqM89m9gHtdKoCNk8u1iGofrrFzXIi3YyII4Y6sC41fc1NlCjVUGGiJVIe1634Qwv+uBGi
KYvqtxS/W3agJrf9XPDQ2S2Sf1MI7glyYfvPcx4cdT2Tuc3zABKeHlxM57fjKQyydYXT29WhQNl0
r8LGI+feTUFQCplJi2sB4d2irSeb+TeqcV+0uivN+rS7Zl0vOmUoFse9bWOjXnNPD3Z+KyR2l69P
qQ0biKWG27jyYdhvomoQ8sQQtl2H+s3xqosW320ErrfWBzbgHraAvfefUsR4NlQXIf8RUsN8hjjI
KFg+q7IkJXyrm03q3e9tJhkunQzKCOGnlexfbxWyoRrLXE+jj25xNRnCHUK6ZPNpcBvJ8/H0IGmz
nk2QiWVL++VcfTXxhzthWfTY92YWoV7Jb8uNENJa8wAey+j08FwtHXPVigcppPrwad2vR1zN1XNU
Z3Mg7Mf/oiOKgjRcvSm9AZ7Kcnn9NorMkJIMrhrrhm85R4ttufFyqPRHap4sRHKfUO9cdOUResi3
MEt6Tcw06f5JOIJY9KYXuoW9oJnwY0zIaqusSZ7fh2Sm4iOg5WTNCy7GFt0Ha3UtjwAwufV+5FNk
WrgogoeH1LpshQBHl6zzOOBwZqCNtsAadPiaJ5CqETheip5g44n75qoGT+tPm/yYs34TUwx0hizx
9xjwi3zhqNIa/F643dd9GWNlwVlQxod6o9qM/Ilfkb9tE7x8jiyTWkUJ3Lowrd2V+IbCW2fytvFR
u5R/DkJPR5DZRhTE8BfSxADCfAMakT1RtH4RyCej/nUveGvo1GKnoh88Bhc03xFg3FsmsbjGdZPT
lRldCggBUbhAkQwbgGufJSj28/pSzl1a8xw2Tkp9qSoIHdaliAD5gYsbNdZD3PqJzC1/q0S6hqOs
Y+09jPAuYXdE3K7aS/4fjYuJaUVSkacpwRK30Z3HUee0eNqwF05oRCrYHsx9ValpsLQGHcGbR5b0
SpeNmVa6ENmuVSLqIESyk3ww+XY9kb4+wcaVVKilZKjkeN5YZVnKk+F6kObhRNRLtkWhP1l3JNPr
LQnrG+3F5w8QKYMO3jkqvy3A9VGfPX+iuUSQwDYVubRco+IuzH63rdhnxCzSboH5z5HieHPICxp0
qT/ousMbBu542lk8tA61YhEpzuu9D+XhJ51V9jPS+3GLVrrKBbzTvBEceQ9IrICeV3IkrOps765b
3Bw1F0jNBz4AqQUrneZrWwPK6YKkT82dcgDas9Qo0kfesy/2IjtnBe9o4R7gDprlZS/Mp7EgPAtt
gZ/zLh7qGCBT/1bjevbHols5Dwr40/z+i1YjAL1vNzcvhtBS9IvOwEGHQ/tEhx+WiTL8DxqVqNnV
JAexxE0ShWATRB2roZl3cJ3KcajmmEYem3xjzRKroIzQQAk2OykoEDT5X2iIKQO1WHyXSgfFucGu
REmjW/EIogDG9hQ4WAkYq37VYhRAdPTV37zqYjzE8vncQZhi2sDYrLUAk27x81hMkKdhIsrDC34M
N0wVAek8WWJNwHKLJxEo6kVYdhwNKn4XVBW+LfPcMd3xS1awWGSVydVOlMGO98N+MHexzbzZeSMP
U3GwwjlFIcf9Bb8870M6JtppUS8/YWoUNYbznGZ3g+idiw5tUtr4BI7W0BkAai8Z51kUc6KEIjwa
e8JDNXF0BxmWeDZuJUyM9c8OCw5aPGGnBSUhrCt0zp0vuAxNZWrG56xcowdwz1PQPwfnni748NaL
HmEKGAZ9bvG7lNQQ1bNIkBLgImwO+beslqV2urju+paq4DingiwRdUO+mZWOmVKa5Ldbw54jZhwd
4rb1jtApifz8rIvUO7h7jGUpQQ3p1K/Oadwh2NIxsgLbe4H3ar2xG7a6U7hBugLmoctHVaehyUfY
MVTYdomTb5UCLiuyDHRnjIgLrWBLZuGXwdrIJiOBGueFHoA7jhKKIsj5Er/rUEJ9FucpRbnknGko
O1HN3yvkR5Bg49x9uXsje5Yq52u3DApQWTgwhWAirrA7AiTIlgCxShpzMJZ8hVsEVPfm/8gsWNuF
PMVbkqOoMKFAlO8uHZXt9kycEospLyEk57FD+M21BRgLMqPK0RpDQZ7v6OCSvlp42qmuwBY4TOXx
VUE91PJo9RTQKMSWlI4JI0wnNhCChsPsewoED+V3HjoLdRPZltpS+g+6McrUSjXLf/qTzEF3FxQV
GIOmgV6VAipxsvA6W6Aq7ztZlmjg/5KubVEhKzs3fuN6QQgk8bTGimglG5u1+2jmWohDiLOFHF+J
prtbZI4OdEzAd71pLl8KTQ4uvb6WmB+B1c5tnjaiuWvYWgP16AHfe9DXBjqXVPjhhF8Sy2gxjMS6
jrKIOIOROfuomb493BAi3Pb0v4wbO/X/OaKaWpN8FVt8ZpXW+j4wRHK/b+nxSa/Sj1epzEC+ed8r
wy9GZEil6FlUrIGoJHHR6qzA08ryPFvTuaN5BKSiazfLr1/zO7yCaHi01KB5kg1qARgzpo9DBz1w
c0aCOPvn/0sEnrHPwR6ocRokNnZmaAjxvQf3lG3IbF3+/c52BWe56tR5/WOyg4vxf05MR0B4euiw
0zOlnaFSup+a2bNem7YvzA8131YkDB8RdxaCrhwlL10jf5v4DJBrc0Bk3C+Y0MXrpSKDrR5j/KOj
08qNA57H6+i91tSagnZWUb2UMP2GZ3maAVNi+SuYi0fE9vp6Hz1WjP13q2DOg+1N9tTEmAR9GF90
ABZZv2fdVAIQ+ebYobsKRXsqPgUVOeZphHLYOHekrkZdcfBCCrBQ/xRhuMrgsllmzgx51Pi5Pknr
iJwREIp5bLa93NALH+3MaHZRkbTGMd1fuIfEG3eRzycDoowBX8RxQwzf/7XSFGT+QehAvWqU1085
/AotGRRRPVFwtWHSGuZkfYG2N29NTOflfOjAb4mMJN4uyjogmEzzIKzNWWtRiab+vO2tWUcs3ha/
3UBiDBvZrj3Vn6yjVc8LlH5+dvUz0uqwrd3qwYbPXiAeNgJ2rMPvjLM2mEvCboAAlrfg3op52/RJ
hgtHHeWJxFJFOtFVtgSKyxn2y3bNa4UYxSnrPku3uYw8C1px+0PywkeLA7HT1e978vv+2DycSGuI
OUpiQHd+biq3J8rWP3dZ/tjXFFw9/Ef2nI+GrBEJosNtURXX63ZtMJLMnfUw5zFbh1Tc2SZLaZFK
VSUtNWMOtEc9Bluhc6SO5zON242hdjAnmUksg4mJ1w3GHaEZ6nr0Jd4HUUO/bGlQW0CgK6BjieFN
W618C++sI/MpSDS8LRxH+oxK9RCayV8hU7LbSG0pIhv2pPzTB5QemUL92p6QGnhkX8wqZDAFMwQ3
N086gXbS/oqSXBJLEI542n7EF0ilkpNgPUIGUiEXCkMNp+nR06QKVALmp9lDyWMRWpSXru/YuCDw
t0gu0PmrM+Vy7RGwkC1emiPG716H4egV0J3DSeOC/ucIeISItgQqMdXbe4/YZlhT49Xh1Y7q+j+3
A7+v/Cx4J4i/b0AuOsrjgyAAb/PD2ov/nT2DKhK1ibnzOUIDLtnEWDW/DT8gVogRrMwqtMmxKzgS
VY+nnuW0fjhr25/q+1gDRIh21Q4iCMmoVPiVbTy797P1fPq0nA2ssrzjkzLNSfvKJKQm9N3SjNxs
O3HbIFVZnKmybtuotL0UZaFWfXFno23QNHc3PUOSgd9tMO38TQbuThgKOjF5mVfblBiOy+HZ8Ix8
hTu5/b8xAv/X9Zkmv6KmfjgMe2SFSYeaj4ThzHjD4w6w6XhI91myydgfTYnXBIaXM59bt3NOZa+F
1VBV2HcWZjazQ8RGT9PhOziSCVPDVP8xCLsqp49CclG7Swjz6s7vBpY5Sv+O+CRgi1tQUzYHE1BT
ZR+33I/HaK69otN+8rxCycaNosIhPvAy09CA9zruzJbxpz7dxXdiSuD0jgZLqwzGumguItONrzHE
+vP7/EiOMPIZB+Qpmzq/1MqfQhVSnreminhEdBoqsssqGkeZ6fHyUOn+rdhsyoGqxNJ/XvXUgTwA
qkS31PboxNvMT+KmBPyQKBU0jpn4WYeDive9L5pQOow8jMj9UQzSWFR+QNOOSnjrkxbbOSn7xrPt
iN/9Bok0yqsNOSmCiqa+s9ypbM6BvFzeBUkF/FVnqBSH2OrLbe3Aa8t7Exq/CjQQu4QTz0FN+M+6
9aGojcRgHRiNfeQAMMVNxFJRUTXTo//F6ochF9BhkDtqxRqJhpV4e24bjzt1ygixe4r9gbMhUYN3
oFZ7hh1Ji05vdGvyDauI+12eXVcMliYjjNNT0A+qPX2057VHGJWAA5VhvOnPKhG2CzMNacGkkzDH
c47ibHT5IbeS3LqEi9UXNkPETTdyOeuDYHCFaHbxnYybQs1TEz1h0d7H6bN9OSlQE0V0EYHEIOk9
DQb6HH1h4TQuZnPd9DlgwMtsWAw6fd3FV8WT2KW6HWHP2/Wd014++pQcfEcybeiFr/oBGVe9o9db
P3WO+LfuinvSle4B1uRcREYYDMBVQv9+52ffWZuOMlRJ/y2CpxyMQNhcLLzlDDkROZPK2f8qwwBb
5LTCErtMezs7WVpMquc5sF8sImD9FHR5SJM8bnXCdmayZMhD9a9Au2GGeqcSldLsVf+1UiL38eXK
t1I5873eW9JsFUUvOSlgTck4ITfkhr+sNE/moBcSHmqRUgDo1hFL4OLnx2yvAjIE7qz8+TDXQ6SA
wPG5NXxat2frgyTgN4IVSwkdYk02Kue2+YFJAZsBRU2RiyKX5b9IXpfSpyffuEWmK4mqE1jUuykt
D+CwOYr/q6/eJp+6J6d0KzxXi0uq/n+q2JJTqjVZpumPrRlWWK48I6571kPqJAEac0rv8w0IVtWK
aKCdj9MHqPz+LZCHHn11ToS4yN11THCLs/LxN4Dy/KJsUUQMDcOBthBaQtLXuil0Y8Lscdh7zsg/
3+/dq2MjpXlfW0kSa6y0ipoVgv9WCBALBpq7kCNUA8KFuHPPEugEvr6PqnEF8Q+IEFXpjoKizeTV
tfy9NKiWjKESBEeJNdFh2M9eFKwXbY1p8elNH31AyY7XCODgQdJJkzs+80A9c2IFhQUCGoTpXUKe
bWuPtlg4YxHmDTrmCz419sGkugXTa4k6Rr2rryh02Z27yoYRuHeaQtbfyRKKnJk4o/0tMWQZMtUd
hv7OgmRadXqbKxlTPflU2t7P9N1ZB7hUoKJHJzMqmP4xq44eQN+Rz8QXBo+d9mIi1Yg3nAWtfUNj
avsqvylArS3YYk2d3PbZX85EwiOGYVogB4RiMDliENcCoV0dnkDQFhC2ODjnq8ioCWAuppFcQWFd
4SUhOFRmKvjDmsEcHXQCi7eQ/hygTnUw2Rmn4BANqsATkM27GHCzFcydiBNftkXr93Xl1M0KQxGB
pabJLgjHQWTEkF3idRh0FivpsMXFxkXskobaqb2Q2vt/abUdGbfiYl7FH71wsZ3EFYQS2kxJscwz
Yqg8W8SM/9GoPxz/1EjeTSdSCLY9WOZ7nrdP+qwHm9av8drjoWjChlk8urjMH89JgcE6uRyw5i/y
wgEbgtk15BJtbo59dNJkUc5mK2+IgPJuXXsjDv7xMQ8/KSHO+0WrDo1O7BbQVvTIvVS2iK0hGiQE
SguU/ykTSsytGOhbecGWif+fm/rIStiFyIm7y+E+8s5yZgqt3nrXAT9rZLIpcjp9biacmA+BOMxD
wgBVrfJgA3W3hX0CnMReSBM1N8EvKjKvDO5nokc4jz370Jz7bV8H1ZEdRKBL7JQSqODhI1g/zi1c
xPkh7nZgDoRESJjnrYwHtnaCKUPXbIRbctQGxeL7JzyUMxVchCWYxdEZyGp90Zt6YmXET1vYN2GJ
LNnWUWD2oRhJTRt8Zope0Y2G3K1icQoJ5w7fzr7D0XDcdBNZssgDE5dCJ2c8elMlQDybavN/DABO
85ImZwbLSuSdI03o8AIkwgJmK46wITQ80bTP2kyL+p7dGCRrO+MZuT8bzxTKh21dWem9Ukiz5Sx6
wTdJd6gGHU/ybZfUoFwBFLzj0Mpb9solfLylXbjUNjRJb1tOorjc+U0v+oPw7F2VPbTpv9Ny74y2
wY9clQH99Bn7+RLv2P2oDLvm80923YdNBGl3nphf/3u56fRFTAfj8bkXSMoTrLE1X8fU65Uw+e94
uf82RMGTVnDSbBAtlHWj+oiTfUOaQaTdjdEYtG+55u6/6RROskYeL39ZgpqoSmcCv2gan2FzAYWJ
WX9o8TjEU+myPUqAbiAoF7JVMsWEB1Kvw8hrjmWsEgnatiXWlXpoMs8NDbB7yP2fIWDeYT7Weq6f
+qSW9VS0tBsFpF445hSiRc2By4ETVNziEBKrH6a/++ZU5XhCWTag25NhLQEGAXc0xEx/yIcd8PTG
ioWmstWzBT5jG639PlN8k4k48UFK8Ubtw4QPjND4G2UcdH4ftO8gp7MK/+R0JHKXPLtB2Pnodovb
+N7dk9zWyzhUceegiJUI35BBIIvslpNGWbBHQeG81vt9653/OuFZxKhv2dcXkMVVsCCDmkMkijbq
RpCsBeXqIT7bGNTOCEfvJuS67R5HqUVBZS8VnEtt2IpBlbMpzx7SC60era9cCZgeEuDlOO7wL87M
5M5EncPwum8nFXIzTVcY8/kYYFB6lSQ2lMnHaBcTtMuUK/PU2Bd8r9hd2FigNrhruMBRGWc+CzgB
F8YGeX6npVFi8Edi+CeZDNTsEuYbKRNcW3neBK5ulysj/QsYDSn/W5mxk91NQrYAJMj14tHvm4zE
eEl1ckJBkOgvSTuud6+nj9hBdV0eiGKMBDkLcjuDeo0whznA3nIEoVgA00JtvERyW6JxuwqU02pZ
B6EBw4JYyTuKajiUsobZa96g1hcnCwQCJLZJz6xZtBivlQHW/822tpgqn7d7rIo9kpvOgLR23wmJ
0ahZIqhnuq0WoubxHoU2acQAyrgsmhicvIrlznNuq6LnlZbnRGmfhN8grMKRYxbCftDkHMzBiZid
ognGyEIAfo9B5y0EeBDgeNdDjw3kb26Tkm3IPMG3BWSwiz5Vf7UAjrLjJFKQy0j+uaGd4EOQf4cw
ErJQHDZ9TrDiVKMjujAnvjx9qyuvA8QChg3S+jyppM+6OLBApJ6V+/sfkTx3Ushqf/oBnOkpDB6F
dnl52O0oSpaYmSNr3FtdebVHuGxf/VuwmAyZXWLaKw3Qcj7Jq+KIxOlvVgw0DPVtIn25cFMPbRCI
nYV/EF8HlMwQQjXOP19rSTuPpA+wHTx4vWD5bL9vKbs4ZP8iqTA+PU2+QJ/zLrUemXmeDZ9PfNwA
YCVUlIyh1NxIkX8l5rfOLf9cbsEj13AaTtrIVy7z+WSJ/BSGmH8FtedJss9/L53/qIbf4EIkr3Ko
Edp0+6GALnwZrbW+2ijIp4FEWS958opMDYuhYtJuaavAV1Sflu1nuh/fvTUdyYrfHpwU++aHLIVk
o/HBwDYThtCqPJmSTYeS11aFh4fE+7OK6MhnwDOQZ1xiYEI5YxyAagtbJ7EnBnglfvql5qo7gcwU
FtsRAsvEWnfWM+MTAQsEctDDeMnmYA5TSolei/lqNp2scxY4z6ukN+GHC7C65JYZYVkY8JZ5u+xS
LWKqM5r1yYUNBWwKvVpKi2erC9y3meJPVsmtIwexPsE9eGTagSrdwpbYHoeZEEqT1RCT1qFIu/Tn
TDg+GxGKt+GS74rgVlmt7G6h0hQwtZWSzk43GaPYcImoniSj2YtC5vwpqp0Z90ocXXtmbulJ2utx
dTKf/d30NWTrbSG13swd2Cn9WqK6vwXSEfA33qYowcNJifQiLyID9VJJtW2Xmt0eWV23kWbX9Yfz
AHOYGX8wQAkXUuiSG0C+82o9hA0UJrQPhERE8kCoCTYl7jxUMmcydvhrld04ck5wShO84KJOgxk3
VX9V0ePwJHMJCOGNvZadaQlD/ZonQpMbwC5Hv//BD7yjWeqYmwdWeBNVrZUYnuwTb/LmunbsDBMH
qZJ/9XSEZCQ92DUauZPJv8W3V73NztdxSb04zphpMlIa+Oi/cYkANDU4smyW5nNzImC+nrLSdNBb
UEd25EdqF6hAFOwynzvhAt5tafFOxhM13agc3d+VaWeKWZsa9xNzRfnJWMq8wF9rVxNmPSlSvCiP
eiQKy5w9237M84v1+nSY8PDYFJTnrO+cCch5L8or7iC+6CAhrypfG650KqZr2D/1DCKBIR2C6CDy
GsPStiiw9l0/G6g6wHrT0HipiwM/KqiP6c6hTe772Q1UfDzMeyamjAei1WMOkxvXD8ynT29mMSMA
n+0Vrcggzjz836L27FO/VWnYihmF8vSl+6wYYYJI6qb+4woJrdWbqoV63JcBH3ZzlyUTvfumyhxe
Z5a/H1kwCHcjnxH3TdtkVBpPqJKzrQ77Sxl9dbEbKYz/e59BDO5DhmP4fh3T0pq2j7NLjoJv/A/j
K3r2rQu4Tesy+AIVmyFmOPTAzoNh6FccbaDBDZOTWGAPXU+QzuoL1hfLQZC4zCu/NVTyacPcZlXt
wqO1tcAYWbcSkC11mm6D/eXmYfSMbEkAunC4ttXkwi9LpIBHxrfLrutDOHOQuqot/LXmxSD97+7X
8pJe01m4nGMlSg43eO/lBgvk5jPhTGPivVf6Qv14soWEW9Y/s8rdhtMP64qrUi4YYSAqAFAmI+Ff
lgJm+AynqU5yqBquI7PwkqHA3DhHI/3RwWUCHFQup44BUWJNuotuEifvcMF+rSe5mk8JszoEGqfR
e0m9DDWJ0u+dGuxBY8Y7DmfRWDU51YPxEOX92WNvNmzICtBWaAqExw3Kx1/jd0mMALao1q8rJWCM
67mo/eaMXDLQtrENdZrBJZK5/3tyVgxx42Ut1WIJ01ddr7Hc3YGKEiS3vay7AEjuttBmd2Q5zOrA
PjvzkNeiY4a3HbgU1srbAmHYIE8n8W1bLRgSRIG2PiXrIuVcqrox4MkV8hzymdS9zcYnXcJeCKq1
4GRSWLgLL8bnyg0wbbuX/zQBVQOW4AV2FFTPLliGzgpOL8Z2cGhEhWxgWeAvuPb7VTk+MGLCqN3q
c5+BuLsu3KdrMhLo9gbYsOWLjC3k+764jKyvzvAFMYwaBrsVVGD0PP2ijaZa7ii9OYMyAb/4aM9n
56i40saXi9oUHWAIYZh11KcHjpgzkaIoufxIeKBQm8U7APfbTXEbY1yZhvHK6xaczmaheYW6Fojp
xaHMC5CSALclAUY09yAzTS5rr7FPgU4aS2HxUu8twkz0YGMbpaibkxLn68sOytoRw+hFgv831Dsm
TnezJm0MLMZ/KkvU2d3Jclf+fMrbuwh6KAZT0hc9/K+McK8ay/b8MNlfTdro9McMqpKA9eUcMfNJ
Uvrzvr6pXXqo5+A+qYzo2W8xnyvFbRNOHxQGgC5LpcFroEE8D8pX11zQKL4u2tgSZpAtCPKcjlhi
cSi1mzpl+k9ty6+Rfvxx+Q1jtXn51rUvAaz77BFmiXHfC9mZlKORgWSLOqm7MameCV9lQfNuL7UR
Z0KL48L9J5yimwCsjd9dDbjCGh1hA2UX6Q+Tuv1uni7p22GhO2EOflzBbSY25RdFxmPfk8ZtLtd8
OkA89HJxUyZO7pGVNi1kqmQB3YbpHV6UrbR9svoHGTVz7Zz+n5CCIYHVZhfBpFDU4sNE31FGhPRH
2isNOPLZYee8gAzRUxaB9UOiqVWvvOBAK0c1sFk1SSfEYSj89kPVLRa6umoogdHmjvOROzKDbkbY
igWvXKQvNx28UaO9ebST1Fs5mgYPhXKHjij+QOtCpTH6ZLQu/EgSJo1TS53aGcfaY0yxhpCBVYCJ
jvoBuHA3nysqzBSRY1D8SKgbhy/D4qxrRQxhxeroSBa1Y3g/AEM4SnDPw5WGkeIzeaRJpjI/ZGGi
9Pb4C4IbxiWkhpVu3aV/cKbwcfnWLCtwK1vs/eKTfs1w1iIg+vAtN+lvlTeFUvZk0OcYNUBmq64N
rFy7fToDZj5LQSTK5gc/9TWQHfV7chFE2dvm7qHIHc3LWt3SnPbB6pEoXWKAxNTfUgh55XJGhMLp
cSYlHPzSKtEhNvtz4DIJlna9SSup2CBLZ4QCh+d03+ACdcNqBBF/Jj2hP4NPHQRLOcgptJoM+HzK
wDanBLqGpIXT68i7iov0Tw9XxGW3TQ6zk1j9opFIYOf9y0o69jjF1b25eSUVlAVlmnnFObNy4u5D
n83GfxfUJPV4SNBgTYRQQ/X4j3MZlJIF0psbplfMKpTJLMNJvp7G3SVAJWo9zrWQGG07hBSx6Mpf
hP03/UhkM0j7t8MfK+IZaFpi/drpLBXYzZqGjw521pIHw1b0siYVa5N67Mz1X2vPa+ppEXamvdHv
6wJdV2VNu3Cb6h9Qru5ljZ10Hk4ObTCZb6qlSZGorW/RrFA/YstgDMfuuZ0QFLJbk8dlTdUvd5xa
9sK7rmh7KrCxuQG5153fxXPJd7ZR6qUnKsVP83B36iXJTWvwK89RL48A8kSub42ZywwqqzTR5Kt7
qzNTZgKXNApBkU1QKl2nt6IKitFGiNwM1wlJLXskHneYbDQC1TBgeKtyj6Dx3bguL6Kmr0w0QEqZ
cPQKuCcl+JQu4r0Lbbkf0i1pULIz9KTLV6WBocAbmBV/nW0a1ocoSP6HJuuqRPfVwB2L8rvJfc9H
wKlgI5QlxrfvuzQXHxU5t6R+bjddqCW963g4/8eoR+lmzTfABZlmS1MkgqQwTnib6XfpVS7HBNo1
RzElaCrt2AmT9UZcj02uO2xX4hQTiDiQ2g1sNetjykCIieuJoPgirGTqvX1Y7ulUKv/2H1eneItV
/5Pw5qW9B2KhlVOLNIGkW6FqMPoEzaC1lYWXYPnw76fd/gre8C+qUyd8TNYqjcQ/2km60w15IMjB
TDs+sMA6w6JQiiDQghQu8RPWWF3daQGB9Nln1uOIxa4OrCVNNL5Cx3jqdyW0Iq+x42XaMpsq04Kr
eNBong4nd/gj6ItLN3MYGcQ2qETllbpIx3FJSvbFlY0y6GOOer3dQC2NkVncd2eo+o9zSqJnoUtf
sxZzr2gjiJ1ecdOl0z0l8e8REKzq2ySs6ia99sf9TlADjy2tx7t7MjEHFl6FrLepEuS9eM7hhGz0
1lWyTylomobwitkgbe3J9VaAzTGPDXp2B83VzV6CNkHQEB3CbHqDQ6JGL2l3hjlaP/pa/xgyBZWu
YS4iHlZdIk66aXcUqmCpGvHUnnsEnndWaRLYIsCbR8Wi6obPOKiM/2oV9xuzAUFfYosoJB8njbkk
RE8DNju5jSuJPrIy5lmbGkIIpZXYlTCELBzwCyrPjPw7HbkkH8QkihkIb8memTFsZEmtldOQ06JP
89/lxG8cR4pSL2YTWa+wPBVcC/ZORbbRQvkI9jmxzf9x6WiapZ0PCXD/ZgOZ9tkk1AH7HxfYNHF+
ubXBeQaj2Et/mdc03Ln3Lx0741Ogzk9PzwUx6GFsC7wcRPUP//M14RoQpDFW1ErrWtbXTThbRvfT
feAys6exLz8SuhSjJFN9DQZet/GSD6xvhqWKnDxVvD6YeTPMYExYR1yjzXU3bfpuapOfOMz7laDP
pFjQHYO2et+teseJscbrP3Sm/3g9gmgl+H5sb6r27eTJdC4LSEUVc/c1F89RMoefIrPMawiqenuD
3HT0NCceOJguN+cTKv+jaH5bjrBZHvuNDGissu6GfuJM+Gv8b85u9JOeAs3iKSu69+iAFh6Sp9vH
73FDC/hMvJge9TifJtwvsUphxQXipkcUUpTKBfwhoMHSmQVFglwqrCsOZmmFbFkLMQOkwDAWuH9/
xeP1jp5eLiuiHhGh/FgVus6pezIbN1VjgFjs6BQp8nsvVDwUqFKw433293U6jBUCvRycZyMVWuQN
rk+dHmRZ5HH2TcVll1v+Uek0E1DpvySeyi49qer20ufhRPUWiAgDAZ0ovyjJApR0An0/xG344fNR
gyhc4jreP82LM52hg8L6h7tmmrEN0ojCWOwV1MCtdx/is1PNTgyf6UxG/m8LnjFVIB8MBUlnrxim
iElXfwTLgHJ+4El40EpIfQ91QvsujCtVIhnjcN0q3BkHUEKDTarCndadTT0OsTzsIkPw1C5tbngw
II83sisIutccVnih8kdZnZhwp7FY7cFi1dcNeR4En/iDns7glDcZndwqhxVEBxqj51eMwkS8RzJX
kvNd5ZUjKwZwtTzt+w+zvmTImvzPEzIhJP/yhi5dHkdh3CTJCwRXfH8qT6LZPzsDXzmBj65BMTj5
MXxyTNSU/enDXHWBgxbjsndOzxZoLE98cfjgePAYJd+mTEaGghs7NTOp3URLWYFjIPffXJRcCtLE
W6zoyiRXRkfJyqVOdwnqDXcESGBb4ds+omWHBWU/DsQp9xSbVrxAehgjelH0aMgjeBiS59zhuU1O
veUNPO5lhqa9MnNBhHDmefLG8xk8RmfBEUxNvLiSuPbwRlWZKJuJ56wh0mJ0Ifi4Y0PWvr8WERp7
Ujh3lYuOBYHDVIs/B7nbCeYpGWJ9peSOC6Ijn+8fFk3ykHk2UnOnJOqkXPQIK9mOB5fjgfDsDcw7
9UMJxUHz7yZOaPUmaKpT4gjxjrN8JdW3zX09kwlkbk03tqD2pEfV4BdnTJLeeRaFO+EjntwXkl2L
99zLsNP+38/e0qCtcWG/wrmJI1E21hcYgCVnV45NamCDYeDO33+bBOtVX1zr4V0WtuHe55SzS7+J
9xr81ryQpeLOkas3L9Untzu+EybgGd786v6MOhpAppH1sVnvfQoWBfNnrM2t+BAKgDTGKwBZFbJ6
GbNYSJqmz6aP4E0vB9qU+App8jYUC9ZlzVVrU7SxTIlr6ETsYJ5NA7U6Vyig/Bn3Bj8A6y7mPQuM
7YH7Cs0qhi7iSwvCIhbk52ATVzw0+D9JY/6+mQCGGv+Gm2xq+/o1COjdNpKOJBaQYu/1thy9WiJO
a5QiDTPl06eviPxA+xNBYS16hPKXWasdXkie4Jc9EylR2RGkOQyxRLilL6zLb7y6okiKStDy6Ij9
IJ5vbGuGxYeeP0RCF1YdKybuJcCGBooEBoJE0RdqKCUz86ZFlNuT/zWnkQFi0neIa6o1dk4olzQc
lPvyvqKtMxkzGppNw+QOSq6qHeebr2x+LQ92pHENgcpb0yqOO8DnNuaukAXl6nvI7V1KV0j/1yt1
rszYdsrF+Jnbv96/ihEEVX2qestOwLLTh8jEULCpUSafCm8RV7hX+zsGSg5eilebRvhHPFOS2pVT
89/tWIDGqy/eaS2IlA894pEYbMr6qRJ4l8BRviuebrlPhsIjy43tApDZR8x5tCzi9BpcyipAL0V3
zJvVK4CZGI4qibpmzjGCdnu5WUKljlM+6vuJq/qeISTYRo2eLyRElzT27BvH2AWnjXDb43PYB1HN
trIIKYGv0+vwJR7TZSAZdAyjenQdzTijaR3Bf3m6QOoZxvLIyzE+axRsQDeyfPhUyx/N4MemWG0m
SkshHQIi2wJeyXGLpmGXj+v8fIgnCYfzfsCBnFsuLyxrxGQCYf87Suom2r9hDruv9QEtglkg0S2q
cS+JRWwMb0NdhXphl2Xga+JWPTnxUwQjm21W5tKimhp+u+uRBO3+jEymQz9ucKWFqSBA66X+/xXq
JcQFTaomxm+ubOqgAXk8eNea3BDQMwpPfXwKxQbsXMFdViZ0WfIkiBvu2pLtbVc8URJvGyq/1jlo
F/s3HeZZpjpPH5Vx85qob+UpQjmXtuRyTN9LDYu61zH/4dh6Ui+bu5GW8EUtayhmir861FL9JZp9
UT4qxXNDP43o6YXifzpKnjyjbkwiiJMhIhqL5FvrgrD4h5w6wAwDJSwGs0pGg0DFVHDeEnGjz3E/
kGb3VLkm4hv3zIrg0YgKbOVEAMUO/w7TsFwpj/16QK4DzjKvnP/+a86sf4hRGESz3d7AQNW5nyLN
OnXobX8cvM1MR2yxWgX6LlKGyq+HVNB9sG5lToWlHmEcwaFqVTcIXOdPdGuw7qfxph7vaTw1fQ6A
pMarSCsW9rH86ItmllY1vFeKMMgSDKK+PysJuiaCmi+BiiAX6TJmzIQJiLCsbp4/qNj9lGUDTqB2
7q5TqZyT/HsvxPuz02ey3+gYWHNkbVP43XKomNtmgD3WCRBugWAR0eY0ZzF+tjjjbV+pHJczO6oe
lPGZ/RsVu5qvNdV5T7s0rJvUDyVWyXX91bFqwKGuNc7/LhE8ZmjSuVRxd6sxwZooD0CQ8l3OJhII
D2XdRNgVWT36MvnbfIRNqqQgEeCbijr8drgYfpp8e8wjuT3pxLMBE6ptRvOg+Spjo6GWcZW6dtdO
r3YG+lh7hRBzVO2+KxqiC/3jR4UTAnl3GQ2P2vsG8XvG5Hy0+oFvyFjLLYqQ0GQuDlSVk/4rpZML
4zmTz8OycD8qnm+G61nSNsH0SiCCWj+QheINJox62cDpUwLKohlyCR6og1H22FhkD/GpliDXvBL3
T+dRzVm0Cwsk2TdEYJnAmvVP9bwb3RC2snu/YTw/J99wSPS/RDIKDHTCHlAC92L+AtY3oO56a88k
cVZj0qpddI9nfUjDe+lb8kDMfzcqsRHj6NTcT9j1MzT+AgZJgfge5ThdnvyYxvMeXdepnhIGnPHi
orVZvJ07Mz/DJAAKLSRfL9WaWnoGAooZrvPL5GQWoLcOb2sBi5uhr7TuUi1TCyvbONOsVPYvtU19
lOkRAU2zGOHd9gPHt3IK4+FpHK6LyVYkaE46slAkP+hIVzYQR9nFFss658PPJ58nENPcngXriYdU
m0Z8FE8bNyW49lB8/XmpGi+NO27GwPKM/PYgbAqG5knM/+Gohy+DgLDqFh0AKYwaDsqUQoEmKf0a
3Bf+zj4sLRa8/uRfyfxlKXXeTVp12FgAIGiMoCQvWwKLpmTanNerPdVa6R/X2t4yjlrwaONwYy6p
SallVug8U/7LokzUajBkrzDtpNgw+6lKD6ho/OZCczz76xQPxOcsCx0X1/3NRW64mCIfqtIULPS8
d4gvNiVX3gDFiFIQx5lCc+oJYCor2cOY+u9WXhnjtcp/YMdv3rtjjBsJregij5wtrGbWflVy0JQu
7JHxufRI+hYHmwMIi1DkoeDzlzHacLUZLpBfsJqDZ1E0a2xhjujduLNdeFNg2LaOI7zOSbCCX0FD
2W0YpwfhNiXgMsfY6xYEvnkW6dxcAx9qlxGJb1Qw3asLlfrViwHatUs8aYcnuugUiA7mGlWIpb1R
zoi/3wwc20PJLH5W+NFWhMOc8ipM85b8o8aslJ5DE0+NVxrZIsu3kvk/+Bt5v1nmb/XhobDna6M4
WHk7hVqEyaSUJCo1PvUgPhPijCapxKVfq0Dr+0hOfOYmmC3oJtT3ktXFRoM/UWN0gSJOQKUyf9UN
ODpSVuFRowOuV9Od82RPB3u1WhyNCCGF32jNuQg3ayHOyb2Ub34oM8P2gYVIxC92U8Etghg8Zikd
pF1lrALzkmzVf+zLyXxb7pqiqKxB2cNMbyQpSe49lntk/SIgrOhKbVyWOfZzhhiquyeR7cEPKlVX
WuHISLiocjg5xKMg7Y07bJIOAVlvTVZj9q2xvhR7lkUC43dTNHKAuKJAOFHfmG8JJ5cRVzoFO6x/
QbtJ0brbJqt9NQZz5/P3pvYjivuwyCx4p9Xqr3CbWo3riH9kuUQB70kJTf8YDpSCq9uwyJoqTfLJ
mcBE6x/sitNw2DMlm/syM8bG3AJh71ZfBqaHshYs7pq2ixdzVVtTsAILAy0ftwryw9eHEBzdResP
ymP9lSNVKrke0OPpn6YP9FdOrsXEEKOphJTUzX9bmTbR685dZm7VdbeRzTdvKJ+gUp2Q9TKprU4K
4GSzBjcmDlwauW5vNnhF2k7IDi+A51uFh9gD2goVEMVMmtEkMeXKBlD0/ZgE3q4PTg4PjMcZhv28
/9Up2yc8Lv/gfi5YU1mXDRkV1pO8bFAEzQqVA4Ub3q8+T06GkZ+fPJycJDKfbfHoIXxGcgASIr6Z
4pLlCBoxP8Yj8yTJWvaewZ3tjwppWG4Clc6Fe8uObRx8juT755+X28nd8Vppx3XQRvDBhU+1atQA
YZnXCF9YzJmbNmcWVXbJ3SF238LQD4rrgPLeu/T4TnnKjFo8yWPIVoTFTHQEWTKJebnHqwGJKSc/
jWFLifRDj9NKK5XQbEEB3i2+tf/phaRVt7Pa25ATxLCsWrINR+/t6OLJuutKky3NruFXcCXnMhwz
Ap2Ca0yEZHyPgSJicx4PS8Bh0Z2ZZZ5Jkhd/y/bHTRW0By8ovIpXGQTJBaeWEQbhEtUdu9izPxI2
JmybQeuGmsFx5UUT4csESsirO4idhM5YVTu6hc8HemLc+A4P2kXDnGFSPv5f6hb4OQyouJE8nKRR
aGnvu2PLoChezPpyTngPPafaHwnjAh/jxb6GULGEYDby+61M8AojzWBPErhQRBXl5NCUt5YOOAOo
noVvdXAm63F7tapjEmQ9nuAcsdsxso3FHcPFIYat9eohCdSqHhDaE4Liw5F57WL3vymo9kjwOk8x
CFb6SwSaxN+++lVg/RMlzZ+75Uf5g9AEBnxqPGOAK6cSmHuyNwBiKCAxgj9iZnusRgkeJGrmA5fz
uZs39cSaet2n1+VNJs+EoVqiiJVJDFugaE5rYCGygjkjE8ya9GZjoo5uam1TNdW5wesvpgtkcMBz
mHQ6BCt+Ob7Zuf4005ZwO6oCsScVlrlsYKb4pj3LAFTwFGDj0YCWOnz0X+fsvVaeb6zIpEtAV6m1
nS5ZTEEUgoGu1Mz6+C8fAg6HQ99ysyD4o7Y9SSUwrzDHdciOgZvjIluR8udMaH3pVVzpLkTtMcHi
H2zlNHObzrdf82apPKAKnoyKDbDnTodjsswFd76aa4PxDny5mh7xPoRlQ0KGEBDXr/J8G02z6lNY
3M9ZID9ctOeIHrq+fNMZJjCuGFAS71vnwoNDp1Ykzrr2RIKnUvsIfvNhBbmM7UpNCJvdlbQMC1vg
pP6kzRkj33KkCQFrE5RMO5ZvwnCEQZXB82TAvSTCiM5MzMSB508pH9ObHwTi0CxpRRMEeYNx59bI
qKQzPewQ8rk5jQLqj5O71c8jM3KBaiD3MsxLKX5kfG5w/U7BvCcEUyVRr7UR+rrvxnMsNCD0Gb6T
22Ky17Vjm+jPAi/6sMDEuJfaS/u14TrqekAgaWLG4u7XD48ySugHrwMEaDvqRBWG2guRUVH5WWWR
E5bIFIrtoUqafRdrOaTjyBM0uJGk7ZxLoNP9GEA7C1+7oF2575NJqQYodLo2QjFIHcv/prXv/pc5
P1kD2JSooJUPrYhBHRNm3ZDvocAMl8USRNEVZt1TmBp8AbhrjtisEHm+XZ5oe6ckREoHNDn9Ca13
ciJcydX+ccvx67jyy2GANIY+JVr9XZCrY7P8w1JF/wT7Eg9NBKg9rww6X4JGZow/yVIEN6O1SnFV
Lfv4Lns1DDNWrN7iwtOJGUDVtk2UxkgVjkYjVSgyvGVR0GYvS3mrCrUIaynl/K+Cd5tv+Gvj+fUG
qy399to93UOVu9HfHAxiNW/ONINh3+/ufO6YEmFyd7OOP/CviJCBoAOpWSsZihMyeKw/75YQ7WCR
/LAFD5XDQ6RTGKxEhicSnvh6hZu+mQYkUd8f0zEOMaL1XCTFvGix5h7tG6qR/lmSg9J1S08/cglg
aWf1M43N/TQxaaQpZCiuLqUudvOoChr0GhfXL3SS8QHrdn9UOnv+BYH6yr0eWwOmhE63wLTMi0g2
pzxwV9FdNOGmX4sN9xHvg/gmd0IF5rIpWX6QbbF61wdl9M1qwarXGgSQECdgzMl5zF0sS/OzQd5B
pXzrD9xhnoXg/OdSeXI5HaAtPDJJZzbUfqUFcM6KrL+A3WmhBBV80lWqEdvcIZq7UXgScywDCqE1
BanbIru866O/7yiPY4ZhgTiuQmqDfc/P8bUVaSSQPydPjHDB1UEK1WoHV6gUkBQuIMA1O0SVWNf7
X2unQc4ZYZbIk8sWarjLmlWw7DZM8MWzPzDMSB8B4lmkHqAT5pJZnnnZ0no/29BQPym8r90KysUq
++GCqk5R2mgXUKMRA4dUE9s/A8iVoCglFySXplL+J+vzUldUUe1sNOo0ICvC+C+fXtlnx6FH+B2k
1IyrYZgWRk42HPwr7ZNp1zu5WlphZA0IAQnNsTXS9+1W1azMa6ihyYjs7D3m7696dC+q2UD+QV03
QKKhsxl1Dpw017XETvZah5W6k2bnRBamv6KcATQzBh4iF8/6FEVh7s5KX5w1qw6O+b903OMlFIG5
t8t7VXznL2rI8De/34u2YkXG9uOfbFnrU8fDWhPbONU/5mYypyOaqre0yQw+jcPj4dIV1YiDaZFH
qi/m+NHYAJaMdnIYFiYR5B9NwmByigs2RuObxON3wqtgM43RqdkBfmlbkQbHONrNRAPK+bYRweQ/
mCfHh0z6IEmF2RCTdTNYLKXWa1r9hbwIgOBez8jfVQ18vNIiOHTJVfyD3OG57pGZjJt/9bKzLKed
uXbiMlowWoj6BJ/o/g0432aNj+xgcfNpJGNX9G8P4jNBnxLkVM6LL+7Jv/JAIqQEqkOKs7ErZNq5
pmSS7EJ8KEYT4Pp7YztU+xgss4W0EVo0SgHJs1bBaF3SBszaM5ILA7v9M6nFp6q+Gn9pB1E+LA9o
bM0vfk09aa4xQTz+fVMVcEe0kn1VFb1ixurJ+1n7VTTDMV7jgx2/4gWyj9KhWz/cSeRTzyVIYxMA
Z8hKyAqkObQbeu8e3rtkYPqO3nA6k4HzSqWyZbp375YAoXFXcwW+PTG+stbeeRtTtsJzCx0oplKP
wzDziNC047JYC125gNPn5puEm5hjArCUNP5YVxE8YdyER00mc15rKsScnLVNsJE6BJDEwZCAG8Co
9RsUNsq3mavMwBisA5YC+0Gq6MBmFb+rUGpc/xyTf0H96qwXWjX0VW9ggd2aZeZ7CqAgWD/xfwwh
4G8WfRyeVjVYJgL1H2muK1r6zxtbdjeYRtQ5cIdijeSXLP40LdCpezgqFJq1Dqsqvss3TEyIykeV
GJpAgBsED//dJgkNHR6IPz9x3BPmFnhIv1jUTkZ58X7gYiUuf/rnsWbxqMp9oEv/SfkU+lQ8/fJe
Tk/AOfCVMbhu9X71yyPkESmWy4F8DzVNzc7LUQ51hgBksWwxVkVfRGZgAYBUDS7109rkDR/Sz1kK
hN5Sn9b2CJ11AgsYASRS4Pn5Q+qeNhCUOVr5ztGREVaQd7NWkiC+G/wLaVyw64ByLv3E12wHyWxt
ObtSPl2SM6QWJcZmgQ7tu6DAG9VYHCgDyvI7Z4Hc78189+S5bQcyxo4KKioWKc3hOlr2rhD5XJ0C
7lVyVM3fTF78Vf0oZbupc6xh/dZAtSTBYauIX+1ksbKcqKXbU+kEzb7GW1WODjIHQ63uztqqbaH/
Bo8o1W7mY0SBpIfm/ThNMgyNcVUZc9Q0iGkTAyLsriTSNliap4NOF1bKZlqfwBfo6RkUfgNnvtVF
Z3S3J+FMeGJ0QCEO/QrNlaQuhWoXxN9QHt8Ecx7xJ+a/qY2ShaST2MlF/YcAwOwx/kwpXiBDX4Jo
nzNNQZLgaPRD+eNH06atnJ1GulyrLgkHu0jUTTj/QErxzplhE3YR5uI/M2u5Id2OsxRYsHfteNwG
v/EOj0jD/3WW0oqcvzaUKX6gJBK5h/RedVyYCN7XmVOwUgUyuUPFBkBxpmoG6xJZsKiWxtphj0pI
V/PbgUB0/g/4XOmehA1ahazSW7AldUQmWZKfgLa6hRdPGwX2UoqffGSaapf+sccV2Mwcz7/seYck
TJQHPe5qwd/21u8X755ggaVv1ydT2maogET+qmMxXeOTwUQIf8o/R5WeM9FcHg1VUPZLEyeUKZWH
FjC6NcPVDBJX5l8oJS8Q5kCe/KIEoxz39H9kna3BA/SkxKAUx8Sw5a2NMwpP6vYbWZg6e9841Hos
WUuu72oiF3QWmWzUdhoLl3nX0Rj+/Gx7QBujlxYZwdzdbbmiLSLbBkGvNS6pbQRtSCS4WRl8KHHO
jKt3tohSAm1B2vm93HBGGu0OY6Fpt+BF+qsGDRXQd1GOYF7zFA7m5GvjDaEXC35beGDpVydnj/Ax
lNyqCME4Hiji1Q8448+LPWmiuOEbCRRP9xDWfN6GVvbeBPYqxLHung92GYnSkY3aIgPzZJd/1BjK
gDlWIZmCAtIA/KsEFc5iNlX6eBqobpWx6vt2cKd6yFMm0kAvxyHuskVdKTz7vLsVzhfq9yjSTi+2
cKc9usgamA1e4f2KO8SFAohsFvUeO8pbwAuOeOc05592ZerfHGiMK2DV64LyeILrZt5NrKM6IGaH
k2JdoxeuTET6BVr+v9Nn7hY19gXfoGDLK0qjYg7THvSWWtvuiwugu5lBmLP1PsxS7wvdFWB9a2m4
hDi4kOqlPWPQSVERd/PIqDYdDxCCzzr0+xxYYcdq9sRspr8m8rYbYigsLsii7hlmtxBeV3iHQFNA
CU7AZTSPqobwvZBQ6Q8Z+gFb+g5gpWT8uV9IizG3IvuMWtkdJR9zWZZtyjP/tL7ZXqtt63QXnZDL
7s4R+GSPU8mwRFwsjXwgn4fhlvgONuyEr5yK+tMgeS7EVbg5sEagE+VgvqMctEcjlc/LkudYJWMy
qzWQv4agcgYtVggfo/+JSafabxQfptjacDdvQyJDCgBjHdSuzTUKDs640illBEUEAPtGPFNkUxsY
+v/vn/6i4JkxWYgyyY8BUq4bhcgVmO/IfsFYx4SodGBL/v8jf+jqoeFB56xgL7tJF7hca7j3Q7gy
0a5NbyNYCqatE8AVNEahvkdQZkXvLjUNEjU0+v6KxxwJIOVq7BdqIMq2rg09s1iWzs1H+IW8QRLl
/zqulKncg0VIk6p9lZRrg+zWB4WzhvXQrsWyGx0o9VW8w/AGM1yi7CpGxV1CKIivFR197mkuiqOD
fAwJCnW6QAR4aqQxOojdT+qRBcZStutLUe8Ijr53JaNd2Qj6zRndsJFUfbASiFW63OjDmYTKQsrW
oNsipZsvQ4sgIS1vraPc7WB0VVUw3xCnwz4U4OGZqnXAfryXc30Uzx8W5kZtUeKiUkwyuSFcpuay
L22Pu938xMbCwyD1MZzqWTmoPaM72BLFontWCWYVmKbz11KZeXKzF7B+Iv10AUqLA/bCVHPTSh/B
DciSuFBTzP65L7Cwvwh/OMdC62TErTiydGJB0JzMvOF4nGJD3rKb6M+cdT63MPQNDehtrvUpqp7e
8cXmR9qB+nkXW45nQqID8R7YAeJWRufYl5qgaVGyeGu2iirNCBOa3jioY61cWyfZz7Pd+lLevobW
sY/+AzTCTNG3mu8XiJYNvbhGx9gU+MgPuMaHYl1cec67Yy4/wRRqo2JdGER6bxLstt28hICgI2Gl
0TbpkvUnzmLALlw6ZLpAZ03cYWjLLFQ7LnLp7mVwOH79oFEmDncwMoo6qri+A+hmbIqiMjhjJ/BB
uKyhnzcnpJZcMdCB9F5sK/AvYA4MBf6WAxgm0tezo/R12L9KA/Ma02zPBAU3RZNnJn70zMKaHb+e
03j/HieaJMRr/8uJ4nGYuLvSv3uHryu3czmedgHH4/7VRFYKrgpmTVig2b0WsWz76GorH61iiLf2
CqmayNysJRXboVMfjlVAq2UX48K987U3tWs+qvpScm/Mung3To8AS0Y6cRHop8wkOQNR/DyD6+Gr
Po9olwVyvA3axsJkNq1nyRkNTwbwAIWEIrieKKZKDIMoI5bmiPMzlLonGKnD0ZIHXu21bA+GIu5n
ltki4tF54J8/vdKKRhIHEZqsqqCSuncsoo2XtMSKIMOhRuT2zqRFj/Tn2+WkQBlbST7n1qeg56lZ
3HMpP9H1fs7Rko0mXQx2cAUqnBBBqyLbSfwj3pTWPkMb6TgORTOroWMNcWdZRiKHyQmN4gR0W56h
8aTD38eJSPvJRMbN/vvzDo1ZoJpjHVWkj5dF35HomeE7bnywQqx32/1Deiro02YBDGf7p5fntL3I
Qffth6orPoZBNPD+Qy2Kno//0aMWzlEodAg+SrHq/dF7qpWspe0jdkzVOUGtIVi3M3czCCT3c4OR
U7xYkw+6MGfscPZDD2d2lVwrsUtKuHV1kvofe0TQQAzwVOSUBxIoDE0y/JXm9dJ4WKG+oRV4XpTV
sfVT8IVcU34lZBTNdTBjh5nlWMY9CTtkaYkdkNMsYq1bYCtFjKH7k/CrBO6YGksYlk+elYWQ2JjP
zw2YdO3IEyz4x8twMk1/6Dlj87e0EI/fYJubRMZWZiImB8eMFW/iw5MPj3ln2Z6zHwD2l+jJHYzz
l0dwn15GzFw/NlB3QAgUSPuxrhkpcYYVAvBR3qCWsA6xYJMEfKbzFCmREw5irKdwAfPpnNQTS/dz
uC/UbVos7nT91r/UX19l3ZOoQIytAeLxNlgRn8aDihaawhIIDO61LHz1/OX9rIJVXMHkSs4sbc1P
kqnHVHFp/W0RZWIWgGFhyX3nWpr7nm43C/G6QQBdnCOCSqqfPCX33ZQHUpkpaTndjLLRyVKvL1Ku
m8Y4FrJzUd4qI/3YL13uC7u9KM4OcC1e0Fd/LJ5FdpY6IaPBylTAekzNVZ2cNk035WFQ18cpxymx
lDTrzYUSFmv9hyTNMdS5EURro29d1Cxy4tvcBT3LwGT9ReWIbWKULLWay+A04YvZGH7wE2THMEPE
UxqohryD1BBFkiWG7aF5RfGxF6RVTxK//CwJAZqFexOAUQkxIhWNX3GQZB7iXUOyxRaYTE+HQ7LW
O3re7gZe72mpL2OT0VNmAK6S7/u0IZCl95QS8UNfbeEWOOEHd328KHzo9sjNOdmb588Xm0IHmDjk
ieHtMxXRhGcJSpsoDRJnIa2Uzakl+PHsJOmd6AIk/pE/7CC8h9Jz34Q91Z78UpL44A29XOkGZULC
kr1Kai4pQ3NfUGTpHV8dksC3Lvdrnr7n7T2Kbkcn8l6toXKjDa7+E2QZ0oGM6NRmurEcfI64+gJJ
R+5J/fAZyZF8n5nd+EQYfljkg28LhBcwtdbd5f2bAgZ7a5dko2jVOvbiWB2LPmgk2hwbnDOJaWoI
HFTbvhJvhDEW+BQ+Ts6aYWWXpxSFnUwhFmkQ0YDj8Dmx4LAFazEetilL5Smxi275RCQQ86V1CWag
F9BDnab1uae1kp55fo3pi9zBTDAox0u60xfzwMDZxF2TFFIxpaGusytbOl65Lo/OAcwAperBP2TQ
9eCmyDVAjqoyYeSNgnfi5W84bN3aysZt07Vra6JjIzE/vGeUvlx4gO0aUGw4YfU5TchketW00YyZ
B3csoAu1uIC7XscKqgXpjuo20ESr9vywjkDseCnC5Z6Y1E+STTlvuuQMngaoUPLsGKbltiD9On7I
ubfxpnzZ3n+OZTCt3jF4Fnl9facan3t7Xmhv33m/nxNMJ757fkz50RPaCcKY6RlgphQQoGqlqSj7
sRyvBEgtE8NeQrmO2E0Qq6eTVbIy28OT1Tyj9AHMnBBIuwiOLKGQXuT7chcd0v4p5gagevPJgp8Z
V+g13EfkC48k+JheleI9ElDhokRA6qwWlCZLOAWidDBW7y7132h5McSf3Z3KDBpXgnfwgw21MiNv
Icx2/PaQTJx5EhJ+emvr4ZjBiNmlV9acAlFFE5gOABUaN8zpUQpi4tS77Xg/evIVpt2TL2h9J+mu
9H5TISJI1K/CEd0Rs6cydI6lH+vyHX4NQJ2G8+TWWfSeK4WFsgqwbJioJE0gu//a2gD8v/NJvfUB
AXNcKmNBDne+bJZsTGplXfD+ViNBgnMyU9B8DLxYl6ka2jRJ9QQKhMFXOCY1TAQH8v40H+dT4EQu
S2WHJatm3jiLlwNcQWX6Vi1KwNoFarssPnKLOyjLMDR3jXZIfTQHt6wlEQYmcL/PoJjWliAMUY3q
HakGFyo+IyBfDlaGCzA9C3CZ4VuCGuOM66MrwxXXq/q2EcMlE4lnSCnjuI/a2lGRHQ8PwWgDi+cw
MSc4MLeMrSy4xnQbyoEpuu1LLXe0ndw3BHOPJcAEPn/YcvyEc4E1dxZpymm4T/zI+JcTD4lPyric
kbdwNUB/GlcaMztfNm9VODh6aw5Q4IR2sI0hwm108HJ5aZVn2a1TJUvRTtY2LPpxaIKWxHlKmEwd
N8weyY7SLl7S72YChUP2Bt5pdsFFjoE1/6R2JFgNfxnfvpmiHbcFonhBf8PttZISRUsg6ioUIMpx
LaLVpASFKvH3XkGUVOjgdeg/XRsMOvGolnJBEXlNTFTQnRYfTCiyvnXYUN2AcYk1kEqGKrMTKG8b
qVCZo+yhB61JRG9kWIOCN5SBJzpYmhfm8mIGK3VqLcvfYD6t1kRA1jsqFlKMnuQoKRuXXanZ+2JJ
9EPuAU8Q4hCLC8N26TAgTyHVmXJ17wOUpRkBVr8g4f4GgcYkHilZJVjXcUARrdwzylstMBXkZntx
UFNYwfTJkEVDFJLGkEgl7MdWz2n8PYUy+4csH3hk8hM4t9BIgp3a0vcGAPvp+HhuGSwOq/XX16c5
qzuRg+QZNEZAWT+pSaI4CfTlan0sIjZdh4OBVF2CBEQWABbyHrh/mrzV20nci397lWSkzeZ19+Ct
mChGQrAv3j0K/RiJ2cApF/FzcprsqOQugJReWv5Z0XbRDmXpa4GopLx5nGcW584xKnHt1sXDQuLp
aGJoZaoQ5MFJZ0EdHpcRqLbi7ZYjpJJSzzGZBP1ibEgVEn5+M1juMUm7HTKwkvKyXOasUlbalbDL
ggqvjOJ6VnNo1FI53mYrvTcg+gDajJKt3DipKN4QlSLNywfvynPFRPQw/iWkw0iZKZ7IfzLQzduH
UaXczWeswHC50lUep23B8p37rIa+oJI9aUmU7+4l5Nm+wDbHKFIPAWsagsmUbyaGyRfiXLpB689l
HAhK3WfKfTOEsKktCCJqs8vHdM7HyD1qCsyD1eykkJo6KKHtprUYahaOLRvzpaozNa155/xiDHmp
J55QqQU6mPanc+IY+V43VvMiHsfEv6DnbB7qf25r1C9B0yp8sEV0jwKP3kL9LNQ4kUtWnQsoQlgj
aJBdeGUDgQlgYngo/SZIee0TyZICkES73yDbZcRXt+5DFySHrlyTYx/rfNlC/z400Mv0sFgMYiJd
3uQJvAj7MN9eZ3dyaCEGQ39BA27sQB3ERFnB/1I0mGF9BVP+Z19ZscaK16XMaW3lbrBmR/n2gNOL
qXVVQdJnts0hhVQSv5wCpnwIg8xYMebkP7B4Xknuezuaphw5quHlaUi1/0JnH3oQdv1tJVyP5zDZ
StMOTW38+Z+ZhOzi1CU/wlduuu9ooFDW7UWsZRwzZO9tlUn8o6tveyA6pblfPngUpU/3tAFc1eB6
oXEFJxulTwJHRokhC4EnxEE5135xTJ5iKi3BND8Ang3VpLpRymySFBdySN/VkqA0+OBj4ulwUSgI
/5F5uzTHA04RERgkokj2xkBogqVosNWeNjSx8AgNSGlvwYcho7vhJUMDXRPqZV4A65sz2p34EZsX
CE59iKKa66YCXk1NKcrNQ6rR0qxJIyYWkhy6I6VcfdJLnHR9I5Fc8lrpp32CG7N9rWF2OwRB6ywS
3co6bLoRHo/Ixh68muBihBrppqCKH4lPzHRIqE0/u9yf6VjRudci9U4DwVQNzXbGi/Q0Ptv8hE6D
BW/YUluRtIA4h+pbtA709CVksmqFAmgA085uCD1yWXgy74XqM6UqxnF7+IicuVkPQbIfONn61bbN
xlG5ifaFbWm0nPoEwuw7VjgYb5CtIY5oeCHxcutLGAuPa/f4StPuNJW9O7OoEntYJqoKacIYi+xV
dCemmoctER5aqomk8N04B9a2Qr7zE5H3PzeObbVvVxGK+7NnT6DE0M1Zgayzl/FvVFRE1FWWK+8z
Kt9DkOQCvPllgTnDBk5qZqWl11pKHFiPYEE/HxXVBH++owHYkSLq5wwIhL4FenQaUIjXfgQo2b8m
MZAGsqz4RmoL82lETVAiEhDDkUnlU5unoWNyWt/2Vgf2PDlQ6ZwxPwQJ8+cb5jdHnt3wYPMla0Dz
VgRNxx6yjc5cDuQurZIM+IVSCHy50VBESgKD3vdNeZNJt+fsrAvpkzCS4sm9uvslGLdAowLULEfp
tqZ3whRFd+UfNUzcRjzxnbrz4NKMkoBBvsb9M7nMSEtxyjva8QrsLbWCECTXUwT66kmwAafrotud
hbjYRgX0tjkkkxiMFE+1T84BX6pw92nc+tqtCtPCtzT5TTVmghQwkw+pSgVLyjxo4dD7292XU0/2
5voHxJuf789A25KzxC2WoD5PxD5Z5uNaMxIEC4IgCCAMg8DZeEqNB9juMIVuUWO2gUyxNZe1PZ4N
C+fXqdrq4Jexa2bAxBaNviHA4+S7KhFoX4WLy9QRGyxA8SJNQfO1pAgB/FbJ5aQCPPi34+HHSVb7
Q5UfrPlL4tsTOcJJ6RME87EPci0A+r6Y6TWA0EmT0kuLCYStgvTqXTUtZAG4hEW2u6C0Gduw7qAy
Bh7V0jVH8BV5DeEgkpOv1r763q2zZJkuL6/0ReLuQEK/fJJJehjrM/HMfDUJtYqFme4BoR40MoPM
WuQ5Ef0yEELTa21AfHbvATEeNX0HvlEzQ2iOA0uHxL9LYxFz/0G4yTxlRziS+EHKVNDgAictOw4g
UzIXh3hLliNXOW9bnHBv6KXCl1RL1n+40GP+Upt9hU422XqR6XFRJqMVpJECZ0mFz1mUY/rnXZSF
ZaZTBq9PDO6rGqYgesQijHRpLvhJ3UIXdWR/LtwAbCg0YzJt7mzl2JC0szfrmv4Se0kBQNqi9+sp
DhhNL9E9I/KeD9BYfRzQA1B5bquiKdJShC3s7K2fMLQz87Vs2I3nDDgT2FNjfO7q0rZ8NCEBXF8Q
Dwom0UXsay/MGP8qBmSjpeW5pS2UUgq3NU+Qea4PTrFiDLCkUwUpm7Pe7hqkReu9P1AJY1g69Rwr
xrjXnGHKCLeyaxdezny0TzSz7jr9/yRx3ocZtkf83dxBVpEL8zyDZue4izf1XyIWWaJP9NFlIKHf
fTH6GFhTftQP9kxLWiM5W40/gCXkY11hFfuO218zehcH7d1ukH6eaJlAmUSAIEjdXddKSiEl4XNw
h4LDYgzr9Jy+7AOYWpOYj6cbNSsS4OywSEWKEhFUCUz3qFnVbmIgyEDWJtr1i5G44XEzephZrLkD
ExMbyMyXyyCwVeUBwSM8svnzzu/w3PvaOW2q7s4qce7QqSdzNx/+ebai7LRRgbYHTE0FPigs7jRD
+I4M2S0K76/0xUIBWyR8EuJo53WpThh/uNIyARl7sztPlHGs00Ev4WzqycUOgq1Vma1mZTL8TozP
pOTVAQsslEJjUaB9mebX5GA7sOy08deb7mex2lzCuHavMgyihh+Be4HquOnRUcP52o0uKgqQfVSK
it1IXj93W6Mtp0vtpG0zBaOkoWIeMJREbRpfeDbp6wHqX/WH7zad2cU5psMyUsi1NXhVJeH9BAFE
bqQmRke8fjScOrXLkIFAI0S82VKv77xzVoM0eFS86v6R65fS59Lvru9cOdjrCpdt1z+Fzhu1BhWD
a2MPkslehCZjylnhIeete4qlLMkux6jKJSW4YRqqCa4w1uZTNhJFoE2bT92SqO0dOQcJylZYgZGq
bjJgwh8MSAQsvodsUSd2eP72OG1EyLfbbZ13VJ5+nAug7DCksACxOAc+9XZTyfy51zLoxgBZd7YM
+X7r/qRE563rolwJIwwgpux1F6abjf0ltWLsrH2WqNP3U+wZFHytDIXQkkhlk18MGAIwPQUw1418
LW272/mAjfQ7I+UQAps20WTW3bJ5/HGT8lGe+mKe/WUSPc4jScNunlQIX4H5rqxGVgT788uyGBu1
NagU3eJFD8mno47WfZMgS5s+TXKQGTDRXNmcW3k2hMpknFCbjhlrN6TECndzqttxiEFCiAslc5vm
7hkQPtJYZI+Ah7GM0P4rys73MMoiMp2SntEToBiKLF2sUpWyLJifMSb5lyLxk0tHuLojxG/5qld/
CEM92WYP+WWCtlRA5utf7//ofzbcCjK0lOoc4/rrdvRO97tMQw5LtaUOXkNZti/H0D7h3i39piBf
S6fqo+bdi54ifCri4lYsX2XVLHvzwjhazbr7c70t+j9ZgQG0wNvyHLcFU6gY9KP5Fe6eAy2h2dP7
6D5DAWnRtaKwYx3ggsXMg3tjrQ/NQ/oHsFlTu/Mup6onOCHfmg/uY2xk8knPCtZ5F4cbo5HfbVKK
D/bVpee2ca4O4sXPxqkKJUiUPquKHDM9mRU4twTaWZM2WeJMj7Yj1SdvO8aMyl1ag8yyerfXG3mj
BjlQ7WAKkipJKjscrZoVkJCNwnA1B5hGUDyOYXjFvL4ttT9CzNZaKt5d+A+DBmzt+t59Hy3VU/QE
kgWxRyaYtUfqt/FBrQyPfQT1hM3TpvXHtXS59Mk/9oxDiBYyylK0BbVAMqOhLQsBrEazW4Hvdajs
MIcr1Y3r1ein7yVxh3ir8IUBgUrreVpnCD4mS3/D1APo2cct/KCXpNEzWbIrA8KZhIBfDwM6uU9f
1SkStpqOAJfl2WReKeckIFmngWUaaBYhghpz5KanV9kSzm/OFU3QaDII/U7MQkfROyQBJbbOcfan
KZPdTQqAgN4cOLHgr3lG/cLHQp7caSA0oNKEPVL10u5q/HOZFRIAwyshJqX7ZKw40lwHI+8rwfjD
8+PPy4Yw39MuQ1uH5iKBiKvColU+8BKbfHCliVKXVXVFSgMvG/LthOybEyk5AkUqQZWAfByI0GxV
uFMZKarXEsQHHqvpLHbNCuLthD+haY/wWzwv44ig1ki0iI8vCbkJ2haFGz07xFF1+dnkiIwETNlB
IXYoopchb48I6GA02dJaJWDYlFfmvpQk3dfPCISSq+XEMD9fSNU2gJFdf66Uol4F+YPFuHNnLCsu
sMqZE4ygDN59qwaIoYb3C4WmkCV7rPRfslQO5qxRZE+9JzPJcRhNKehpoIwGa+UUmC0jVdwt2A1q
OPsgJF6Od+3cQZcmcXPNxzw3yuNnYEDpLOTDJTDQfK+WSvyEbN+gzMmAKfAXM8kI9KgXg6F5WwLI
Cd3hz5LOeiXqZEGSMuRJu6rnTnsCjQJ+yLFnSsqxn5MX+AVn9CN4oYUSKlDWs0vL2DxIhEqV7nIg
HjsYaoPgz3AKKRkMZJqpTiLVaIceMG9AXDlfZyEsVUyZl2As2xhhAXPySwwY+sEaEhSBu5v725rU
vwqbMTokAWn9cHaG6HQe8H6zfyftLqXXNchtHEH64dAK63Y7XWB9hZ10Lbut6uqhAjpDBMsdz2Ko
N+RZy1WAhce3GCn1Gwv6Q4OJaffif7ZYM6Gi9juofUvNPXBQBQ3XXYbrcMkqbUIEvVMqiFcAYWb+
aesMHZc7rlDPQYu8yTbXO77G+jDuRULoQEFImwq7YhUDBEcePYqG5IuNS7tfHJIWsyrkXPg4QB7d
5TE/nH9xRWJMmY9CoWD6XWfKDQUeylITMLqqhookgtf+ac/H84cuN2nXHn4i9fd2P/wbwHTaUbRY
bxPSlSLhMDNIRhGCVQft2iEiJyoZ1lilNBfkNwSn90g9PkJWxrtC0rB+On4ujjrHDy9aSn3q0Stq
Z0CqM8ySV6heymwAY8njJAz7nVnjTDnhEIf2KeHZ/XJeOLNAssOICN6sjqjEWTHfDdoPYH9hucEY
CEJPLZX9NEmX5zN60nxRxr+vSOmaHx3v8ptRpf21jLubqM2VrrFAU48GjBRfs/fUTMR/WfkHk/fA
Sbo2LeDgVdH/xud2DSIqJqnLvfIFsF/OMwgrWaK9pwXAroNfQHvfk8JgbWIHw15Ikp2GOqRUaSMh
B/T8Wy0QrAM+SXuUQDQUP1aPNnO3sWVULubXmm2+QoQykxiXxI6zmGEsnzJR7d/easWv/qdmQQaD
IUlW1g6m/q4I8/ZJuAmge8VL9uxHyb2dwQIxK73rXPCahPQz92bl+OLVvfiJKEqxgMh9Imc/V4BF
gFz8UZt/WN44FHHCX8yHKa25zS9raNDeh7176xbHhdTFJHsXGv/kBtXUS6e0Gk5lrr51UOkbdJ7J
9Fql39abhExee0ELGke1hgGu/tkKYU594KXDJiWTn33HJSib8AApdFGg6N6f7zxviGUKOJPE1fgW
eOuRZqarN1e8xAPJK/fCHoNisIQrcDI4FZVyeNVE/4hw7ZgqGHzaCV3f7xReM+RhymVeBhsyKkLC
x5bjmNHWD7nh3FT9U5C7ukfW1xNzr2sy58acfO+NSDlZHEHwcJafWOb4uJW/pJN9nWZv3qstVJik
aX1sJBUgsAzq0ao+oUbIngwURekJRFq3C9gdhuUgoq5fitPnofuQJy8JLTtfdsf2/vwTctfh8YnA
kUM4HoS8ohdx+2cUjrckVRW5981KLPFaBuPQ05LSgE2sp1OvJIoiBBl3ABxINXGFcakt/yAkLYaC
N+0QJrL2yUqi6LhqUphUqRzUynlFhySxcSjcu2Og1LUerCnf7aqFaarxRANDrXiCoaeg9diLhUyz
julzmXLmUNyf1raBO6+XJJJCCd0c0AmoS59ik2KHMFvJ1pbHIJG1NYT/7VjnACT8t6NlnNhPfcwh
xEnmQA/WiLKg3FaeGMH+Nr612ykuOOJOS/C2KLJqNUQqPI49PooLnBUN4wySx3TsjaSvWL27L1KE
M5wNGajAIQjkiQw0fqWv+K2LpsiliTiPK6TPnVc9XTpwQpFH7pbab+5T9r1vXHfpp9+3VJWCNLFe
9DaiaiZW4Nv8UWFrI2it6UNIG43mEX8YaPtS3IQtHHs9E1RUEd8K+Acv8cF1TRownwVC5/juJQB1
pPmQVMe4NbRyIwtBgb78bu8e2or/CBCtu/qBaR7RicyIn1ZtqoVTPG7LQAq0LDvt58yEHjFza0Co
+XhqM8v6sfWAI9HG0HCWhvyQ447PCUFaHRIVVNzfyp9Wf4DJz19cbquivMuQetbYZoQylnFVbKb2
9mtWu76PJMW4LkE8lu8st0ZyoEkcmpN0tA/rS6JK5gss3LQnyUW4sg7bjXFw+Li8SOufKyZF+cpv
vasRozV9i6Ijge7Mg66qJqpkFk6iIGgkDEbubdz4vY+LYqXHxfKYiF2IzpDLxpYWfSYpAMLR1c37
6d573MSw8uy/XDRTSM97NyAW6HohzCTXDy+22Y5XSIYmJcSIDB0AUdQ6GpiRExfXOacJOsouyFzI
vQFm1ZPjmYuqjdZR0vZAzcDTf+Vc9tnNAMbgFt1CKh82srFXKsE7iNptBk8t3S4WkyKk8JunvhJ1
fcHefQn60D5UKzP2pR89fdPKMW1Xqns62SxG3e9Wzcej2ch1mSJQPWDgYUjZ1PEdVSOXloeoF6KL
vHffqkeB3a1uxnQ7zzuCduqoo18fC9t9hxzdtU1DZSbfAjxQHRBjnRG6wL1fa2lX8yaWb7ridKoG
7n0a0RPJCr96TKGkkItM5aS1CjErW+AQ8bfaWTUJi3afEiBoOjwo0habpmSP6tLcDV2tjIe5dLTG
AM1MeJijuqtE6SA6x4PvV1uqgzfmIRN600nAHFmLrYx2/Z2nKxAGhLJHNbEMvm2/9Gs6L6iXnTgm
rB/txa8PCzMmcuXT4HDEiEeaPVYwQT9TsxLtdtU1Gee0MyjG/hhmOufA8zIheWr3fVyDCRhoQ83A
I9wmSzHgKltysw3paPRmIozdg+kIU6Zqp+Gnnx+exBwAVShuzW9pvXWPCQFsJE7FPxdk1PBCRoMR
NgL43taAzlRsK84Xf0f8qNIt6IeMcxtez2AsV0lO5ML4N0K4+pj4uniXcpFNIXf9lDgznTylkMmB
UkK5mT7En9YrTUYD8ZoQqii0cfAJ7Qo0BybCrcCbcixWncGvdhLPsbrPYEv9Wc/NW9FhHpfFSUGl
u1ofmBxdG73Kv8k1tY+4Ib1OHkr79hN0ZWn0asqfwB16pYrcW3TOzTgw9tmirHaGGV/VHaiqBeTn
OzP4oPtvH4ByBBcymbo/m2V/6oluqDE2/5dpPxRi3wwuUeHjOw9TPfjDXMK5i9zspU77X2nN0ybm
9x3tUi27gZZX9UbqmmEkHTksmdPrSb7AQ5ovv2Ua0Ylchqog+I/SCepKjsG8SVLmiNe+W9bSwG8Q
aYlmlAroL7lKxFJpjtAjqYXEbh86QA2tmIBOokJEtFH9RDDVic8z/I6QzNJjttVUZLXxSrkz9tQj
JXVy5aOoZkPvp3YUrn4lG6k1hEbE81p1iAYHItFyeuJvThkpNbRwe5mNW7Y++yohZu5J0s/qhANL
eZ8DUUf6NOy8jMvNcLQEe3VBx1joFR8dkrYq/xe5jSWruPIn7LIeZVZGK5xAc8o8Vl1Tp9MeSEe6
9LDOGMvLYuiP9Pn0EgH2CdJ/XGf7mWPwBtcVfAo4VosDFdZwPv9LEQ5shOZtCxetHDKIcWJAoc6S
4owgTmxQmyMlim+g1GWHSVTSvuM4w0rwNgHAEdDVJWTv2ysgqT/KwBJfsVQot2/dKH7naQLCqfFq
o6pVbootZM+I2jgX4EmxmClGmDnG8TUoy/vZ7/dBn+L4b0xxZBF4YExJ1eQIpvPVD+I6R3ueJoFj
SUCH3KfezEr8VS0mFVTBE75q+gBjIaVZODT0X9nW5x0EhKrSA5QF6bsgPzthjmB7TnQ0JD2YHxEt
VDpDLbKcZ8BCs0rOjDtZG60MkOISf3UVXMCWoaZnvvPVHiO6Hv78xq2hexh8ToP00azjueBuRCaV
pXR5RB1uUGymbQlucjrmQKUBsZNLTGpOWZVc4uqAwComHR+wHMl9pDe9bjJQjfrh9uIN0LZ4m7J1
ypdEmzxhmaUQTMnwsV60OEEBFtSqg1dubbwemUEHcCKMGlaPfo4vvm7iUNIMito5lMTjTjcMPgOr
Qs8bPudY/sywaCa3Fx6f8cojhaSGhvwXjfs/cy3Yb5WnaACK8lCs5CwStDtTdJvd1z4R+Ur0yqPK
eQl7IaOLQpK51tZj7c0lMDa0QoIPyxwu2C1F43wWZytpmzPqRWnh5PoSvul2WDVougO25+rjxF6V
ZInHzuLuCX97JzpD3rmrQMeD6c7rVIkQKSyCGnDgHdz4xcfOUyJnTVQuqiVsV7Z37HBh6ix/tk+r
1FOlTOeTegGs4YexhBpKtPf6W9FojIyqjrgtchiVBU5lJF9FObFM4Ial4hraTe3z5axlMIEdTOon
w1YeyyuguY1UqF87Jlyg1DcrFr/IowVibBck/FLuFdxSIZoYdfQTdkIJxfcHRQo0ZByOsn2gxJV+
/oaEUY4tK+pXciQl7d4M1v8D3UrdTNbzBzbZ5rZk5KS/HUY2L7eNh9D94fBTsUflBeyfQYrKvEUr
QtAzUHFWXdNWdzxIX/nWN6y3STkEo6z17rCBVw7uXbhclxs+t2ObKJRUNvJ2qyEwpIBiEsvrcYlA
UXjHvmxyTtn0/yXWucehFZ0aZ8zJWAnb4YhceuraEg39YFKcrxks6MQ5UK2LtKeK5q4RqIFA2AfH
fsYeS4EJX/LCXUHpwmZtCIchZRurRrPLiBqClwr4hS2J7gM3wU8UTbo2H0XSVU4me37/DACS9RGM
zlauHOSMJg1jptfK9jgLJw9fbzZI+oGIDf61tRX7KUzfV/9/mFcPreoxd7HfDrL8yyM8h/JN9Qqk
gOL6rpk1iUKLIPA7BcNW8MZQOxvFynA64Ozcydwd22OCv8SfWSyfnTYCIlmeU+Ya76nNP/9JkreO
BXGysDRGoTf1jGoGUiSrxYhYlNowpEcX3iz7dJ7r7OgmJUHNH05TTWAXrkTRXFWNFPF5H55rfbJS
k0MWpP3hC9NgKAN7jG/xIi4fsDenO2/ZlHc1/GHOZ2B3W64a2NZcEGeJaruhghAXvyYved36OKIL
jegPmMSFr0KLTfTvFPDSx4oHTw89cODnCJN7DL77FE27nHCJADKAQp4w9C791epsOUpAEM0q3wZF
8oxJoAYZT+9R2wB8LBhXmmLMiDCKSITZNk7ohGw/yCw2OYbBAE1wCX2hdvfEaopn5vkJvVBuU8ax
sCwzoGEOSSsne1sFwjelvmPEJTMhOMn239RDLS/Kwr/qcxotv61lkaLJQrgLZ1IsKqxwBMMlKlak
TgMAQt+RMR92cna33KqdQ4vn/LfZi0QIiyDu5IVyNP+4MJmi+wx5whPRqaB8HVnH2J5Ec0oeq5jq
P39uLKQmDWRFP0yRx27oPlG51o+15ZI3KqIzajMxbaMNIM6hzl64cuj3eCHXeLK6H85qk6EtL6+r
B4aasHcwISBTlQvxDeZckcmiMyZffCKVG2Zn0SqOSy2bgWaRml0DodqqhHROwcAg68h9cuJSRr+D
1K3f3BJGOKRqHJexspAqhMzf/KmILdJ+jwaEvd0TFmoogtAKrSFK3v4W53rWU7nwOtDeRcwxXEm+
bodLnhE6Hws776ufLVtpjRdwvU/7IPq35mPCRV79AykvvLYVTHtEkHkwAceOa46sXgREckGgJkoC
2cOuFy7LZU8458dek3Ct5XnlK+H9yqNvPbb11k1GMYflSoCZqL3Nriaxvd/0GxuZXZ2Gib9GKrwY
Q3PBxFCMZoyKpTUmWiD4wytuMDH30BPNbPKcbDCP0T4jUort6Z2g0nC52C774/v8Z7q3ROYzKyzi
buuwSo3oEAo8Rd09JGGmRQRKyVjghUSuMHYiEpHp5eoOI2BmjpJXanTw89QKuwsmSRNN++7NaA/U
0sOtcn6/w9hUdb0MGZSIDsPMKGn9aBm04C/QiqJDA+fX9pKNiVbVVU457GdBsl1LOTKVZdd426Q2
RLeh1TAsbIdGgJGMmVEiYxB6/iRodlONXTLDABzGB1BgXuHIzh3Lg+xDlvGU1N6lEYzaLFUnAgfV
7537NRs3k0CkyO3JrEPXK2Pzs8HnU+4xTs0h+c71PmN30rAbiIOkBkyZ0mHgg4eGIOizqqbH6/uQ
wB3dlACpgXt5XZ4BFdXf8sRNwQ0UAlXzjn8+JcUyzKlToljLmAqax0fPOL2hemyAeDuFmyhrl7mK
Yy6wzJhoLwWptyiZZ6nROO8T+cIbzfWkGdTl12G1YfFOJRGgOmY68pMSB2bo9wx6b9KICcHgnI4y
p1SXxAFypX3SF2856DU3vUQdfU5kmToNdyPd/ORUFsrGp4wJUQj6EZDGeeCWPQ3RlaLmRorMI6Zh
UXA3JGEIbMXQIwcFn4DnNC/5vTVj7B+cC65Ueji5wogA9m8TyrodeSnAsZdcEWxR76Clj4xaF0F1
dkbge/XpStTUxWn5UttKbJzTt6zv6LVfCkjicIMOumcVIYJtq/hvMjCWar8I9OuIePTjKiTjEoUg
P4A2DRiAV/sjCPfwu0oHZFJ+NPFO56EBErdMbPD7FO7HHKbmObcO56StIIHbpkHITAHnm7sofuKG
9H3r6zukVfTEmOqcDqDlUtxtgXVYN2SqYBEOaNdwWHU0G5JynWfBTNoaDEucr1OkhYcucRB2uQIS
bN0w4Az2JVxsjUq7tIeYWpQ+Z1d9sJyVZOsjoLzssJW1ry+H1raANuMlEcpSvT4DJdYwNmMFwa8j
5fzUdL1rw/YI2vHal1KcX5wEOlrSoGgLViNjs9S9eJuBKFys2Gwmm+M17BtJvPjEJ+fq1HtHvHWi
QMiofsNcWf/kHIaD8hcLXyf9gH2gUKrtT1RL2Ibdr2mw22j2msbjR73EeJJVpFYsJMvsFzzMMYwk
qKpeXVUZAda6J4D3LYxB6KrnKgOIk1Zpc8Y6Bfg1Hwzrvvly1IAUBWINYrgFst7iYlt2quihkRNS
Aw3I2z4nC56cjjX3qLpJwSdI41xGDSlGrphSmGYRp3wjGCqsiNPqb7og83LNxVRwtxFv3bBgERJx
vDdP1Yvnr6ppZSeqloPNmq9s8Tz60zQd3+iOkt0q9J6t0YF6EATslzWP4eDkMh2vWd9J+6vVX7SN
Fze6Dg7V3DtWwW024t9oANuluiQGr0yK1s96WBKlx7EuKYYuXtYs66KRUZorF9TM64gorHob6u3R
2mJeaH0mUeXe0qefvJCHjhqk0FvOHBhkAxhr4d1aMKAjVenTHj76fK5pKuV8BQ3oijlcQyv98j0k
BojufdQrJdFLaqk7srE1esy0WlYO/du5cUTz2PJszbrCJbHvE6dswCNH976bWNDdprz6VeEwrP4N
qyzG3VVOv8zAJ/7I41Lo+w0jjfElV+c7Ylj+XW5M61R0qp5PJ+qjWIjH230VFl5lqR5eDH3eSpIl
jPASEwZr8J58ERg4+PGjLddLXDTGneYKG3DP1GmEw6N2QQbRbPzHGSDDQVGGm+zfyVkrnGxvCmwm
nvv5HCIIjyKcyJ9cHZuC0ryfdtI3w6UryQeEIRDvjtshDtcfK0osgrmTVrHWK1tMmo5tInK2Daoj
L5b+14Lh7ZEklxD7CXnld/GkujXwFv40cK2k+Ti6fM5uf0BeldgJWmaq6olew4mtJ9KebOp0IeF5
/I+9nm7REbwH4yNC+cCUNvYoOnevO3WLZiVmyPeOU+HjVS68nMTwlRxa8WtwuGc5WH0kFKCGrl2X
PUnQgNwpp2iTVDLGw9FTPmvocWHnRTBuEPfJSu4qyNANxierbNiAeG6kBOB1cf/ziJyGyzrtGG0h
OlVGX5O3epB0w1K5t9cnv9KVo0SLLXXT2MLAcmzEeD2ieGA/8WI4pjt8IYpPFnu+sq9bGaqGJFuR
m7yebpGChhoZFQvW5JTPtL+NMk6lFus0YBOzEfALzMEvw6di+HFoMAwhsdHUQBa9wpfR/4yAR0cM
19li9m0Ck5zlTko70kudm2doTkiwoh4s0sWNMJzefkf+FrdR/BIuLeEeN5pbpS+k5lt75cOS+q7U
2m5grdor47CcIPoqIU92E3MulFC2ejfuB7OntY6V0zFJ9jTsI6Vc9N0vu/0S4QUPC49fSSTKF2xC
zMiDNkTOvAj4n+o375P7FNSwtXV7QPn2YnQgmPaIhn0FrSXPcdamyt0QyRppfj8Kme82t2Nz5hK4
J0m6uUWf1H1GVXl8Mk9Y7qIC7zLDoleg3W6+xPbRr1eQblHUmIZX5KFo4RwRGb/kuSbKZ0EDDI+o
NuMAfc07iA1eMMEH/IKZqbiwBTdDVLmG6Ni17/4UiPlZ7z/uLNMH3Wxzq9MbMyu1zm7vZLxCw8/2
S0UIal+Xpqmh5nWfB8v/rge426LSr2ye/xEnvdp6sx/n3qxrnlwEDWTHvMi7iSlXHwKYHJ4DFIAe
skpV0apmOPuMVK1pKQLVSQaW6PXOqiAn4sVGPfo13NgaGzMJwQ86uo9r1b58Vezn1tAz3lbfpKz+
iOfNfh3rrFdlakNOEBQ1DFLQNikCbIeCj6p70+sqmQtMY6PNcmbEI3vuk+MbgwaUfg3XAMUJ21Lw
6g2ZuWz6kKpqhntYLAVklHbjEmeqog34BlKK5WDZhL+tc4v40/rR0tu+rBl0GOdWWBP1UrxJkbGo
Ip++GhnN3Fp8T510CXi/c9Qw5mahFECdF+z1cESmIy3sEw8U4l59kyN6veAT9EbbmGnNqpOII5jJ
pR+ywxK/KwTT2i3ra13We83sC6uc5BvqvQUqUP4UCJMCEq9XZQOm1iHETvy0QQM5SIqxkZJ1qo+f
g0APxILPPLWHpxFelQKL5lJR3mIcHaG6VDo8oLNCecnNHoTSz/pxfkT830PiTkKqnga2AffccFiu
xH5aiH1W4Zo4i7AQ+3C+yZRS7MLysI1b8+rW6WDvqTzyYr8y7Srqks5lEUqTbmLzUD/b76F30sso
HZTkqO0ACkwX34CpPZKssCoi39o7jVwW9YoYlmk2TQQNQKISuTopixELn2qK/1aUjB4zsWSRI1VO
HgLb8IhaKYb0b6Cg2MUfoDKCg17svMBNFPPy8Cq37GgsJrVN7pLz/hsQCVYx1dvOGouL68DjDgNp
fi1WuEIZh/kPRrbLrpZaWknJwSZG6P328DtGmJgjk1vCcKomMjdM4MVxhlqHjUkwyNzCACS1L/r8
OnKdU7Pp6ljerXvUa+jd1kSRKBThpMM7zXuBLPjWQLMMcTzSA6GlqUXVQP6lDaUgIS0uqp0e1YtA
LggKmzQvKGYXk2Hnc8fEsRjCltOivlaQjsUxN347OxemDcEF2XhcoDphO7QigMzLN3oUEwsiz4ly
smX8hDzLLtKwZpZRrQcMDFlaeDUEHGUI7Cs4DTFa2yAApiYwoLAN9o8oDN5HPSjFurWHJgSEnBNd
vM2b9af9zSn5cmqL3HdnQr+1791DgBZBzakaKb0spSHgsvtq9Xhu47uwHzD5ezhJEETda5aTbyPn
yrXMd9w/zwLXQP7n7g0bxl06oZPr9I/cCJFHYlkxjpsmjMGg9ZWXL/s/o0SSoQwM+s21neO/utOY
7SPqGWNEGLVaES+JsIQTo4HsOBbMmcKN3nJ4Y+2f6DY49Zu1GUA4wSgSOLN2FKNU97Qj1vEC9yVg
f8XBsH72+mbTv7a0nXh19c7gDIyxDrDdwKx016+ilfZlcU1qz3e4+ODWfdedxzjrajGAdEnJR+bb
/fAjLkMtdWKX19hFPyjQX08lgi3/YhAGlAGkvg3FHLnE83Dbzq7djewixDGr7NBUgyAvvRmqU/rs
ZKIHxno3CkH9+hV3/FWC5ZDohwHdpgaiF80Ubt7ZWcP1mj4QFHJU/55an1oYwVFG+UfJIPU+KSd+
KzPE337WrCvF4oYKGtGssFu5PLO6WI5bDckj4P3968LuwLPuaurfEi3i7jTnSxNSkgznPdrlO+re
26SuwPGNqsLFbQvHGhWufVEiv5z1zL3LhF3ef6ZqI8E4uvwJJ8MZYUh5590jv5no0kN0pzIOEQSn
HTRLFbqEm97Q0f6eaeTYoHyKLuu0lBhla4WB6y17deQqTtPDzH5FPTkwkpYx0RcrmhrSstauhOqp
hlixBTp+vKuba7lNdrBLstw6QNbc2z1+WSJFgIZXu7ymLhyEe5iWJm641zNayalRSans7dow+AHb
GWpfrGSIi4L5vI2YeiOwEsSqumf6RvuUSKOOERlIMqDt9owKm8/xVG9VvdZRZMzuJyd/N/5NjqM8
5/OHUbUCVadaB5vKTP9tBjaCZ/anZSRHJJ3fHtcqYx/D97JIhtOxBn+TouHvQkBN7ChFF5+NfrMF
HiNjlfGE/AM4AbyE5pHxM4y4UBYU0HEyzz1vX3buysk8KLwYdorUaWFPPPsQf/GNHNqdD5yWjJAW
xC07pvzIFUvLleJaYqOUI2Mis0p1PS6alZlxoJu9HHEFplrX2ZXJt74m1lpBX0GdAEqrDXbqTJMY
kf6Hq/6xjzEug1AP2cNGqRGfwSV3/qofwECnR9FQeO2kgn2b7yJ7K8xTEdLgpATwJwfRMOgv4p0L
NFGnboT6OQJWHz3i47mkEcpGYQPgwL6pESB/+Kl6rXM3Fg9ZJFrh5CdqhkoSBgRNyoDUV+84lMU1
lwC/L/5kg88OWLGomHN44K3LDq9Tey18TIlsY5tvDfP84cNqOOzcV+HwiyFZJFRvEtGqHdeL5nj8
L1F6IG4LooJUNWXwu9MxWrjSDNsaDBKFX11onvkQtOZ9778GkeJob1gEN92HQ8p4Olrqv2NBeNzV
Tw1wPwqpqOpz/Czvx2q+3a8axBChYviH6t8bIX8ULZxQq1T3eXczdl21kZ4i+kylswebcBzLXP2v
1RAXSaffdckOZ0XAnHpu996l93dyqrEbZqeiY5UMWG8I9As7C20nqaFvVotnIBeIgAr5YbDl2IeX
+uZZGYCbpU3ZM2+4b3J9Xj3SjWrr2ftvCs1F8HumCLA6P6c/ZVNpeb9h76NhjosadHwmmLSjWsN9
HlJNhhjFOp7btjesbGMZ7mW5ZqCytOfcWNCsY92/xtPPly9HfIyBkPi+IbZr+7eMkJkDCGmzhkx+
UQUbSfQ0NUgN/FdJ560MIf6FC26+MhRJ/SMJNpCDlP47EbXovQ4rty1JMGbSzvhbw4ZkKE5rH7g9
uMX5mI/7qAapspTKSEs2d6bGr8Iqc7+chLASM8sADrPFObLRzL77SbH4TlK7qkGBKdUelOwVgo2X
Gb+23F4mHifdoPdwl47ZEJwaG2GnBTTC/jNu4tA3gCT6ltjK0WFXJSK5+Mh+pUz5/pwOTB1vXe/x
vJDPWSSExBtZDiL+YDwzcpnrQFuPlJMZL6Qe0IsWYGdxUF/lm+PGk0X4GIyt4QJpnCgJhmwAtl7K
hW/EAG6yI5nXOddBRYW796zju2iOfQI/YQ99NYwUcQG9BDaI5SZLVYXhLQAkYWRA9FtASrelH7fa
E+GnEOgJD7M2AL1M0t8MFO9tWc/MZ3w+VxAx1xpdPD952g075JuE7+QnLgF7nxg3y7ha3jdflyRB
hr0RM5aNfjG0V5B1KEb8BYvxpdmp6sXXvZlloK2FyL82xlMNXk75k+BJcUhrfOJx/EMwnoOSVauA
okl3ddySkc1LgmjmHNLmKjtpW1Ir8H82K2XSq+LXJbzL2o7ZvIvaKbq3Gzlq9Ha+hCu7lEhxzYx6
txWYWNV8cNqWM45hteg0oXTTbP793CK108Lj220uWGzq3YaXATRzQqVvccmlzbbUOeMrvKYM7dUo
crl8ah1DSglCdC2iLsy7EI7NGW6hfFrHbMzNPPquEtDWG/ftKZxo2oWpxKMKD9tBp5N31CbZ5arg
SANnVvkvlMyysbjvCAgUcVU112W4qt36QvgXAG/1kos/3gZeICqGaoqD+sFTBoN9/NCENcU5PtFU
4cPQmgv3jcowlb1Xczo5WaawoQL4PWmWCCGvVR2I9VO2OEOqgDrm5NrCh0O4fi7fywIuCJbBfqlt
+85DX4P2lErKydwOkxFVPkJMNMG8ZzwLig5xjdmSbGcOTE44qoG7BONv47yYWibYToEdefdfr+B/
svbuvURRyD3Do/l5QIoeBZxX9Z0wsmdkaa19UhyEx/6MyqYrR+WlHPWvQz6oI7OvEMU2ZFMk474Z
Kp/UagTm41Hrj8x5Sh9JU+GAWAq0udKJpWGtmDx9a+rdVjrOIVRNdfyRpmkRHaJRl3zIEKMutNug
aWp4lU0nuR4B1r0IXuZMS+EWPs8bXj8ebjJvy9CLPrY0Ya7o1lriIHCWJgWUXuQx/KDQXG+11ZA4
ZBfVHn/PyBBtkcc3+Bok1tbJI4ZgZWNXHCxh0TMpe7p9qBzMZYGdUY2/6WCv1zvW/OtvDSuZPuCM
r4zQM3GwPVS7ChccZE5vDMueBgLvdKg/UzdR/AdkFZ66hbAitrc72Q7bCzSntvPnPL1sJmWqHMrM
pqjIPfXdK05aBzFAgDnCwylymxtmwlIF4yrNEcpBS7huJJoOjIMzNfXeWH6ZpT7USX5ZQPwVp1K4
73n9RWE9FMrigJoGIjHDX3BkJLSSbIm01ozcd16UZ4othsb4pevGAN/YaoxHNBfd0K93rstbw+br
4jiuJJaEMiXGZyIgByJ4O4kTF3Lo/SIPjSPZM/ke0PgwY3aGXOsDd9BjnPLiMRiNtiEWqJgkOMlP
6Ui9lx5sjNqUWPQ962LxvfnvRy+CFvj/oOSoPNKXOkmefkKIGDM/Kcl4UgDPuJn1JIhAC61wdFlp
Glz3N+GtwcmKFaLqwoSnGmlnMDuCnlncKAVA+KRaNYKYWgceMpPJ7wAz65Zgr1Pf3o/599Bq8nze
zFlec5yMr7bYW2TrwryKHq20WaVn0CaIVnDnQBvANIilAHJGw39WSZKr+Niw27llhEpwAFpQ9Rc4
toF5e6147t5eF2j3DWWItaea7T6ehXX61eb+/blFpUyqfQ6wUPatLVG3eVHCWhhIPuTVSa9xvrCz
tuvcPdNT/i+q73P+I5zibtCb4+HFkNpcF2yaY1KMwDETzhByrzVe1jZ8BeyFsVeLbUkzEe7lKLkt
AbvKb+xTq2cvZ6oa7IGW2yqYR2BpoouRL+YXhuVOKkuCgYp7PKWmH2t0VMc62TeuWfFd9DZ7n6cZ
UjUVBeQAoeSjKLdJ6Oe1sFKuh/ZeY/lujn5e0vyEdxW3siCKVKS3cqB8zBkTAuwJKvSESjWeBd7I
M2gQhgte+0ntyMMwVVpEFfGdnfJmKEej/D6LcyVVYwVuGP80/iZKVkxEPG9Ge4oCoa7TkNWZ9KYS
q9IKTNhrm+UHVjm1Eco1PBgR/daFkjJM1HPJL/DgsS5bJEnNF9TQxzFurOsPgibpXyjmROGcBy4e
KiRHXcvXN+De3rmOe9pzjizIxs6A7n+6cvQMnPR246WO5YdtSRAckpu5U/M9OxoIpkT29hmVdTb+
eOKS32Jq7lccv+fDNAFds2R2A9uu6IfqL8g//zX2FdvkMc6BRzat4Vd+CZaRjkzAJNPL3MbMk+aj
6OUwHeLxNwJVJP7iVJeMN/qCLTlxU8IXqRM+Z6x6cP+cdVicQBRZy2Ntm+dYN/p9YE/OicDeZr22
MDTn/9sajfBtGctniz25YkjngaEnQmneGf4HlAZq/5laojrE566DElN2Om2al3rpeaiN1OCTpPcl
L3W/5TVrqAXazJ89Gdbx8ekEahZ9ZvCN32RbNeh0Oc3SnaiJ8Yl8wKnzfkSG4SnpzMsee3JOfal9
EAvylDkAMOyuUJ2OdGJsnCfVPlOSyMwPUEq80Ar5xg0hE14KUiPZnZpeMgARpdFrF+V1tIqATxn4
5rjWKL1GVurO+nt3rRI+uQHIvDX6HJEW9SCmIPtSQOIg1IZY2xOg5+9xh5depmSqv4OqiqeUh+Uc
66d+HUYh0sPsYADO511/mrQ9zj4JBySfh9VqPxPsjHkrBAuoBhw4P8Sndmyvn2V2iLblEYw3g3K0
sWsHgTAUHX9GyMGj3isZpUKs35dZoDJmHZKjq02a2f7d2uu2RLV2C9Mq7ONtpVn/7FJmbb3DHnvo
1jqxHaXNmueUgp1ZXNQU5uuBkvzvsdr22x+vkDGmsWUMWpmT3A+Zc/Ro7DFglqwxU5wAFG1CpThl
uid4HtJBQBab2XHm5rbsgMK5YAnvQkj8z2720iR7WiiMBAGzVgKK+5VNPD4T5XUSUmIJlFWB8z0G
/leTFqRQIzlFnG+jhjgq9bBjmPw4O8MI6f4Gk1LW5ceQrBLZ2x7XsCSjKZixVTltvrmNbShOTJ7f
k7ip59jumCQRx1p9guMmF1gdqfpLz6/bmJ/UtUtIHVHaaY0aqOqsvUV+NTlVhQgBowYn5ax2EmZF
ziHPLu1MH2c2POYnQjqX7+quZ+QqBEaWf1o87PkPhT/4dsx9Tg4j146mX05oeQ+uwIaxScLoRC+5
zT7jeNIZiPTug0XiaJ5smy/gvVlajkkTqimUuMLTvcArmLavcMlMN220Thb2vQNNA5hRAJsOVnAX
vxWipYXZwq3/IjmTJ4oTn3Iap4qJK+vSUyXh8KjabA8DZtzUUkka6i7+OrhVVg9f84MClAO58Q3O
NUSqO46/LrbMgcGdMdZdwj47a+RyIAkLW5Nm2uoWBevpYPdqmaEBZoHbgCkW92CNyfcHhOboY/QZ
6Pt/NZNAsiRBMGKX7d+9IBn+1d6yFN1BE1AbmKhjX/Jce/hqfLqO/4Pwc0OUk8KvfSkbhiFHvIx6
jHKbL1QFsb9veApCpSCmdXQ46RN7sa+Dl7+G0ZUK/9WqLyzEAi4HaMLNW19rBjxw2M+p19nx1tt1
SCSiKz/S6wCWqcZGCZX02ycKSMjracjd8JsBHfnGj7T0MKRkYHGeTG52QyqoCiYhu6kD1bkb7cOr
NVJ3v16m+Mlqr1de6Z43vqlnHgl2rX6rL8nbRu9fLiqVFsxNJqKEQpwEPdajSh/S03vNdmK88Lvu
bYbejAu7/kA5suWN01sMp1DtqXu1cGTxAu5kEZGmLyTZM6mvYmyVKycZvQZ8o81yy8WmU+tUnNxc
J77UzbVTo0NNmGWXUMFswDUFjl2mgI+AUPnEvQtD4Ligm0BUVdSi/7h/VN7SwNeUXbKF8z9hngeG
PhhyouMiR9YX1RNN+WZmwHv1mBqs6uNEuRZDeAUYUKGTh1eornHmhtUJkYebirx/rk7WY+oVehBC
7JuQwN5qfZRxXBjoAvO3iaiwS2lXv/Flwl8Ot3VEg2bQ7njFfNOMKxdCk4hICAuGAk4czVt2hrl2
6NJZk9e1OxCuJdM1RZkLVjiH6uZxpwW8k08WG5B2eSGRYXzXTruCQspIJS7uPc0DUA550FU0xEKi
3X9nOcLx7Yaz5mZ5IRqfbp+vlhRiNdgECjI+6LssTrZvLyK4qhK4F+1OF1cpVjkv98h5YfDr625W
AAm2ZirvFYACqvOt3i8jQ6Fx58bnqLqnAQeace0W20FlwpmE4e8FwRQNeZVQlXJkV7OleILOZISS
4xtY+j2paLQE1JclcIvoc+GNcr06WZSeqn4eUaGt7KHOEjvs05W2kU8+mo752MuzZpAlydznuHcI
HyqKQBMmhwH3OHXZ0CgfBoxBf5K2TLp2gUioDKmm3QNT7AHoCZXICwh5v3MIBhdHJqObsvMnxvE0
W2Y1tCCk5x6mawY+hqf8PVOD98SStg1NQjwF1QuSHqze9hn62NYAkd5sZduF+QmQVklFDnkrMOHM
25OfYiW+oRadwYpFJ5RGPP3rb6zc0Fh4DGuRlZI1qcxl3gUATkfZljt4vXnXn5OR4Aq1gfYFtsGC
N53CLQPoDuT3PzAi1/nrwoR8OIpc5+RlmCauPDry4kOjSmntlbZjS4FWQLNk8OPp2O1kKkW1NROR
cez7HpUUBmbDqML/p8dQJ4gmu1SPIqqgaqeJgVzQY7ztbYQ7bw/oBP7IhAAd3G9OqhYe9wE0cxqn
ujFKbXANa9sZXDpWLCy4m28aet0f+IJ07WmA3bdHvPmiM5rDhM1WRsUMjmKfdiWw471SNU+eNpma
Ysa0IdVseGdxv/zihzXd4xW+citKccasWzg7/N5w2X1BDOfnwe8uAGmdryUm3vrrSBilc8X9hAcB
A/w0KYGwIIOmxgi0rf4ZKT58XUrAYEYtqPhrpGjTL3pMd+zphf5BP/FfO7bkr59RPqVU9f5g4BEp
B1Qp+Y2q03HnoOKJv01oiQZbVpL2+VhtAtNXUBPbtMqiUNT58BNGqiLEo82MJy1XpqsLGHRAAibs
MndaEfvgLZs5mKyZIF8AGuEUeCSgBb/K7nCu+LT/aB6i1bK121JwDmtrf4HmhSz0hwNRODWk/WGo
9mue98YM1XlX2cpBvAiBda3AA+t0moMgfpbEJYX50VpMIGdw9veF5PQ4/UM9+j+XQPC/1KM8dcM3
OpYO7aGYicFxXSmSCpgkif3ZsO24KyzBucvqm5ufDMPKrPRgIbpkt+AX+7B4A0swyyVnSkczH9vc
DmN0DByVXcf1k8QrHuwfqASeqKMFNCGc6wZQkHekopPVxiZ3FZ+QdhMB8z3ieICwyAB9LTHhXsRh
dsmDjyiPdNEZSlu0z0Opd03HpWM/ICeFaTIyfTxJM4BnePxl56VcG36Ytwrqfml5b5fu0KnklRaz
QHcWSPY+vPH7ReRu8a6MFGB45H9DvKSiGdLRWipviCXVchciVcBLWqAJzEw7ssLErqkHuKQvKAV1
ekD1teTmIvo61T7Ax/HThJCx/ZoPHZRZJFdQ9/kJkMX9nYn73zwmCLTDODHRYdBHDMYv/VeZck8g
X+J+QYnIdtsIFwImkzOjA1oN5d7Wr7v8AdBSvX1qx1D2YDDXGtQN5fnJqYUKFoWgTmJ9xyeE0U4I
x72T4qMFz852zEkiXiDrfHKIOBV3mITIJcuL/6QqObXw++zGC/vFjA6eya8gQk2xA2ZbyI5faf3O
wnn+3c4nTMcgUTeW+KHMM8naJv8JOzPLkVblh33mUXUyM4IY2GRwiS8ytrkpe1wAmew7NwHuY6JM
3zbEwoDqpQCdDH77a3X0yaR5MHqSwYhITUvlTg8E82Z0QcLQ6kvAQzOKdPhT3aZd5fSDjc6YNvr9
NJVUwKEjLL+JfxEsl80ap7lDdFBsdMWOtyrYmLedrm9wnKJlwoiNy2DNdJ/Uv21Hdl1ofR6mTZqs
ADMvCXKy/XdpfJWgbJvyLehyI2s2H+DEDKj5xlhbwWfZPzq3PUsuIftRvv8QzNdum35KG2f2jd2W
NQKeCr9JjB9PUsvG/UsuotT567jpeugtrgYrCjB7kMY9N1DzNCSgDiACbn8k3sXfv0vYVFMvdu6F
h/GMI97PFPG+HfndW4PDaP1G+gh/5VMHATnfc3V+s3GIiMLqlZQKijLU/81Es//sAi183ZaRoCGW
IimUEPpM9LC4MD2x5Bp2Ta1aK0L+ht/5pQSFNTtoj0ONJdk/w67xMLmbP7N6vZFNR8jsrBISTU3s
4tP7iJxJEqhRHB/7nfNJFvAnfobMxvbmrQpDf5J5cRQvEGRTTtXToHBgWtCgSSVBsBX+sBC2zf6z
YXwcW8U5SMPHxX84ddCz8A3QtaNyt85J45XmmVsqNZZM8CogMokwRS0tqFHFL41vGG5TkByJkf17
5+I4gCZDyFQG9E8DekFnYIiHoaKdETRM8cDdOUcBp5evFTctDJ5xVZIM1Rk3VGqsUZG4W6azN0GI
/eK5ANsA6kuosJcA3wZqFrXvzIkH9IEjA5Q8N2hTy2T+Rr46ysJxygur8V1oJnVy7bSiNVQCmDJC
YFPaV3gFl5Q51JvKUZ3eKyRCSJhZnfe4IkrO470QYZMdEeyPWJTA+HtdqWZaUckDtUO6TKag6cNr
RDbYzsiERbSGce5tQplrR293ovhNu5WObruVUOB1BP9EDCPZEpm3xtNb2C04WmLL63xcw85xkkzb
0d2HNe515IyC/1dKbFTwMVbxbbmcbimoTzcSUjTes6GcebCI829hmYdRxFcbex5iKeQ2IReEb7gI
6yaxsdfFoJ2SXJofr8IAYAy1DIlYTlHeeiujWW/SwdnqogJ+B7MJpE0p4bhMXaYppFlZf8o5qlZm
7T55irZQrhPeB2R1Gmu+rmMXFejw/IHhWIL0hTQFbNibTOSTQYELB8k4FwW/9VmDIL6eRAEIhkVo
OEQnwbAwXMbcAJEfePZRA5cn2/3lq/cgfmk2y4ahXnNXiAq9Lc+x1frJNkvZNS+g3rK3evfPeIXL
JSHPQ5uFIawHMzlPnDjhf6GJAsI6pLVWcFyqPovnisnEudIJgtF7IRH8giJjWqq0TmnzZB/Vdbqw
NjDSxPX/E+iwNvwEdgfpuk0d5kW4W0msxe39f/6ReUBo6V9McE+0c8dBTArMVJz2IQdXOKYHPpO+
16UtWQHiGZ1+qcgMDfXlOwSrOhMyh+yI70IzsWoUa0gHnx7BlZE8lgIvzi3PgV4KXZo/3xhoThVH
5luFQa8LXnD3PbfTjor2Tusleg4SJRl9DysofySWp2mj9LPqHRsHElsaHQ6SkzIY4YUF3yCQ05g8
JmK6DOE4qTZWMJakecIV60kOuWHjSDLnQO2ulHeWV9xcfyzL0Qctd8Cs5rb1Cl7DAaW23tghfNTb
NEcQaIhEhat5Q5Q2cr+560CqVKnF/gcVEbt7kSotSTtEVkdQbk8wbCOkcPQz1K52UJ/91at8IwUT
DshryHbDyWLFA0ivXE2TDGRsYPkIOTeMx6M9CRhfTmvofnBFkS0QRkY5coUlfQNQV53mNh0J5uQS
i4hKj+zJ2shLCqYUUvQAa1DQQL0ddRLF7pJA3C9ig5YvEGZxxZUN6fGZCmIPkofAE1cW8mFbJe5k
wdv6p2bWCL3/hrSJsLZt02UR7bfsndfs+MTEoo2jMKK6px7yZV7iqvIERIlkTe56OYnEXJtCCsr6
jkh6lH3CxFlfdA+5k5uXMR7sHwhlJ+GB06ByRey06+c8s9tOJt44mglH9ocgO2a4zNa5wIdwV4NY
61E/tm6jpTAxb8uRtsYQzjzPktDIMmY7v3x1oTjsPvQ7atq4D3yG7CCVRL1tchv89axNyqqhTuWW
Bt3y5hZZ+GoFHmiW0tOMPGPNKG0n9KoLAs9veLYG9R0tLnc0KoV1L6yuG7a5YAnCdGGbf5m4Zcmv
YoCNoqkOvRqoGa1ikZgurydBFTyLWGR+VbOJrqjW8HNnpSVFsk0WGMmjcygF8YJlO96utehk9vIs
SL2nGsY28y+synWIE/ZcIofW1k49ytQEjttM2VsGFiElYD0jeJ73e6eNNGtlcc0lAjfSkMPBQIuD
4vu4AoYL7kVBoE9cPnmTC8QCick6lh7X9zUsDDUKPeb4kWdJ64f9WQrX3eWnB20hCPCda31cr25n
sm6V+ZWWjeVEV26GbDoI0FJs47Vaa604VYVhzPP4B+2+/5zwKMpk7ufbcwWd0y8iIEIj5LQEz1fN
FpW25lTemveFbu/cTJ2HA73yFVXB2K2DrnkcnbAgMNbn1l0gR9cFthaGes86h7kB0JAe0ouQ7DOq
2APpC9Y5ueOLJKfr2NwRudcUPHJjzbrtqAMqHFGJnCGvofyJMivGojtK3X7xbo98ikHgNIu7BwYL
8Ezw3poOAprig4c0PiG/e+MJYKkRQKXlMYm9P7OVvfrZuBT2Np82jwm4VFFRX6POPPWyln8JVeX9
rCvdHJEixLT1QfDu8bYljNGCok1YbJ/YFivoZYxWfZ61y1RaySJHDL/i7cUkomTyssUtEtc6F6wZ
RK7qVkKcg5L6JfgETOeXqGnhNnO+bba3GoBtP1+mMTxvx9uHvYr/6BLtdI86q7kw9YQHoEZFxdEa
Rex/zCXsHxMzDne8bhzA0i7CmLkw4+eyGuuGe8eKdetcP1SPrpJX8sxh8IzuwEdp65doeFG1KvdZ
Z/21Kvtav8yNcLjRPxgstX9viPS32rEYIqALw1yw/Da5Ed1XxDQYLAORVc6mFPcCovX0aavszn7J
hJN+VHC5R3eIHENxy18RasSP2O0XTQP1J8iBMldseaL9oD3mt5gFqmhns51kDeRgVM9gBdJ6Odwx
4ctxniyuVx0VXWxIuJ+5ixpSM5CWNv3Blfj9Eg+55g255qlxevmAsYgHFEa3P809aGmlQTEJ0cgY
z0tqccOUw+hUgwc7Aqby8m+d34Q0wFSAompMEMT1zRGbEyCSqTXGSbS6qXoRBB6VNL3jl185rgPm
7V9CpSPnkaRU/gtrlPvqS0XULCmnrIprjct7m59uCpA2UJH2vViWLUmUBez19UzeljZL+U0r11TA
9O7CtdMV1Q04t3d0S7ry4gmAkDpdx019WJ7NrGMVxPh+ROkvhEtPJOhTTV5neSlEibo3PLwamv2n
Rzzg+X8o20c2P3eKH4/L3aO4UQJu5cVQfZTpYXOLw55sTfdnXcLrWlbmDSLZ0gUZ3sqRXiFcKSuy
E7Gk8SIq2wt7axVISGPvZ2fR8sNhEMpaDQ0nwiwPCXOK/xHhK5aBtqGnX3BmTNgvE7/FDMuDnYWY
pW/h4X5/b3WsNCNKPtrD+Z7yq9VhnsDV6GfGEdaRkwzM0jgjnA++a7V12s6gw12Y4LSkIzSCdnni
94IWnh20Zt87MJSE83o6DQY3D7IJQglNUeaHMewjT6hCsojKJTaAVstRgeXzXlpCavN59CZKIjTu
jU+lPLj+izgDV/wtuMy+qNTZyShCAOY9wDyLRXxFf/5Jx1EG+hcFfrq0wgsD2EEhjprVfh4ne4g7
18xf07QYe9vhyNw70ENtpIp54FIVkKdyj51ituw43hiDLBe+WmT61GHImf9ckP+5tioZ6ECNSHVn
TZ9Hbp6Vs0CoqHo6CdBbRAsiqLsgH2IPRaMl1sXKBxF61rKkM4V3ex9HSe+HVFxof9qZixTDrI2a
VbS+ZmMXeLR3FEbdGq+2lSak4la7x1uRJlkqEvodXnKmGXscNBlhQGuQ46srlC5vxAinql+hWVl9
RLd1oaMAJITx75uv12ZSJcoVsi3LS/lH66F28Tj2XFqAwt3KX8awOpo0WqqPtr38EITZHsDEY4kY
9zGjfwQ2LzG+knQ1oNKXAS1SgJ1wSTe1ePn7Rb2Uc+4qn361L5jKJRQAKzD9xFScaTLhIWichJ6G
YlCB7VoK/kzRXG1N4lp2sQuwmlLaQXpYvNKHqG0nvdFFBIhKJuqGPVHNN0Q3THEtTyeM/tpsNnV+
8gb7RFMlDAX4ovs3ulLrqaMNzy/ZIlq8MQZiS67BbPK1k16ZUuxwV3E+adG37sxqu2R0eUjkljym
DXyqVmUIzbgxJ7MB3UwdRSD2OGDioLHaMc5i88xo5sH1GN6rxGzhEC05/E8w3PJxNhdcE+YXbe+i
fUZqIalmbRVN420Ig5Ybg9omx/cfyH20TJlI0Ccfojm52JYh3kVGO5URnPnDXCdn2C6Np4FPbHGX
sDA/ywQRkJxr1gQfdvL2ljJ91L3/iB2/57oHW4feX9tYo2yHrdNoNkWdZlckKigelzUhBRhr+ghO
b8SWaPR65il/W9nATlw3WYTpi6gqT226dfoj96Xxg44P141rwT8OqVNhcmeB8qnc2XKfs3lss7qp
uJGa70yFLKBGly9ucx2h7TaKH/of07vq4Wtltd2EE1LHnvfr7d/L8deYlSdo2TACTTX2NtrrAZ1N
4laveuUM4+b8U0V5yJ3BMmtMk+7AAOYjUHFOVNML+X29BeFFbh6ic9iIC2+IuNhMaExtAQtHB96J
kjvV+vh5xOtCM5GeXTIcbsIF/aSEzdkXTz/+qHV2Md/9cROwKqnJwCKufQ6D4z4p+EYWjanDdrb5
bxEa4H3iK8bq1rPxhmafPsV9hZjCzYrXcLNn+tSNNh3CPw2DFsRLz5fsvzh7/xVqkiyCiuKOpHbt
g3bxKjZsci6hIvCpZvNgOuN2xSmEHxHgCCSRiXNpVCdEcd39KEWJVRE6D5EAodERGzA3bIp7W/GJ
zlOKph6AbGEIR7e2Hzr1wFVBNhGiVYZhIgqnZN17uhKaI7PS4uBGgkxKA2H0fxQBY/YX60Hxtk7y
r77q7KhjTWWMoy4B/Kas5sfpIYqMskHDhvXYA4a5eIjFCdXe9mn9pznby2Ctdyzwwhp8w+wVNj9c
4E1rSlXW1247Su6lLnKcPaGXc58kFpa01ttVJPJbgekz0BrByjhfuwV7MjWGd4/m+8YhRZ0yxX+G
5JMQ95cBlCqF7Y/Z7qGSDN11yV8qT2cdFDlAQyfLa8O024MGTlzqXFgn7O406rQB5dGNZw0pqThY
qMevpoaf+Rl059thtPudKRzNGZ4fuQrooaL9TkYvR7VjxF0M/6KDZKZqT+ItsEhLhSJBxT711H/r
jK4eJ693DieatiLNSbyuwjAGLoYsBMYmDkM1SSHqjbBL6eJHS/YUSuGq+xePOc0TIXUjFH1ZRjJu
GR4hgvnXU9lLSxousDeT9uWUiv4C1eW+/d3n28lHqD6d8831uTtRVo7b7xBxcRlJ569quPBsY4Ei
piYXLVXUv9d00BJOChegVl4Ylu4NihFu7R252tEaC8FEC1/RYUTmw5TpK/X6mSAiyc5sObuCBcvI
iuDdVi5mLvTe+T7oID9yLYRSjoZ4vIMZ+DEzSAXKLYIKjsOwcUGe6yXPfpGZXfT5oB4tq+CFklEt
qGZ3ulqtzFGH3T3Zqt//uxbUG6RE3jUYxYy5IrB4qru7gecaVAUR05QkJv7qFynGNlrsJBZTgzCW
K1CvvHW8hkgm3AWK1McwvwToP7lvX1CnjJzeWI+ONoF7bY7oH75BV1QWms9uxtRR/Le0APSGzVkj
oV7obALChN1bQWm7JCqA7nnEOwPaZ4RvlIwD4w/12GVPAcMJChYtHRs7Y+9murcpGmhORmPpeyH7
6X8DdklwOcZU4mMtZKUqP80KZxyFAd8AYf5JPLWCC8BxEpNPmjaPn29tVNN/5CkrM4eClxz0lVWs
b1NBvg4Vs2YkHrut1HzLqCQwNe/jaJbIpNGXwwRqqKrSGCPvJVhmwYMu53TTj+c6qqnoX8cZVbuc
EjW75hO1n7d7JDQnASg8hcq09G+Bt57WCD9Fntt4/wbAB/c/1LUxhiAAFdf8nQLG1Cm/vxW1AXeT
5oQbYIyP6a87wb+5JpfEL2KC+jcyWHQGFVDLoFzpeJIqG4D4jjoskIx+4Tk5d3bahrc30VEd4Ban
Ism5CK8pAvkRNph5+ns3HVOfrghBpG2BdIGA7AeqjBCwN6I798p8xEWh4dR8mX12Bvj02YSvOA/h
C7/5gmzCgZpYsDDgLUZ9jqWqMh6AkahXQrepOEfxMgh7wmVy/al+WzVW1MVPu7anfDXOZXFopLsO
L4T8dg2yn/9kfwEA99H3nzGIUzniJOPGRajtk9+nuuvDSfjThIdOU7SF6/j6GOv1pyHzdEjLW2Ve
4ryFA4qrqmgPjZz8LIknyDQ3Po6ecqE0Slm6LXWCeCUC0J8MBK1xsI0/itIvhQvJ0PlmkNlibd/B
52H3vo7gAYNRi8bhMOG+wn6mrlPW1P3K2fkg3pOzW5noOsWMlcKBUgk3apExTKiY3cKXrYDoD5ih
Hc7BVQqdjE4KnjmLe7e47sA1ud7Xv7v3Y4z2P3q8VWNcqIXN7krkIUvPCEp3wprbU34l9UjwiJuq
RThlLUheEPH3qf2VayxsvkPw+/+cuUm8pRYasGFkXPYYjhKSLUiCxyIAF5r3WiHow5QB9oLjh8oE
vVVKWR4bHSW/C4fRQ2NAf8dp8pHsB97NCsPEdtnoF0cvm2Apz7ElB2RS6emg9eUdeyp3Tkl5r2J8
HgaZS7OW+spuQw52OTyFyDegLvMy2nlebmPh7i7x00/bnOCPmV9eLJjRls9BeQ6TcF/jF4Ht2XJt
Gsm1vx2RGDQ8m9lMOdyWA+ZzRBXrrR19qgJhKq8q2Rm++MElpcYqnv8PDQyUgz8NEhGx9c76bVOq
6SmJveXQ51ljjvw1+bKjcNzuUKcKn0fpwZAOltmBHd9vCjaNBZgP3m4wAkdqHr3u+/UuJZIyyKsX
sjk0VEFhuD/U62SfS7K/i48gUVNKy1hdP7Ko0ij5Ce03enXvb0wNCAVinTfTnDu/LFRSZ4nkqMAP
fdX2G7UBDfuBOqRp2CQSdTLLaZda7U+eW7OshA91wtjv9HYO4IDxjPT2VPI07Q86j51oWpGh20jH
zMC+4Yg+s+VqsxdmsAR+3aZooSefBuckOEHHC39ggR8glppEMdF9NfklRjC4YjhodhViOHdLSpk5
S4SBRs4oq0dqVBXOqN/Cb3dXXr7IWI9tJ8WrtBeM8DFlCYP3W5QAOfc6io/MUEK39DEVr9lYvkmm
8GxXW4cb990iFDyeU0dKYHDQus3WOLiNgqehSmTVWGhFbM3WXiu5AYa2ARBA4AmlFsPFive9uLmT
FW8q1AxmxynA1oUz7t6GLsxd55T884BSonwXWCRQfnhjzlEdtkClTEjEjr2JI93nXdHzSTku7uPp
W+Qet+daqZ/Pit2IJYH+dit/mKUthPmTE7mahQ/0+4aos9511FKU/m0DvToCFu9l8nCWwkXW3JE6
rUWiWWsyIKugvhGKSi5Gm4jNLkhdXuRwoeYwXg60AX+ug8AKUClJiTiBehBcgkwZWgK5bVf0LJqQ
CpvZaxrUKFxkAuUDn78AlFhD1qtwn4UqwJPWEhKqa2IBtGJWVasj5/ImCdNxD+Uu7i7wzuytTBrV
zWUvhvTNj41s9SNbflmY0AGhBnHON0tropV15OZKID2hwkHS7f97Nkn4O6w/SnG31Zl6DuSfFKUv
Q+G1bZboc2r1iQWcVb/IcLnbR3FPoJJzlF7OwjbpTD7s934njQFXGap5Dq3daPmrahK7LLljHovs
m88tZqFqB5CsE6dTBgkiOESehyQW/AUXZJgq1E+iijMlCdS6V7WXBLOEnus2US5gQ+HY6o4K1w01
qh8HtN1ynYnAYeMxRhu9D7BwoEdZ6zJsI7OfgSy3zbmXLQ3xfFmBY/8PApbE4+uv0D120XZKMr+h
0Ib/FWHThjCUeLNMb39mlHTT4WBSXy6ytbfjJQqOkBzhBN0bxC8W+olrg76hFP4+cRYFs7ZpeZQh
6WZBNTjqYALZ/fJc1nXIHt0QcEEKiodv6M1ov85qzgEY53UYAtEtWK1tIlJEo3LBE0TJkkFUHRqT
H62nwxfvqvrQVo0KF1PYqjNgoD85mZnoBdXeeZApICx11Z5xT+Qzfyl2ygKKUQLiH5cBs19npmca
0MbkCz+Uaweuyrww4QGFwouNW1G7QXDsxq3pXCJhPd4HgWzim7ln3Q4aHS1t+mLNIdP+JX2HNagm
4Gn59UmJ51NJJX5Ptn3SEdtR1qJ/vcCNukydmpPZtxq3LZQvQ7E9ZrIH3jP8BQWOQjCNAO4qw/aP
lbIb7PSHwYZEHJFPBPpX7IhTq+lZH7kboA7M5kMB/q+b/TntbJLaS4uax2k3H3VSm0HZgcYpcvI5
Q+ug65xvj9c6dyCRd3KeSCqiwdL9gBrLx+HZBBKIrk0aMaDhlPvkkJfJpUNSxk+/SZObhDMqZzoQ
q5fikVJ5eqPIRlbXMq/ueCgNNNDEJ0i0GbNKcYdweGKI3CIWnIpwVaSuNe4eEmU0UbclzcMxVLJY
D4vR6wO7MYGoK/mIoVBF7LkNIMdP6Tbcx1FHOBxlFCvXlWwT5c1B4kshZ5nnJVGgQi9Ps3Q6393F
8O6V97rdD0Yq9K5TJPvOvajF/jYFod58Tun3J7uE2LiRL/3KFrwjjG/HeetQ1hDoFyTQxFLykolp
Zf8rlhqLRtkq8Pz2jUnrmwpaAM+6/RaXNdwRPI2EsFODAPVAv6IC4HgQWUKJCUUjjOwngMhFBHka
Y6e7L+8V5vjPhz/qGvTH13sprrulOozq2Ph/mXp5fAD5aLn3rIH2pyha4ZL4u4Yu1yL/e6MmQ9tp
qEqKa4jJ/6hPkrNU3YB4ok0UyxKJOne8GCherhsLKUyL6I7aCjjvFG0fHfMl4Z0haHIoG/d/Yz4N
RxHsr+ZLOIfyELFlgyhi0S1ZsyesUgpHYrHMLwGu9NkXT/rXdkoUpwdceDFJp+x1H8A/0ROKepa5
y4awD8KMfgk5/dJzR8NKjHEywBPtK/w+369Vjds9VK2kuzOuPyOdoUa2L+tRm6U95seDz0tjLrTl
7GUgJASwmGfKy8tVdovXm4xPrNmjjdJ4yKK6gUE+QF8iHBYlJCZdC+5KksmVC+MZbdRG8IMuYSH+
SvOTn8TRVqwUkbrUBOC/r8dhdeaFIHHu2EVwZUhBEUH5gjqIJml2J5T9TNrsKPRO0VvJsRO9zG0Z
HmEsNVCszztkTi9wpXvDvKmKiTHzQlJ96hUTkEmw55puWd7hH6mBh3y7FW1r8IeJRt2ms9DVDbCT
E4tVSkQ1xEH86c6+5OKVpvH7/GjuiXo/kl6ZHrbf74tFAGd7j0ZOqoyzzm6fnc71AsxKxnI9KPIH
8iSXACdUQsuYw17imLtar/CO7KTGVLNZ5iJySZ1k7s18lM9S3L6zddN952/nIDMhw9RXAT2JKQ16
KBm5b0IcJto/imT5PVFMFhMnO3iQ0uY6yLPD3SqmXg2pLxG5YqAVCRvNRwgkvIyHAW6oqJ7JGO4Y
IybSzsWj4OGERRA32xgvmDytV0FuTM/og1PmKFJ+xxVVfeKESfH7EcfMeNLvC9Ksfk97wquzVUd2
x1EHg0yYxqRQR+dV2S1oWmu9/RIDxQbn5Cv1Knyu8pqZPtR1f43xX8tQpUsllNmR9UYYGq4KumZA
7LGOQWJUFdk58QQI7XIRtd+Ci4BtGv/QsWEJFx8iT1MhAnNprajDR7ywNkuoNu5DWkV+HLB+KUi3
8zAbPGm2sdOwzLhxVA1ljNeNmrHinU58U1n1wbCN8mMxfhSAwvnHsoQYntgsgQzD5tRIb1G1rO9U
LBa78F56YBRlfbhZyhArPvB8sh9dbo9oFXLknDTmZuo/pGqy367Bm2g9QmVX9ahDlZ7AJQr2IPZu
jp6bNR5mJCksYcz27JKEHP9MscB5vhTJfpyWSahJ6md0HEq0AWvy0tKF7wEbJZe8Di2lIajcGCGJ
v/LkJ7s41FKkPbk3FbJsZcL4X+we5bkDeyyxYPL8r2a4xkcnjpLPywxJDOT6j33RgXepGaamcT/A
r8/6s6F5b+NDT1QgN6Zwwp18A053u8e1KWZfwgginhVKShL41xKF9iZfTROqvNotsYLPBiidneSA
9vjy0LO5yNuRAI+QCkoMoYQj7kK1hS0zAJBEbqHJcKd8BGkUmB6qtCY3cndLqz2w+J0BSV50pCLb
U+OHLE0GHvpEBvXeQ8qiCQMq2sObrrgZKbNFOTJu+EUzKaqoz3/WDQNl8xp0oRCoPfkeAynijQ+B
dKTn63l/PcdNYIzUSVxF1mwqJxNw18PaAMfVFZJoOeOc3TJQAbgkogdKAO9gE2ssKEDS0GEiYN6b
lpEVJ42wX39j1YXH7RWp3npoXfLDq4dwazLz63aShoyQSj3qiwVdck9ioWiEU5eKhRrOpVv76IH9
ms9IQbg7FMeu1ugy2Rq/qW2hdSd33S3lYwJY1WPvoc6liB2PgeaBEuSq6GC1NAuu57DI8cH8GGD5
ObLkiTSQBFM2HbJYHW08EJ3QNTfm5qLQV4w6LiurdQlZCtbNnrSxbdx78tSI402MwObBOSUUvO65
alVrdnwrZX4LFiRHKBCluiZJiyijfMBUfE4B2pReAhRqbbDTKzTWL3GXk9hPIUexQw0wVexKFsZ9
tWMk5d2GBuN6NOt8O9Qr7aOtj/NwUfoYy8pR3MG0NK6PuMYjvMRZPeeAOLMjZihbXz9tDxtjBrbm
AYjUb3BF56aMKRY0RDtmkY5fM2ArUSNr+f/5jLywo0JHkKp5/5BrnlyJ7tNBYi3x151uJznOmdlS
C3XmoM2w4d+dSrNZAr6T/fvakQEFwqSzcKVJPVQWBtgL1v5d49i743kdHJoNRpUGrMSgH2obAVw4
Ri4IiKgOQ90oArGM2aEAfBWwDKn5R5oHp/7UyQS8Y50qMb7YKsEATpSlO85mwHNSz3e8xT25VL4Z
M9cm9Y41vEVMvOVCBwGmx0j8w1Aw/c5HtPUasluQlWCuLLdpNvUYyReAF/loCGSXKvxdahN8MXl8
S0/EVHqhxpIpBiA9pVRhOZJzmjxSUT+DcnEGblN4rkbw32nKQropLiq74x5kh8kH0toIjQn+Qa3J
bxf4Vn9I7yEvn5NmMJQVR/aGbpTye0HrveFswzKnKcfHwm72ozzxuS6sL8QnOOa1JgzriF7wnT/N
n5OT+S2qjdRNhigLOEwBVu3S7gCt+ltWRUyUva2m3Z+SW/oA5R2SVEKJ/h6JGPl3+a1l+pmyFBE/
A9x+NCLMuBs+TUyKnrr1N7r9b7xdOzkvfprmLg5zKjsWXcGbH0Gh4wM3RL7zezSDrOuHL/nE9BVe
Vlbwq25MSUi8VViqOBcdXaP/0oTArGegki8ZNROzAACQfmS+snuZPOC/VIEw/40YeZbYbFWYzrNa
ZKNxqddBPX+FWkDTQVj1Jr9fI1nnrhLKe30y1+FYaKjLV2rfyBXV3YCDGIodH/MDSpftEBNmdAPN
IySaFQfcPDR8zcukxFLz1kxIcCoJG3wxFgsvVYdwQhP8sYJxNY02Ww6ZR9irjfr7H612viDbmRYU
4WtJq0ESqCSGyztv/7RKupkVeaYIklvXbkfBjC4m9JjnwrEb0SLvztqJ1WWIAlFQVEu/jK+vZ3NB
5nPsZhO1mWQcUIIhCvqqo7OEQZonVzuQ3POaOP3aKUysycAnu0oxtp8JBgablfVVYUuZZOvW+Yh4
JAR4chr9rv8fEzdYFcT0MH6SB8vP1nfP8Ee/qeLIhHpRNIfVDD1t7ECV30PqurYbzPN4nOsQ6jye
m+nSRc/bmIMeXMtQ7Jck2Fp67q2Si8BpK1IJBFNpsKP569n0QiibCvS0zsvR1GmenmkhZxEieP/A
HJMJbsHIkJ3U3kQFIYFUw37sgixhaQ7nHcFf6hkkTyZcMPrhXLCkRTz44pvUjwf6YDX+O70xKyPB
Tw1Maf0cwEF3TJijBM2aVYm0385b3CTzGefvXpvmRkv5kZ6+njkjCDegcaD7JXE/lBpBHmvyD2nJ
KW3H/oKQdKCJbL2Z65/VUxTxRkL1GY/tUqdbtjTIvMHgCOtRqT7VGTEtuk4Yw4k3rIQXtMQp3d62
vx7f9UFQ0mwWGWDF4QrafOWcSUDBI1QNW9SH35rYBK5tBG892S8Ppw55GknLVmevYPU7JBaSUrd0
uWY43pJD4SXZk6Zu5rB5YsJEv5qnrVtZXiBLDSqZueQZRjbWN/VEZJvZi7XTg1GUT9wh9D0/ZlQz
Vdcas25hvS/avUvm+Jwf/ZXYXlOcyxdvD4vlEfIfC+0xfmvvZBHfC9zrFoe0+j2btOukcM/OQpjn
xNGH3rUk2HhbnuvVqwiQG0Zh0O5kdwzd4ac8KupzceTPYCXg9jsJ0EcLs4JosCJ7dKgAxuRE7wF4
OM9SiXDQzpALfmbUocxruP7hio0Yh/2l69jk6Jqv9UTJnil3IQUwcS5BEX1WGx3HZI+wMUVLDQum
4yUj2GMOKL1sqFwBxo475/rktiNaeBFItNiXwdX2Tj8QRIyO0x60+3K7Vk2SsRtCHM2miUMbpc6Q
6tr+MJHUox/WNHQj6TMeAy2nb0+h1kB/gfmHV7cWjArwjwhg9FeOPy/N3f0cIlW2d968NGS0/HMV
+NH8KUF76W+rjN+cZSFovXeBewC0TRQLka+ZDm7p9JUri6UKXhgGmKN/Qh6g0MgOxJovx38v/A75
L8gPIMERGhAY/frsHECaERjBcInVBFYahAJT4pYutPfj3Nqv8rb88b2+C55b4dc9KYyITgGktr39
3osnm2vHBwHQFPEEAbAsvaS1v88ZdCF6BbvfOG2YSPDHwSh9iyyMSHXJ5e1rMAgtoHn1YPapbnsb
qwWObjprhw53CUALB62TbbwAYmN4BdD4qLhfnXZtSvN2BXZ1oXXLf7PR5dMqTn5egphdAGjCrJse
hFG9gxPxy0wb0InyKVvDPwgoSCYFaQ63rstomvgRizF31rYsM42vYtSWEHFnzOPgEdoCOOkMCNaR
WU2Jf8BS7MxjVshnR2q/LG1HvvYg6IwSCaiu4Mth/ZNUsAnoMp+RYqsjPEkjd5M7T/mAXh7yCQYR
r+kZuh/u2iRgmfXZvq987YoQuw3Cqfj9Ia8C+c0xQpLW62MzPH2Bv24QqQ4jAVrndwdxqbGT5IAq
o2dOEacoaXPd5wQYFa6cbPfStxBmbI+KCmBMnsNjnzCcmBl8aSt6xe1eNuISh+Z7A5hoPBUaBH9z
2oq4iJZgm/62O+QJLM6KafACOA/NBymDuUh2JTp0AA+4UTJThy+ArPfpLCrJowue/ovijPqokpuy
mfsarHkUZX5y56K3gmc0SykxkTB4levkE5p4TpEYm4bhDaql55K3YtLtTQkttTBFDl/rqcIkI/jX
lKvXoiTGRt7v7sN+qjZtG5zCuamcai6VHZd7DMgiK4CLYwP69MZDc0tz5QeWjxqIds/hKhmPq8wr
mwz3e0pGGftwJfSGd5RzB8YQMyUPivdk4CE/4ZrzDTpwq2WnsLUr7rwaIbobWKyd/jQopdAEoirH
Sa5/LJ2XjwHEae98EL+LTrATaV6VUrTwtmxLvOlYsWUoEOWqeNbmuAqMFFDkJJKslHDMcPApru6b
ussVTKPSTV5Zrob2zZ1urPgsTfOFUEm0Yj6l1yVsbFZi0t1Xwf2aDRdd4bo53BYBW7qyXQ0EVkuB
/5pwRkC/iHsKqXpwMBM/oS3nq1J4Rt94TccqZ3C+XtfB2lcvO2jIGUQZdC49qlk1Zmp3gkuR8Zrb
AzI66U+KoN23xc9QAT+mcjoR8EkdCzjkx+koM0MB5/+D0KmYOqBdWFxaN21x4CACxbiM87isFsvr
icw88jWJdfBVMq7DFs9Biom2nzkNOFFQqW1lkLVLroM/gC82Y/gf7aHiSy/Dx0+I4JdGvntCPWbv
Pdxc3SJzwchQZaj5AUh0wdAw/cnPkexj5cCCls1mOd7UggyMzSAohlwL65LYXDUIJTX/LNocaXHS
t9bqtSt1xOLOxRSZohyr8fX2Gj5exu0MrkyoGsIFhznIJRifx3r7PCNCzHJBIsVYFjiOGoUbgA4X
31xKSUG8ZQpzBS/4bCvKrdsb9lIu/3NTrY05dC+scimZaRNPInir8LOK0yJmqgjuQr5AuUhVaTBN
NgnUoy0A8uXv4Ynd92m6XkTlThEibGDE+PrumcIisXWWADBf4mLQ+c5GjP++vlxmnu4hzRMw4qY4
L6jIrsc+zAzwjgdkO9eUwoIBxNfk2McW5nAs1z/zIKH/quKLYEwZy276QzyHByTChpZkCOvF6DBK
mgHKptCHAAt97ZnCglxjsMpniWmBGurFaStPbC7zc0h/c7mktAt6IOl+dnugZGMjpcF/BXZCrItJ
XQWru4iJumV1H9gRlayWMamRthK6HwJtZJYbr8JJ41PQX10xp1F6t1BFDlXDzSWk6bFTahv9F7EM
UjWauD7jffut5cd6YC/vNUfXHa2FJUGmt5VA5vqEi5Y1IR2QCgWTBWKxaHsLRh3VxQxaDnVT+o+I
UvBacEG/FBoolWjJewPGjlLLz2Rgg3bT1uj0Nt3HY5y0g7WqMt4YOKBlNqD77LRiRaivKYkdfVXq
VecW84GvpFECgTHvckUY072zv4cIesuTHwClEAaT2hfhn9MzCapj0KismpagaNm9BJ9GRXfttvsM
me1naCQcbbXw3boM51hzKpZV0cw81DdGFD3ihDuMvfYCrGE8szFyYi0/sgCVgNlfW5S7vC8aYkh+
75DGZVGkz1/stOuCohlBDmoMj6GqGZOmGkL0cPze9It5BXVYvUkRIE1Q4jqybmufA9tPeHKJxEKc
kkwg3VnCzwxqTaqW5cUwM8LG0W617gUpDE+32aeKgJyfAH9esY7WTjFeV0moCKwYqlLkX+CKo6NU
1/yeLP6UNc1vuTa6uX4d8N/VMvYDZ2vJZ8osrlN80JEXiq/OMQzw5sjF0Wd/Pqr4rFmnvOc1bSY4
Nl2t2vZuBxqKrRCJ6xL4CY33+dVtPIOZ5pBd5ygoEhyFdPAjUJ7VkZPJm9nh6b5djA7C5B9N7KeW
jtRbkbqwC8fXtjpo5eqWpdqcGY7fdy3IQvoTa5MtfmZVZQqgkLyfRPUNS77j/4bnYJDNArTL2TuQ
mSu9hOkloZ2HwsxgsHDVZDfEQp1bsk8wfPqsqkpR4geXIvAZKn48IxIuG4YtY6ZyesfFxe75QpEw
lr5Qp8cYp/rTTsxqMguN0vqe1TLPFY2jphIZhoofmClcKc3trstclTsWBXspKC6e6Bl7hOr6fGgW
t3kd4nDUspBvWkQxtABhKMhMgHuePhAtaTcdmgv+B+Mh9xWYOLCi6RmI7I4jrrm7GD6KV8qwedWv
d+GcNIPYMQhzXEQ3ygiDZYPObu5BLhe7l4SfXOjAETAtkOzbUgCIjCKW8u8yNLl31w3XGT3nqRvh
QldZ6ybPBAMe3mKZ7RD4nkGD15hG30bW4sH1EiTgd1bNAJ9oqI/dqB4zQlbREvGCZDIPjkpIsoLN
Ig8xDu2xP7qy7efIisK9mtQPfpqxNxzMeK+ZfGjOitMzB/f6VfxonJKc0LvL3Iq9GJ5MVf+1B18w
ENJBSdpDAAv5D9U8juIcWlCvjLYbNTpYlpr5OxxIsbzpWuf8CJsgY4w5QfuK3vAIImvYlA1SYffb
XiPVBsg76AqMWXLT6yw0HXzswVE1v0s4udRyycIsmBy0LeDbcHmX0eWfvzQlKMq8vP/2l34o5crV
5LwFoH9h1ybh5Td/AQGECq+IwRlQOEfcR16SLHFw2SUj0KHyQwB0LCVxNDmY8LrMM96idLepvCOu
tbJRXHWn17+QnqHY/xm5qZAyKTWuZv9ZEClB4a7m7FUGaxzabSWBMLA8bceaiSlIAJHbbNqLO9wP
/R4+jgLiN8GCr/v7pG4n7WO1N/kOFLSZo23/RL8TxdTZ9bHZp5S3kO7k/+SsVXTj5mZle/NQDolH
Fuo2zyGen4Rxn+giVypL1yZnVsTbfE1q6AEZjZRAppkE44+Rna3yLTrV6cB3c80vwQELLr1eRGM0
A/70jgtNaC+YZEN7WVx981P/X6EdMHz6j+vaVK4sJx2qq9pl0t7zziB2ISDhCibknzspfj8d0vG+
8//UGjgC4v3ro1glWlW9fP2qcgx1YDgct2G15naX7/x4LJox9u43BEwAV20vmOojV8xkhwCbTsbA
f4S1dg80YX8PVy9wqH55R03q1a0SCpht5eUlYMuHULyNmeX6tPeLHOMkVrjEniBFT+/qq/WpjfQW
n+J2VW+Vyvduyo9T4xwhfAc+/w3kNIg+AiyZOAMiu2PSLCgfu+PCb4yHuEJyqHR9CNcKyYsf0D71
xuxK2Z3fqah07D6ZKwoc7LPfMgOpwCL5TbLgbzFDcZfAsMcw+LDYEwJ0E+R2VXpNgBYMc0H6p/6B
eFWkg4VRY5cSDor7K08AYjCltPKnuwYIPsXhK0QPdXDJCVHuwDh3XSqR2hVBaWAOBeWKezPpvumI
Uaev1jSdzn12mBWshec/t8LnQqxSHtejcTqMDSvyBhlIk0iMZafEoiiKAp5bZxRUZCDqFMdJuvCZ
SeKCfVyDK+tI4yE+399x/k3i02DqV35F73bqZNRW9hpNlH4wK7N70atYiatH5OkdY0w5OyTZzEUW
KA2gDSGBAS0dV5nsdXFXWNwAClyelJENziA6JemzYX252b2TEuMEWxrKQhmu2W7z1n5P4TBEvmHr
pgXWN1u/t7RdeF0j+79P3Av8Un5n7oSh0tjComAN1jDOLSpfBlkYR+9fM1RFL0vkfJfTNBiQ/zN+
DX+6RO86YXxKJGDDQM0s39C16IJPo3OXAnOdtXMuA1PhaGahuURbQHlS3sZdQrriDYjZIQ12kDQk
AZGaev1QviW/qGPtvrfGFDsMHbjsnVZCXrzqphPvl4eI6FCIJuUVdWCNKGj6P+D9bYNdcxcuvmX+
44J6KciDm0hmsvrD/ynCb7kl9kJzoY2VfDgZfffJHuSYPnS2S2b/3dXDoAnd28LJ+7uhC2KFjVFd
8czfIFW0Eu+BUMcqdbFmA4cEmpBLrKEizDx+PrEaTVGOaLZOLVjz/47dGtOatKxineLbk0l7tCxh
UX0FIZ8s8aFcxS5gWeF1wy06tGeePLMRcxTzesXU76GVns9XuRr6gVzQCYCYppACZuSpuQAGlhFN
DdtXwYLagCcDPpRDCPzj1qs6DBkrAob4urR/kP7rBrua//BxdMUslvro+8xTlItEeh2/AHZkkjrQ
1x0ytX298lM9HFKc0qQG4Okv1S91Is/P0AbFDILeq/mzxbXdzear5fHKQWjoUILB8gJ7djd6TX4p
aQf7FVbNYHemFJDhtJ+t78U2c7RGjvBw63CLKIksW9uknKJty42tJqFo4f1alNlLfKBgY6JBCuY3
raIAF9GU++CzIKDbCakg0JlC4wWWcuS3OOVdfmb62jlbSi90f7QMZdVvta7kxICCyp2L0nL9pUhR
VX1uYEKn0vlog7dk9aPMu3WxhluojaxEImAN/ajZtjaF3zjyaRE+TsVQtyRJAveLsE1H3xj4lYqv
TKii8GkuiNr2CmBDuC5/EvHThv0WJLGYUXZ08hGNJcgyBPJS/+j/4m7QTr4CnXcomKOKwGxIzfGL
CNJPiVY8xo6b5k+0gtEQbPVawYr8emGCLNN/esHqxdzINUYVLdA9S3GkXGhd5KRAtxfAXiE9RqXu
qjfbnTbF15ODZntRE0ibQpvyC6Rs/uR2pUCS9tRQhRE2GvksZ56jO65euorfq9mXJWLu9KQM/5ow
1lsQivDSgm9/aKV9r0BF9eTO2o+GogzKQ/6IzU38XzSfJZJuQiWZ8k/y9byqDYtrlpXPrqSQHKQM
w/UisDjiw6KO7BUKszpZX5J8RblztrDOowVm9WftxaswtnbXi7fEA+CSo0wEtPnpLSaK09l+sol3
8jbDs18N+0bjf7SNHyl5aWPJppvWdESTrRLqUP0YH9AtskR/PX4it9a7/KE2OUqBwsnb99KZ0v6q
LlLNxpKIXk+BqdXLvlsECR7kgeoVM24hYhWghqazovzkPDsPRJvuEGQTcMD4X56F9ud1loMShrmC
KPsktiC8jHPLbH6q9XX5AF0Bzdg8wPVy+Gkpei1JemelCTZopMbml08HJXNTQsgDTYXykkrEcD4R
ehQkK4vhq/jRhG07pAtfUVEmcxzNd5ziOTXX7Emd+Ihdmh3qn+TU1ONySNflUCYMzhsA7KajDlAI
xdkbbeSwpVs3jrrlkLN1/FCTn+hUylZZfw6/9DdsRrR9kH//8coJ2gBIX5iriys/BbrT3wofDUok
bgEzA5XJvdkCRz4Y3sCDA27MzUomgPM4TvttJHC0gvHdQwVFN61j67qhDbE+m98uT3tsPMDCydgM
h9kbduc4Pr+bmxXmaHanWA5x0s2NyHmEOQJINbVWuNiV7gTYoujKnXaa3fxiBUckYUs9G8MtU+bV
1n1vIJafEanxYHVkIC0q7A3cEszhM9iYYCddyMFyRrmvLOl/+TT88itR6iHMGLxNNJloL/RBKqWi
J9z+Waz5ix+fkU0Qq47pzUBlmIZy3kaDvnP+1bTT7+cRgBgnZ3HGj0hYQ0X8JhUao99HtiG6ukD+
gVorFre0mjpDFNb3WCcHAlls5ovSFZawSZrwgUPCqraqRGLpOOve5Aw218a7sutQwaqNVLikUV97
PS++qTvIK6TIQ5c0IcfQDCLAxO/zYAYyOFeG1eVHI7OgC9e8w/JnzjsE2YxkXj/5tF6kyh9S/MYq
gvwwaBkWpmuH4NLbRyPj7gynnbsUjW92/RE4mPAghkiN+xcnPsOAnzIhpIMrvoKpjdyNpbJrxfXn
psyE7kl/NpTkxSD+e4KHBeWwUtrZnHS+xK/LkI7ixJz9mkAcve0KTO78E/xRIrJnux5O1pHjh3UX
/mb69IdFp1UzQtIQfMNTuPZ/4MvobuuU8FU/4R5ZlDpXeiHG0Y8bPSKPY+EIeaJVnK0qhYU8nkBp
tFLW8kUgpTMTa42qB9NRAWURNcaD3xdkJuPMuhzNEc4DCD4Z4wbLG2dfMPHz+wuQUDq1xAN4t5Tq
T9zHACC9PtTqlpz8aczm69JkXNo0EwsbcqbGH9F5+MqNvZ/QEDfzX6rhcPu9pLOuHkomT8+pOxE7
MoctieT0yHWkQmsPoWoeu03QyVx9CKfzrqs1HTyHKfWynBEAQ1IboThEEdYrUtB1IB/7MlewT9Ae
8ZKSfECQnE5aFrbgYMcvwOU7g2pFYuo2yIE4cjOTn/qlkE2mHfhgXPGasCSxE2X9kyXX1IylTp5Q
Ve1UR6tHzyX6uepWhxAvaj2v3wK4RKHQlShw/SACKzVOT7WblwZSCM76/dUdf+SsTLfzdqS5bi29
nuIlas4b7FH6ec5oYnPPD9Xv+eXq+Jxro20+EMyv2oJV7SSF/fdrIBqxn1mCfqRTLPAvDBecLDEU
prg5WSW/rgXHvuzjJOhsEhokPpKUVyptmv9HI5GwIuOP23k4q9SEVmFpbRCSwhP6Vl64mNVQALX4
sC1UlqLCCzOTRd5SSUALmduaDj6gyvyGYzjx/BmDs1ANfhvOwui8idDF4ZX2gLXvutEPW/jctJ6F
dOwzcFbrA9h3iQb54wJ7ui0qaGmEnB9nZCEpXeLbm0TCZUf1hPvgT6Mfq0Y9TgKTdh81I/OTqXXJ
Q+agk2P3XhRpmjKhFbEcJ2pgJw5ZYhhn9ToXq5mLBOzjoUE8Tp6u4pblw7dHFVT4xquJjrwZj6dI
RgYWXzYjD48PSZAbKGQR/fDvCOcQQnA+I4WjDdYbpPckylA5Mboy/U3j6PIr+gRy3iiMtu9VYgqi
ZZNCTcwt6Pjp+musrxzJHTvTo07KMoJoadoalhfR7tKm1YycYnsvp+HBSAV+K8mB9hnRPCr/VtNT
K11/aoTWXTRz5ujZujrZmXH77F5Jp8UFt67vpCGDerkcZSK+IdmX1iZ3AFMnHdZRSjzsLHPJC6UE
/aLHYnWyoQG8JeXazTItY+aVn/6cV0AD1/ZYW5SuGPkdarKq4ROOkeHegL9U2zayLo/oRufXpiua
Fl/Jzyjpehel2UGAod4V5jd6Jnzddi9dKv0azCKGO3POavECZhxsRfisQ5Sw2H+DmM+Mrr3Ekge3
shx06RbRJ4v1uQx0idYljZ41qysgxqJ8HWJebdtl9Xh732flMoas5Sw8zqvlEZ7WDd8FgmfbcW85
v5xdjo2sRvhK2OjtPutb0RNuHmOwVvbvhiWvuhzwPcqTKGRTpeOI7pGGmd9rmJyWdI55jjwU9txW
UO5kv31qGxniaLBm+Dytf6QWmEHl1jKlTzjq/v4r229g+KLyDHvzvgXMzlpGbaWq9fHbRUleBVhB
TbhnEbcAwygbOmQVi1uBIicSyqv3eIKvWg3266qRmu9yArpausOkTVE4oogsqHwtYtaCicMsW5k0
/uGYaBq3gvbz2Rv6ZaV/L25yH5c4dn2Y//owC8C2h4zLTQ5rC3I3msYAV/AFRmWhBJh4iiuXtWAG
6WSSQIUsR2CaBczC9cMHXoznu251IKzHgHs6r97S5tJO7O1R8HS0kEXj/83o5dxG1/wADl2W8Esz
ZtCLdAmjjos1pp98+KPVU2Rf1g6zDxgdE8HEjKYXNo+1EZ9S5mdHfzcP/hv4xOcAq9kghu5FbxeX
QrqgmWqMUY427Lh//LhRVCTzxgzKE10MDjMBliKaB92g8+hPcfC0RNMN/hFqNLbWLi1pL25dLnV7
VaetdkafYY4ofMrd8FPBiiql1r3jGOwuiSoA1SP11r8CuKfrP40ojgJWKWz7rhw5syIo/FFxtfNs
Z77QJLaGqAlCHtLbsT9pFJUMc511BPrdjvpEyQ/V8KNF9QWDYBxf+Ue0Xrq5A3oeul+6jZkSp8a0
QEikYMh6RpBRckwgEBUYn/B7ND2xewwMTk+AP1WXwgV+jyG0v6MXnlWlPlJwvd73s001exsd5pCU
UyxK5RoFG2+Qb1viet8v2+fppHskp+6zo+JAUon/L1x0nkP6i46PjWZmAhkOB3Gcz9qveucQ8daZ
hF1SStUl1orRaio2a1hqyyiXFIFD/rMpBNsv8tu4/Bfs3T1F1LVA4I9Bw2L37/EHvMOhOahUUGxH
5E6MnaS3Y+jqPKOn3Uo0mdKD9G61P1pMxxfzFyz802CXBur86M5OeG8gQSLqt5hyjO0ULbjuBIU8
taXhpbWovm/wYYj+MF7gCcA3Ci2XR6K3tN+TGDDoHYY2M8oIxdPN1xUjYlc3Sqgka5bSZ8mQofcb
NvY8D93R0tTX60zMFGC2iqtrKzaP0D7UtdFR6O69SIQNpXlq9LzmBI977Tl1IDBbr6DYv0Jv53/t
8F6Sq3gw6JiuOrsk4TVolTu4jzoIs7fbjlBGnwVe8sNlzD13k+xzZiu4QPYBj0U7JDfTQscEkZZ2
IIeSupdhzh3lzRoIMElNSuI5Pp6NKakv5WqjBe/oO92J43OvgMNySUc6lYLTkP6qSn0mvcAbjyW0
X6MSaaEXxenaxh4HYSx269cQhJloi+qMjtO53xNs6OVMcGA2Ix7V576cT7XxLjorL4LcgO+XjQE4
ljvzI4mWVz0B6VUWPQm3Z/Wp5XIsb8tMoZvNDAx2/BzQH+C+aA9VhsFla2qtDz0soUdeWBu6xCrW
pBhbNHw4nccyqO3UjKmU1jrUzmV33KK7uXwX4YPLPvSp99AyYEijlrL9con2ukv3Qndo0q2fT4ST
70b1SCXXTKuPvPHgIk4j7aAnZ4wdeXHqaIftjWDg+LbzaLY3BUCBjlQ0HAh3d2OOvZ9OtrHM2Hwl
1DozmgasI1mR89JeuJGvDh8zir17hm+fNy6Q7q+3XbMFDLPmkhABoaqPiVUrHpvbrYGyBRO6z1e0
URHkBoyc8/p1huza5SBLFBphiYxtHphhifuA2B7+ra/aXH0Ppsb1fjupsRXYNbnpXeUWz0JN3RjP
v+hoLLOTfB2lLk9JicxxsEHYoM/3MCDSwOUL0RaEpGqrMyvgstALU+EnkKuFZmZ98dJfFmt8iOBu
xSFgmj2RHbi7vsJGaQ5o3DMmZmbeyH6PYuEPxTQEe3rX5n0g7SMMP77eNPwqeW30q0s5ZWl6bzji
3jFjfgNFGld311rQUHkowxcFoItaWkGKcIVcAGkYePXMNLAvUXFff1PKAjr0hkaRN6I5B/qv7aYz
AK/Z2H7UmMciAmkyiGJ6jHv/6FJoZ9AJh/9lqPpvYmc/LOiCj41pm6+Lp7myIf+kLVoG7GX4xnLw
Jh0cffoBrh+OWpyO3+oDBPzx7HKVnyl2Lv8QlxvhZnqqhkjhAUcHkZswS+nmr3QN/GkcTFwafohM
SRc09rmlGf8d3FBufDRawJlMJq8gwa5m0M32K+XOGdNkgvcOa+ndjsD9h0OYFzzp+g/eG0Zlgq+N
LKeiWPmEtncKdk8LPZXGhFJmivG/1iYTG2el7DiQgUsTUOoaPXsF+ibpYVuucduEqipvM69+BWPa
xk+TxU2yKZCC56z8jE8DbG94G2lTlYlheYvsQbJgsiPGLY4MJSDq8ddyhkgSLR4ZQgQYXPw09I1F
boHtBZTwY2hLGxryiV289NiEbrMNBbkNWPXGgkx680ZjM9HQVuMtBhBpbWZR8wJY3Tq8wi4bgY5w
4/2a4NmPXsh/rBj2wQcjLEvoB+OQqgTPiSU6iBZs5+xpZ22ybkoCXlKYrVXB0pa/TW44Qh+ChbiS
NkgJwhoPC/ck26r/W8X3bl6eu0AIYqBz1oWcBL+3sOjgHjh5CYEIo/yn8p1gt6pwreuqyaVBtncL
kWcujxBI69WCWf1176LNILqm2nI+Ok84kJ3OAgoG0W+06ntx+FPAs4aGIHgC1NfAUV3TyGJsulz/
KPBKzRD88xE3LRxP5guzB8pFRA1ukrrzob91CelfyyTvYL3yMJbEQ6sif4/KzFXuYelacZa/pKsD
rbOUCiG+9D6UZsDK9J5RtFTMVRymIV3U+706Xj/oXaeW0/ZZLdAFZEf9zPWcn3uBw181c2hlVcLm
/blSYXB9wWjWz0HfPVEiSH7Gu993BS9EzyV3xVyfwXONUDNRdBDchk6wm49NqzmbYK7xRmQSmrOG
fantxvd+OKTmF6TXRCdekbJfLIpOA1Mk7BmQ8FdsVuoJpzizX1wEWrP99ciXSvOHxbaJXHmQ7iJk
7NR4m8TuoSzrjqusdAwi+YRumCXxREnk3bV1ccKzW8Kwr8OBR3diR8ivxO8RIL6AF3a3d/i547Ix
dddqvRmjU4QxcNyhNoeDK9vnZylPuFkKOdZrLIFAwJ1uWaHVp6/+Oa9s8/so1kRL0GiHC37HogTJ
/n6bxYI97HqHX4fLmWLyGJ7gn9aoUXHbR6TnY7EJ0VlKN1vE3znvEtKyjAt+MqyyYQ3usqKmqFDr
AjsJcOKmMnJL0VOQqw4YmMe2DGu4s2ie2CnbenQL1lIXzY7cPKlygC+WVr6U2sqGFRy0NRdcOFb6
p7qH2snhaoZB1fTIOT8P1UAQ9pjQ/+f2BGdE2De+/4iqDbe05nxi/AQDd1j+74EwX/+UdEOgpVfG
9w0hWQ/Q90vp2GLfZLUhgRKJMng4jMTgPiLLcNm5sgHePmIMeFlftNA0HVOoHI9HiGTn1kiNzB37
yZuYsm1uEcBmskNQ5y+JsB0IOR0QyhY92hAAV8vx2EApEEpKAT0gcUXjDOhJ65+I7p3VtBC4OzOZ
AEAwcj14f7kdhDKHfGa8BCkhs7CD5sManJOuHRL25H362ZTHTKqLIio916NlxYtxibg2kf7Pp75c
Y4CbVZj3L41AROSLH1kOIKFsG9UOEt+/rE3DijqxU80l+7FL/kr5pD2T00Vhlxmilu9W7aKxidFy
x5yZ98ZLtMNanmg9RmLQqOqJ90Yi4ThbeRFYzdPQb++4gbuTN/t6qKiBFXSddxMPjpnRjB1CZcZ3
8UwluzfaRZmSsVpa/+DTZc4XT3n3cQTT8Pup1CoiwX+gO49XLyrQJVn69xEOUuUyGkpB6qs49L7w
TfgD5k0gCQoYyVObmDl6yYBvMsF4qSK8F/1ivrmh3DXOLvhhOY4Xbc1/NxjldIz+OghFbW1Cag5M
inuqPBCpUhYeOl1oS/e8mVMeezNKgWNj9D4za575IYNtZUAw1XyL49Ysg1ts4xOX/lDBflA+IZ3G
Wn+gTdZE4978+5Twr0oSDiSbWnN7iRVzXDgtKeZcGZV9F1AWdFemYGaNeEyB2GPhLcI+cMUFs5XY
5BRNXxtyHTB1ddbNT3m20OcUIJMrnESj+stPTgt/I4tFHDIrX73bL4KB5jhVuGKK62wybLYBH6H8
nA1Jdh1FjpF3j4qJ6q+npijsOh45SOI6PR+enm3I5dyjivJ/z0QoFQtwEgvkQxj7PMLN+nmSoVh2
W/Tq+USm8Dwgfgm0tKNVmuy40XxDxSs48xIxbBHMV0dC6OXii4l2i/KQPdLDitEwKHeQ5V8pLhIr
N9L2zK3RHJvmpdCrE+lSF+Du/aOzWgUFuoHMPQVRFiV0GnxkMPt2wdRpKeUgZNseg32KnYpatf2Q
MO6fA5icblPuvTvLpva+LBvVlmj9IvAbfj7OyHaxikL4dj0r+sepgclWvPzUVSBW8EQwOPiRfg4w
faEQ1FD7M1IktqHo5tod82xIOpfxlz213h1ixdeyVkrdPZ0P5cnoiX5MtkkiSD4Ju1wfKuV4IwK3
L8RalXncrhpS4FwtBWZfphTYq5GFHvunR3di16q29Dvp0TcxtDJlIVFBfc9b2ITmL8Pc6SnwXbGm
ahK9f01vGawMlgDWKc9cvnBqQqCC2TPQG6iPCM1XXsxA6vjCJ9FthqSZYDaokZxOMCXhJOoU50iM
ZA7p6dT5x9uIO6LGUPPYLOjuw4BVUsaZCzJa3Z147nncw4h7f+Yp3z1bs1+zod1SCpt0cux2zFrL
woY01hGVRPuEWgXyLgkWW9ut7FVfzgGweq5S3aEMp4ggPovDZAWuDU/HqFlE5hSvIFGkWDtuuKoF
51AvwFo+Q6zVRuB9AiCDRVe9UDtPxkPcGu+T1zTjZVXvQhCszg1ZSWrAWmmXrEcYcslVbLn7S3go
BT0B9D3HkChJn+tdB4QL78BxDSw12Hu6C4PNU56MIp5ddrrca/caePmG2HMHVlbD4YlUG3UTV8i/
eZlG6Iqu/S4p1uIGDHcPQC4LWCoeYw3qoHWVD/Ma39Nv4ckSth9MGuoULNDXTmfIAXr7BWNfByjG
eM3rhjdI0XqTOxKVxYLhqBO/w981YDyDzKMuMNtakSS1Ct9aTaufAXnhbRtGHKyDkS9pnasEuvTf
mGtHvBYcgGZVYe9y1BVEX4HwX5HffFDJecrQm2yo8lY9y09DAxIS50bItf4AKyYR6HpqQfiHEqEK
U53hVssA7GuBFf0nj79lYvu8vsTTJvFyhb/8S9KbdiBAcSE/4opVAOO5t8ysa6hQ37hKlCR5ARb+
gNbD8N1pr7IkVHkZT8SMejBNBKmGwoJDEImxQFGjRZD4rlJ7wFExQ2vZOOe/q90lNlzILZ6icTex
PpzsznfgKmdAvbnDxaRKT5if8X0O3nPUJFVNDfs8tZH0COAQmOm8xjTd9mY/xzWyp3DwMKeCpaBO
UXAJnJX/hw+PW8JI/2QcOhtXoORgqbeRRRdqZTCg8P5TaggbXR+i0kos7cqV6QziLGWV17r4o8gj
FMmL8b7xn0uHdPGVjVowF+Rb/QsNDkmtvTA+BCYMV5hxh8U7oybBFSo/m+EitSiz0NOoaX5Xb6+f
EaI0asJVhHzuAuz96gp/ZC4f2uH5RrDmo0Fcwv9AOlx89b60lxoqblkNk6+WR6jwEx6zKfk1b2ul
lK2AWdnYd0eczc24b/Z9QTM8KkTuDrjmW15GwSiROK+TrzHt8wf+jV4CCmF5a5g4KCm5NLuNp+0d
1Ggs9acA0Hmzp51d5qGjgc1Hd8+MNfbq0nkeV/EELRsiBImiW4DW8zcTNzUhHy78Sj6JXCWgHyj5
QATFHJl4le8x29jN08wxH71S5sH53yt3w+vVohgtvYxU1gsH1Dqq5Z0L9AKjjH0kBGLHO2SSq2zl
57Qg+E/ORL+4UCr4/tyNE/m9L5RWCpbj4X3i6WBRXkJsc5LZvQeHHfkLkZQiuGXg/Xv6Xb4GV875
2KbYNW/pEOX9b+oGuV6vw2CKHssOjf/wtVmFSa/YuqjNGhmJwP9z43eNT2yvzddgZuaGYq5slmlH
iOTtoSWc1915GA5XbqLBBTpQVtBTfT29hymytB/SM8xrF2rwNUX1wUUdIuNMjEszhbpRXH9AmpSl
GNjppU/Y3O39R3O460VCXwvQmv7Y0mae35VxAGcKKzNcO6MOg6op2qCYX924mOkzFRUXW9wT5ZZD
ukemfEaN7p5XUUigJQ+Ev4dmUK2rMJl4lYfO9gPjcO5clvn4867je+4sbjzXkaIDUY2k5wbDd+hC
ssISPuvPnq4PY6iJzSQWFbD8HjgWnHreFPnkNBrC1MZ2X/HQWD8f1JQxLoDq2mvhp9zeP5usjA1m
aQblSQ6pOsz1psHIMgHBHQlE6Na6vvtrmc4JV2t1yTV92dTYBYIqeZF4uOEGHrOtLBcxCKRv9NNc
sBkRUVgm1xpBiEIiGluTurBVuYIMxyoy/syC+f91WBvFHZa0Wrhb7/QQXxtI4S4kOFsELny+v8J2
cisMeUpqGFiwx3BIrgYga87Pve8b/xHPBkHJCPABOB7CN/9pye3j/hs5AGGbcqTAXkLFkHt56n0b
OG7pc7EhoAtrC67fKe9seJe3O1ntDQyAlrIq1XlzpbyYgQwOnVjASDfdVPARWVI1iEjHo0bQaKSu
GmCOq1933b3RgcX8ZJe1hnMA7qG802Fy94xKWzb3NzpQZ5cGwNxmKV7fUyzKYa2SB25f1mP8CuWo
/XnJK2y2YxBNk+o1gOYijKyMBsHseI8EzR1HGjL/uSU+K+uFTmi+m5drLExaFliAhYErnUXR/MrP
0O0kL2vwMz4vu3TGoA+b4TQ84fB70fyi6Pa2ru7T27l4KTqryQjomEKgksU8AqfyhCBt/1Y4uNuj
pUhud1XIWEueHkzalJ1VgsAoqrAFdORd2p845RG01VNzm15GPSds2PhaYwe1h3nExV8rj8t0qt0o
BqFfXSym9l9NE231x2ErxpXIPW23NCPeBL3V0w1lbL8YqahkcUEnl4NZDzLZyMhzEqRuA234Fz7i
SYNyf6JJqdZXmTM9Jqp3aKtuZQtG52MF8RiTRveRzs8cBUVqW+oucrcmplqISEcnsgN+tlGzspKh
pJuIdGRPDIoctrwTahUeu4h184n2Apr1zgaM4fViAe4w+jrz4MTnhsRh5129qFnfL+ZUxr+bMGQL
8/I8vemw+OQftFCjCePLm05OKhoIMFT6Mks07eXEzvPf/Q6ELvF0croxpba+at4wIfgUx3k9QJtS
2hs0zrKv0Vh0sSA8vfJKLYgKk97RvBXQzS9pF9LdV8lxvpzcN3t10NH7mT+XIcZk7NL5a5rIFDC0
Rg4kOscAOylbK/HjkpDoCXrMRzuhtjDeTFiDZ8NTrfvKKZzghS5n9dFtHFBMDndE1oc0tDIrOZX4
rkonYPnU1R30LMwRk8XDHUgvOZh04H9PgSgMCfXVFBLhfHeo9lXwz3ruoUqbSRl+JSYXT1p3rjbQ
GCe4La15H1OnJt4xOEHkRFvtWQTMCC6flWDrI9KqkyGNfLqin70o4EZQ9ZpYbSb5t5bj8RJbxgAO
l9ADUGmWTk5B20FA958InhZSrPJS2v6chPyEvmcDLnEp1ikk6lW4fUgXY/oGT0dhwe9IhOtCDWC/
2yPFJg5tRe++oE0PB0sYg0OmqnJnaEZ10DbJ548kHxbaoaO4ap42CE6tXJi4x4ezRW2l/DDltn4y
yG85C51VlZbVpyW5SWtH82qrzE0hcrmilOsfW0pdCd6c/srnwjri/gNufCZVXDDPPDmEKBymIpgX
subdhJrJ7Xeq0zsBhpK9wlhebK5TqBoXRRI1Tgd7qoi+SblVk74xG1cOHTlFq8HZv8FNzWQud0qw
LW5z13arhxJEF1PBFXf6vy9y3MtE5Md1dNNPn3Bg3NJHjxP5X2jQSTq9k3vbMWxjb2rgfszsOgid
th7zTEq/XtSvBILpV0umjV0EjrIjiujC/lOG+GlDtfcCbShPsvGmxGX0yWxqgBqBbeH2YfcPmj0p
LpRlNiwXUfnzppDBkHNf2ZuCs8/1T2vX7HWVD+kx9dj32ug0B2n4qLqsaTXYTYiS+LQHvMk4t+S1
eLob8hcQpDeHfN5vb4mH1BeNA/1+XHn2IKzwEmK/NWKn0KvDP62Zmci6Ocl0WMXNOMypw8eh+exy
mnWRLbG36hnxjUtECLjArtPcWIMDlnDkjF73a0FLAevpMgIFiEPGTryA2dNn+CRBsJ+n4cQKL0oF
41Bk5G+SXdvjCqjuzDJfI2JQGhyiwbq3MFMt6OBf/ITIqhTf7PFblwgRqDqqhiOl/Wtni8z/mrCt
1bGL0s4ZE6iSULzmTj1mm1cWzbKJY+boCYgDC9PPR8qgT4MaJGc9CgFW+MkPdT22jayPk6AbOFkV
OAJL61nCnHa34uvtm3KQDAXuU6xwtjS33Ml4PKGiJZGDCZtfVu5ru9VrfLuuAzCECyT94uU/S+XM
HV2BZ6ZzpkUJSRIaVad5Gurls3JyWnNDSF2NBdWxOZtYSlMAa/aVIBPneu+3UE3u1zKtWKOi3oqc
E6rRX8tT7CqjC9OjqPtf4U00oJiCvu3PL5WlQBo4+2/WQfReojMxeg+ogTETNvte38rjp6pgBNr8
o3KmHfDeUV7ZgyQPi0OgZ/NkryOJUhCuKUJOMobrMOdFuPELif1xUtRB7YTsJ6UbhkkrcG/OFITE
8Lrs84jzbzzYjDanBoF/Q7MytKny/qeGi0RTxTNrbeRquM0ERMGRNMmNIMTMN1VYNHSeiHjhru2K
mzNA9AtcU8ByEheerKBz497U8mstXXxZbgl5FikU5fvPrWKG3GHKQaQiGUZtDSyi7ivqv2b+c/ll
wGVa850g56FNQJCsY9xPejg9qHHliQ/G+cUJx20POcVDjeJ5jDqQQ0d8ejDeoUcf3OKXzOSIfy33
8KtdhuD41nzlfsysP7tclKb0tBUbCK7VjMnZtWRYz0iWPqO1fe3JJeH98uKRYpF5uZNuYk2VMHWN
OhWU67VHI6c/kIK3ukGjEro8bNxRtGRSjuPtKhSyoq+KK5YJHblXp+7QziN7DUti78lNioKJI6ZV
k2aYBx3rOja2V+J16w3PZh3wGtyRZY2Au2mc3vfcGKEGsAWQWK1l9jKro1RZcnaG6/wbN2lXCwaH
dbtTDn3SEyfqPgNG5m9cDqH5lL0NBRCcjj142huelnBi1Ymrab1vqjqdD2pKIiWE/ZTcgN2jzAKe
cyo3WXPpOwceRe04SPRltRAyr7HvcFo0Axl5upR4LfDNV/GzVbqqKS0uh+j57S9RgyZ0b7/Gm3pH
LdVbSA0LjHvmdCYJUvdle0Jjtk+HD++Asx8HvaDJuPcVy6QesY5lyQQulBZzjgDI7EsHDdB2FvpD
NDfzglGRug8btZmnvr1hdomw656AHuSDjr4pZSsV+UMyLsziscrOdyRZ+2bqXoCmNXzVNkXnSRNT
L1K+vSAMYvZo1/aRUJkeJB0/Eht6yUS72yMCTyYXEBtqyft89YFwnNt1mXqIvq0wRJ1fwEmqHqiL
5lnkpJ4nWI63uQuqhOjCvafxogpsDlZANFjx+z6h9LogH/jgMgPMP8cwb5KXebhrzUUQZmA77dCv
XpSm7hL6Ln09zk76lVqWBy+gdjsRqIN1u/BJ3aOd1V3ckoSK95R1dmp61bVkHtdKgi/9RPAqTNr/
vJ8EJD0JY0aSA7FBnHbj2XRGKfmYPOmpeZCwm7XmOdr37I47g1m477KN7c2irixkjSMI30BATuuK
oP7M0tdeMQ3/6dRsAHnhUAlHQGrSEb0b43mhL4YHWgHTstYeFjpWN6Ebl/dZSs4tYG9oOeGDA2gF
4sAHQauSwnl+nJxgfxtl091E1kpuviM6Ci6elOnrdWHeENBDkc/wXGFSVUo6RzOANAT+BNnSdEhD
MC0MCl9HFDHMECKdUfPVIuok4/ve4/jf5ksB0c2h4/t6nT8WFJJw9V/WJimB6d73IoQmVAFbxIWz
u3/gQNRY2c6TIBhVUThK/4jv1EV9VmZzIe8H19AnZ8wL6+bnlzuymXZZFA/IfavgNBJPWA3BcuWa
PoS5NQkp8aRhxIsIabxS5ClDEPr7Plwp7yaRZ1BkXNj/396RRcvSr81SuyI5UhiyFKg36fbFCM0z
ianJwmyuRkTZ+nBYGCQt8KYDXb7cOkoUamC3Qri8/XsifwiI9j424DLw0dzaFjnxxPr3/78b3MRZ
ZUH+AtZEwwr5JSiLBCqx41RE7+ko47SwngSYm9c7OQPogIJ/09aMv7M9IyNvvjKErW299yOJD8Dh
92ga+8Ml5DzvEwAhvxis1nhAW8mypgvQJzwpYO/KH/iNxW1seTJQNeiCYn8xThz4L/zLYkvQiFz8
aI5NRTGrxf6IFV7IqQ9BP3q+HcSmmugNVO/pP5HJpOd4e/jw3Hju4S8NyyEiVEk/KJXzOHm2nyVU
JUlWf9o17uj3oUKJkXrzbvUnV+IU2Dweq4edRfK3tojEleomvtthVLohfU5AF7cig2MCq/ll0WIn
QN+jx/zEnYYFptcdN9VNAqeQQ3Umx6Ii+UWhgiT3xZMZV2P48j2/zx8koyzVrMH+Fh0rNy3H70Ol
xwG6gUKUxjXbtW1FVM0vpCcCHL0fMndDKC02/lVCfZgSWyJZxsWY5B/i6oyBexOV4J24F/HBBqMx
cs+ywojxg5bY5VtUhch4crWM++ky+sBr08q/5OnlzMxdiFAkVjTsqfncmv4oAKS/jsY7EOfKgsvd
LuGlTQDcNzNIuOIdnC4kruPEUXmPpB8cmKOdQlXz+0MaWS4gGqwWMqEGTpr/vmNWj0khA4x3/hQ2
tKMtIYmn4awXwVSkDV+n803UIwN0Nt4iWSEJqiCyZO8eGVp0WgOdtDRJ7qDPp2TG2m2EDQyFdZZ6
WGZtAJkg6XpbpJOQRF2jDwwrbow1uZMSWR+KwKXUWWzmQjG1OFh7uiHrMxLmZwYx+NasKY4pimTI
PfEJCBvZTHSDUCzYNZoBAdoQpAAARogjOJFeTuAn/XY0xQBYOZyfMjh/SRJPOfGSPVP8rmeKm3fe
XeQi0twP12Wn4K+ZtZ1kN3w/+WlmX8bK61C/U0gQjK18bDiEmoF3uZhUyiX1PEFvKyAzXOck0tP/
rmGZ4SBVbxHHhSfj9p13uwnM1BnAWlVKKQYz+2ozTeblXHD9KrfD+ydgCxbRhwkAx6ABjJcQAUXk
ckSWMn1gdEVq4U7hfUECQoHSRZ8FcxJmtTPVIJb4lD2cE7CQdhCSee4+rV9Z2DqW+NzJXUH+syQp
0RfmPN2192Jumm5LpoYk5eHbh+dKOeaVZGNJv8Sry+GUgIzE9yIw8GpkFfQs1oqxBD2YTcOFPNVm
mI9/taLCHZ5igyyMIhAZqQwsP5nBRaH8QmU/9Qry+HKCtH4VonIiUYSINqQWHqv8wheT2eROs/C2
4Blt4JPU33w5mxCT+CLGapFmUymq22JtybxcPoG+EBH+pc+ZKbFhjjFz6DIhZ8UE0FnFI62aXZ7K
nYWvzWU0kPRrVXxTIDqrsW8OoxuOTAMpM6W5/5N+2EiLm2hkalpJeWgO3+fLwkSe1LzKvWatO2UR
gRMzgrL3gC2zkBd3vycSjjRxlAMJCIAhO7/teEFae6kjDt1wNmKEuBptWTXd7gzcUeaSkLrBK0WI
ALC1WpoulpS1L/NQReEdAkGZPCWLXw+pVVCv626wbOl2E60zuWrKAmpjI3K9ZZcwK+qZvhfmeuKl
bqVqTRHijLRSvG/7HtR9wOhAXEUmRKNSD2kZsyFxejTBXTKT4KLO3G881B2yu18lKKdE4LJnf34l
CA0xFtjhNooYNJwidHh1ucBEgLTVDwrdSzZ9IFZzRBWvu3XndXf0BnKKgY7xN4R4n2fmUJTYpzCR
0FVq82TxkyMeo2QWbNg/HcspLwUrrBl47VKqrOxX29mDu1y7XqsC1cVXpGhUh9mI+Y2gmp7c40w7
WB+P6ZGk8Jo6JzE2j4pl2ogxf4aTI2pW9OCsJn+LP9PzDvV3V1Z6wd2XYdE3GifvmGiK+3N1VmF0
wdspms9y9/o46BU3Js7P6ZW2ZhTZMdRX69pTDmZb40C8o9iTQEncwFcH5nzPA9ZZOcxzVY5LEJQc
7ivYingDr8Bvwe8KfJp6BBPUOV8ABXyDRNZmN2sGa+pcJiNXAkXN1dJLP6qmCGQ36TJMDIs8l2qe
tyMXc5a0BBakKN10ri1DfYoo3yDzzva4DC0HvMr1qidM+aQ/ZpPfqzNLrBXSNlAZtgKRKqT55j1L
twiSE3E02+gAM3lgGqK4QjhpOdwbefUSSGSkN60zLjHk7GY5UsMkcJ/v81syHN0pCgNX580DoYQa
tckA6XvpZ2cHxzDdH6iMiCyL8Ldcy4/ymxsBq9UW7tKduClfUit2GNv6xzY7DGWrBTnM4BYVfI3e
24K/WdGzVBJydvY8AzxkjMRH99mHcKBycXQAlLmXdoPAKDCrK9rMAE97RWOGPIOF/A35D+SkMrcG
ps+rkBr9pPWZQnXqUONTyoAO0L1B58mbQX9uA5XmOZLD5p1toE6JtrC/pkVHhcMQPL+SauLw88b6
rvIqfmzecenAmlNwwDFCbNG8W8aIaFPZNqCkW/qfbeQBCpBbiv94e6tGczgJXgb1n5YC/o7kwUAe
7GwcRRcvVFruFpy1L+jzb+YhbOWDvSWwS8o7Rgw7UY7Jj7Tz6hVV+3Zq3ADQeX+cV2Ixm6kih21a
cTguTTuuQ3S3TocoPw1leCgBBdLTXjEE+pQWyo8ud+LNh9rxWxlTlBSdin3BKfLKBgYzmWN+Q3ZK
eFochRZEA3514ePa47FHQybRvaeSluh06WGzVvRB3pTObeIbWZp7szumXgORkfDRoNEqOHpUP6iU
Gx0Y4UY2MKYLgp0BgPWYwXdY/HG7qrp/FPZU/BT/RLw9t1bMxoL/GNYBcs4IQD1Ft42uyMB2c+Kt
otwRLRy5VxIIp+nlqimNLlIjVRUZi+/fiW8DvEsWONM3fCoiAnu+rK/tnanLuvktYnF1LAztm/fr
MpL+eRtm94AIfX8XX2V4Bku5Q0GiouIsMZJMTKTYCeni2Y/3fzaNg4kIuD0A7oMjF6Oz2g9S25Xh
Hfd3YBGxQot9whUczAp7eHDijd4Bg6ks3BUIij0AfyhKzJGfSGDJg2d4iPr0ZNy/PY5jMYINGz/e
ZMT66k0WhroWkG2il117peiaY7h7/sISjq0stwoi5hRfR8UM7FLB43keDkWJekPZle7K8DUuASOn
Cm6iR+8o6Lepa9OgD+s0MASSvNJf8905hWOuvrqb3tbdm7WXU5YUd0506FY/dHjumGElcgLe8ucp
b5mz+PHnJkmDEeCwDa7aSPvOL9+wQO9g3UQLZMzVaCDwUMldBDYuzzJHHn0oGSi3IMxXnhYlY2V6
cqbywceIXk0baboh+y6NtmxV02en+2AyVcpDeiLkSX2rG+dSHWN8IjzIA1bMS7mHIKqiWPyFcHIb
BdecAYa/l9Aubzhif2lzncTVXIfbFzS0XHTzid40B32yqaEb2HD8PslVIcy94CRWwI+aduZriaBN
ucdoYT/vnzmZ3e4RRTLz7UiB5GW6aqvB4DRMYQjq/zXfkHEwRMrsL2wBL0p7ICFTNqevho4hZWLd
RunuVFa1zBVfaECUA9hz6rj9d5rmTLvoJfFHkNBWgBth+Va9YbyA05Azz110bUNs1v69qz7cPVtG
CYvRnKbU/RUJdIqB36SvPkIhv5waNC+HZLwrRe9dbuJHIdNTsLYYayiNXcSazl4dQ4m6O0DM1ZDf
qxwQT1A6/eTSkv9UZQGu/gbszMF4/8nGUnI10G9/fZpCLRTvJbog6llahkz/Xxe4/kV0sCYSFi74
8YXfe2VYDQyVbHDV3suSR0viFsi0ClhuvE+75iGesPcHpF/4jrIjoNdpbTusP/8p5bQP0VaUF5E1
gUPmgiXy1Tj8Zqc7xpw0n0ZUBefMnGvnYvDAoAe8EJdFPTIDWAM7XhnLrwbu1XrwtdglZkOzyBBR
GZFHjDUP50/RJdOGxK0PjW+htKZykDtpgk9RIsmPyDfmQHV4b/kHFOvXp4MPhhw1nMuo1z95WPG3
EIb02/2s5FlLq6C5wbMug0NQiK0P0REsfX2r7Z105cRo56gsSo4Vi7ksZ0jf8TnJWmToLh/9cMzr
H9Xx/Tfd5NXfeSR0QPNk2JMAMwAAo8/EVVZzdPfC4ccUjDcmNmlIl8LB5hDNBKMPyvzSAX7WXt/G
dK7EMG7odEvmYpi1RWIUQ2On65hUMI7MpmMotpSte+IpsvGfpWkKT6eEgd0zoPL1h/K2SdbmVh1+
2/xgIDp8YQ01ktZNgcwKJb/Pa8xNRCI4S9wokHaWlKx/+8mZl+RePNwRAjuIz4jA6ECSVm7abRxD
0kHCb122k+H+YtSfIjKVoj+TVwrAFgH8XcUZN0ySxmcDYxv1mvDirJ/FEt64NM4GFc8FTjfzmvFW
4OgmScLKdlKGUXCFuuHFusJnxUNie7b1+J9+5BLkuJxcxsA0mfpnn+xDlGn5/PBkgtofn07wUy+q
rFqzR9p8XmoN9GPtdU37iGZwX7GZZaQMc2V1Mn2aVtoEVDsosxPBr8jgvGxC/+zZpXKBFXbGOQ1T
XEO38ilu8VYDG8OUvpCEBAyaX/REGMQG2HA7VBarlaA9T9IEWEDQGSJJhJhmuau6Bc5Gi2sL1NsT
Jm6OTyQ+AFrAEDTc9w8ChULmDI8m6ke3IcfU3ZIdtKzF8NfecUZp4ulGGvsrjaECpdBGIVqrej4Q
na5aRGASHULzgT0/k8xzZ7vRDLS1B+JPvfuPzKTViRqb5U4K7fJ4jyuuX2U05m5vUQiNh/WCq2NM
7LMyXSv9VQZ7vhFp1X/vn1BQ3TieGVl7qHxitlTAS/MuERzPzNCW2+NeQfRWK/h3JRVEX5gckYJl
oY5pT8gFfRjJI+C/bTISk4tBEeWx+KoW6B2WHvjiq5R6yWHMuPkemETfMBBaOQ66WLQ+8lbY1yvJ
+0S69XRUg3Nm3UAkKgtl46jiK9jTWJCbW+B2RMPqHz3R+N/Z/5n4GBUE/Qwz5alM28ARP5npyF+N
uRg+UW4dtEaklAjGkRK8hQruYAR1ZTp8YfyObUgCgxS/UngTODtuentL3oei/5UuOD+szRlj0ikm
dy4zrKzx7VtR33cOGQaOAqhgmqeHbNZs1KDv/o6WC6/Z3rdc9Ft/1lgyh84/eZpJkZ2tMOj9cihJ
prrM4a5iSMdXJVSP8w3YcQZRkw5XBd3ZljYblHymdwkg/IVnVJI0LApXE3e02boYmuYWMqrYO5zi
f5MYvhhv8bsZimEdw0J0wfIpvC6WFKpNd/pprKUEeG+hH0LLANXCzBcW3Tn/5DhgJHs1UHRtP6gg
NEyFjgjxO7hF6xrzKACbTwCXMIOoEWmHNJbEIYKeEohXbvZqwerOmpCjjgIkmM/WC6dGtEL31nnR
q3Im4qwjbSNVrngEgJmN0UNZQHciDiJ2xHqeFaJYpSKM1+zSQxtVQ7io4196BjI4x2HqLFXK5zj+
Shj/GAupWfB6DhTItMzcPXuUm5yGRO8rsCFUEIlF5YCMqnWquqbYmwBecWAZKZVKgFEMpYHFGpQe
4Jd08FlsJMthQwsF6A1iQkQtMffkG2gF7JsLRDp27mYInMuVGTmjDwgdsMNSnuWLG1udEX63Nx6b
GuwAWMDZ+q7mMMiBIUlsSvVpEDnMROfan8BNb9FEOd6Hmq3cOfE7WlxubLE2FmJxUo/8G9gGJTDK
y49PwF4QI+krF1TDNGtEmbl/PYSQOTd6zNNLaVpeo1TseBRUjWl29EVWtRBZeOdi3dzQiBA4+tR8
TQWoSUu+BM8E0fi/KWTO1LwFM7OCJ23eQtCTMqyhm8HAOAyuOujMfAWCgEdwwIzUtFJJ2YgKF9rL
fSqUs9dJHNcC6Py/j7vraKtcVuuin0loabmk7kBB1KhdgGBw2/m1F37oF29qTYN74BEZi4P79KbT
qthrEhL2QsNZeIgMWltkf+z6YqouqJlB84S9LFx/veoYmwpxl0DGDR8eZx/eHDsPttnc4nP1Q9Rw
XHVXw1h4YmMHGRhMoVjv7LZIDA57qsV1FEqvuWTopFiAJPY6pKKzvCvP+4RGfwexzYF086M+Ij0f
V9HYhsqLVUNrA9kov4yicWsyK3cdaVl/yp2iHFiCZ3DwZUoxacHU0asJURxoJDHeANEbEhs+V5l/
A6g8gMTuGEzW2X1UayPmLHCN8dm9gdFPlbd/C52pP0frEQPd9QUuvnRyHlfK4YOgSB32yjTrS63I
2WzuA0Er3USJSym7Z3PZ/8rccKNUTG85P9t5xIfaY9fBklRX03zYEfQpZx2FGwxzdiS17hjZ8lzy
BmmhWzJlUtFn7J/5zSD9l5jDBWzHl2LWd2IApIgFWFEqkxkU1p/3TAzTkQVaCl0YISKIYrJWn2/9
bZI6jcFoyXnx/CYMJFTjPjKnJUDRx4/x1Mg6Vhx6i07qqK5AUARdV7lLLzlIDNMgP8WakovTtLQZ
3Rai7KGhZN18NHbB7oxD6XuxzDyFfGJxCvRuMH85v4Axk+gJqW+27+3yfor3lpd9YV5vOWcX0uGC
9wXOCnqmsmSt0bUkfOxlaySk9zkrxjbjRCxafQLY7r4tVsKuJm/VKVf2hEWFi65pYdscFSfq+vCh
AZBuUcMcjAdCgN1vX1GiLQXiKHDC3HXio3vq/IA2vCuWutqraGxjE5KpqdOJzP2ygKEswQ/b+F+K
ouRlk1FfkoBOUpABNueHDFultZMcJZlcxjHG5ZGIy86oTzDv5UlW3wNkCfBRRuCeyGwMVYB6PyDd
meW1MBXBLwBMpjzzxy0S0YSNL+HRm4hy7eJXCnryb2U+hXaT2q7Uuv9YdFtElZGFc2ohDDgPJKvi
Z3bzHvS3aEp336QOp/lBA0wseUUt830ZdjFKI4BwJM0K/CWYehqzvW1yZjKL/lRx+yDznrtcFQ/k
oKSyy+5GaGlEgjSfaJCf1vkcqas+sHqvunBa/95phUdSe70TzWt+3+/Xx28sYi5LjMp8nRxEuhGH
tI5tLPoOEGOYALFdZP25bTP5yOVOEiTh7F4/BxvBi5pdrQytdprDQpgmrhkyaT89Lqu/wdX2x7Cd
7UHLtu/y5mIG4kJGTlKjjTMRzWzBIx+qdmUHDt0WYjMNQhJeudeoE6+hmLwgf74P9dnuEkgvSd44
yFHvAnbT5izhWsewNQG+eecxCP3/7/AkeLuTS0QkTinng86GXAtx97dnQBgv6AwdMom2lj2ynar2
cVZ1mYpTrXnB48O1URYj4Khuqf7VxDo5cNO1L6zDjY9EbXkhusCVOOzOHUt+XwuWdAnf9V0GkZEv
LARuLWPlwlm9U46TwsqsTrDgtz0Lqi5ch+rZQIaANA5uZTpdV7q1OhDdFQax48ZIcxIpsApdAqNQ
bJVf2uxjLBEsRKkrx5KlD5D/6OsLHFpVSxRtq75nFUmgK1TLPNHrnqCtPL4A8G8l2cIvt6qLNEF7
LJUCA3Wq8BpJO3L2U1u75QRsNioy3RSIi6j0KONUBTSMvxF1Ozuick30sCNvTKUjTlTF4fO7h6mO
i6ax6dPAznJ0zGZyTO6jJQV+diOn266UulvJ+1bCnKHUzSdLjQirGuCOJ32GwTzBBGYB1zMZRG7f
lxa3CSPrP0HJWoZ8BhJUBPuEhvai+y82qQ5yGiKVL4UQSs9BUtp/PCnzriz4ZoyM+sf5h6F20tTy
sR7J3PuFKo6TFwXuviuTbvdSOYPgtvW1mhO4hTQouX/mljt+P/iPKQwy3MFGxbY3hwYlfDsvCMpV
8jfBfyhEXiErRKgpnfZz+K+/dJusW0smF4vT+oii2Z+5fq5qU97rOKerbIOfhlB7qGSg1V3KZLKx
Zk76if8H26A7aCmhhwW8Udww8eATKZDAXfDEI+b+rgKL/LYq5mkFJrRBMsIoeCSIPYg+efd8Osft
X/cXz1j7fEB/DfFuB00awoFZ2Vt+ylYvogpBlBKkjPJU85Ce4d8jbWMSzDN2lOZjeIGKsxFQe6E8
Vpzfb3BaAhB5JQeBWFsmL+ZUglcIS83CWvZXLXemoGG9dvpNa2EMvILBb/MjPOkpmiMfGFqKBPFm
tXnUdLxQaSyJ/yqQMDN5vt4+GUyyIUtR+C3kvNYkMx6cQtkYrRcLvISlohnPrGStoHnecAAVA1UD
ZRPTLo3V06uJFYFXT1W5SPHBZcTtX1+Zh9BDaNdpio9ErqY6SCUILB0L6AegL3I9ndCibe0e2i6P
M6pSb43feuq4pnFZaK/UPu74czFaHwDGOciS8QBiroaBwPeEeGJ4EqO361YtJad4GthoPf/Cb0Cg
otSCaQdI3l7SCDxDX9RdP6HowgdB1ifGVVHrCus2iCEVewbfXmZhoq+l02Hq+v2PbBoqFaYMD/yP
TQh48suoeS1POJhIZw07fgOvbbg9ylkdvD8W+XXHDhAiQkXyi0PeGv0NDM4BO7fqxmJo3ngM5uyd
WhNExongnjFddcLG4MlQWdJSZNfqDesgV0CjMjzg3Jn1BvaA8C2296mR0m6njZFAO0bOrrvz3ZFC
94XypJM9O33ijw3MzSThqCAaSBaGQ+B0thTRGP0ZGwJ9G2tLF8ILbV1QQP/NusiXI4I035Byz6m2
wJp0n1RF5FqwpEGGV9e/C8PljvH2sP+A0S/UKXJNElxTS6oM+bx3BVbO24cSG7m0/59j0vBc6OoA
mYvoGlYXkzQ/blj5VDcctl+eQnppdcVZvu1B5jQFsfNlDLyqZy87RO+O55AsWjb2CqMjVDGfMRvr
d0mOSNPJiFfDMWM9PWkz+Rd9POpeuYuh9/9XKmaOJnsnhyv6p8bU54mw+uUQjgL5BfmoEnegpJ4U
+VO2fy3t/6EMTD+PMrzWLLdJOPmioxywWcCRohEPq/P+YI0ilVWglBDBPKUcfXwNvCVv52PxRvex
lAf9DKkRrJlDu3lcZ+p9EwnNFAlbA+qu4v55F8G5GcbCjTPB5IRNnVCQw8eT33Vh7UVcyfRbTHrr
iYlhOvd8zumK9tTS1wnSNMhGvKsOyUOG/SW3QhSC5YTLl8aEu+Pj3Hp9GrwmUuMzMJDLvuy7dPsc
Iqw5J0eVjt5aqjsCJnzdED8xXKHqLLrVmHLFcOdse29ErIKTbsVFy8Oasa9GOW9ePh6YigdM1PhX
tYYNzqPPgv2oWJYMofob/ieUWga5Htmt1DaDrOrY+ptLBYt7TLhFHp49KXzu686c9oIJkoJl8PpV
XmyWQ+LItb+c89nJmQdb1DQUExjH3uUDSzdJvAtZRpUNXpFrTy6UZXLZWMQw/3JXg9s0edu1cfhJ
SXQrkpuKP6cEzG5dCYKvIyAIQminxVuKaYGim3olSNh21wACHm8laSN1f8S5io5Wc5BCWhN8fKvc
t2MZztXQ+u7e5iAMKvAsIKEqEwh4wn4MBosVaKdO60bwhsbKRqX548W4hlo9qN0waz2OEDCpACaQ
dqh7hzbnNj7Q+dgP0ODwz0/0gzbdrNCP0wGLhMlZpF8p0S2UK5/oXvutcbrgZgP/IlnmInydLzfq
MBzJxO3uLBZap5QOblu2ry2JJE4IOosivq+tVexAZmkrUx6R8XUYGVrCaMmtPdIa4J7BI02px17S
IUBoGHbYcRgqzoh9yL3iDvajrlk2l9Y9lSvAa8trPXdX2M1FNfJAYqQOkHwZ3CilrHISYNA1e321
CZFqrhdNhzcvV15o0wjwf+93TkMNzLpPQqAqK+Vc4eor5gBHirwisOrmONG7dGgM8e6yHOf10S6d
2vCRJ2Gc+Br9iQe48XLsp1WmlZk7E5NwljYnTbD+Kph82Zdeao+J1B0w3m4lVeNHtAomG+TQGiDu
8Decnqg+/e+/ojcnzcBc1h8tLgYchWRFeiOQpsjaNwFb6g8+oO7b+s/QcgTJ64bAFOqCEwHGsz/k
RkWAkwWtOD914yfJJsoRkUSRrhy8xJOV4Xv6onE6SL8bDEr/htkYAai9xP09Y/L3ud+jMeVewylT
NlK9MQzrCKmaqM+Vi1+nMzzH38toNQ3WjviEWfab4Oo10GBLEJ4w2/3zymoQpV5Zedl0a2P3L8nl
TBUUXdiFNsOjfuUEv8BBjgrduminNKxZkQHuMDhwO9hvAHeKbDwod5liJ84xj/Lvqg9oI7ToE8L2
rWhGNhbcXyTyG/6EccgfB95g1ZyEIflBkJh8/Boz94YA9ZmYfl6YfL57nyTRrT7BrLXfj6hDHRGZ
i13De/9QNdLemedr6bIXpkIdjVFbkyQT6aeRJm0I4Uwial1OEAG5E4o4y6YeaXYzUZzXdiEWoe3m
fdQD35vd1PFQahKBHfzh3pOHUHr33sWTL5pFUQbluDnyYZoQrMcrzsEfANa0DR0zSAeAONMZzES4
ikODrD00ZWKyWyQMnjjr7CzgqzeeLVo+YbBp9E6sQ69hsKegOK6+bYHl50wrD6l72JOG7Vjtqxrv
DODshlTn74nJ/x7mWEbAnxjfx8qRlq+GiXydwWCPvVcRMFbhPaXguXGlzj1phyFpVBZDqANpKrXA
C1GNZgyIUZh0TbFRwPloQEhRqY4Oew+XbkgrAHFsm+D60gPKe4Wuud3TD+jS6arTnF6dqjEoCbku
LMmczBH2lL2ff2PufIZNg/oV0gBEgHNqT0iZ5HBtDM3lXfmgwfiK0WMbzew6LcjPwUGyRuRWa/oh
Q66ZVV8jCE9C88wnsULTn9fNm+H7r6rxdlUfKNpRQaiInIkAOHwhS5FirbVVxcJ5I0PlbNAfTX7N
4xMhIe5kaVQly9DQt/JHuOAYO9jzWcYTLzO8f1AO5UGcqOUOguPZSm5WBMWYcCQwGT7EULb21Ed7
8n1zmf6vy1fFudKTX2hrsuHbPtUCC0KB0P9v4NGhWxR6CFQQhbu1/W+gZ1XxfusA3TeF81N9rDSY
ga4FPowC4LuzkQZs2ykdEByUlUfDiQnJLYxHM/vvH9BTATQrlQ87aNbHCjiKOh8pr/AQUB1gMfFQ
vCUlFjs+PsoD8qRBYjmkVGvx3z2sSkCFuxOn5abhwrUUAdceNP2gVAiE7VWYIi+2whDFnBLo14zW
AzWp68flrqCHg8lJ7d7UlI2zparP0QUzk5vZEZ45/FeLzkg8nWPUKFVHGqS3UT4JA8RVjbiuBz4R
bEgx66FQY+fXg1ZAPmSe3S98VH4m56YCPOd3JXJ3hLWt7zaBGLbClNiBb0gT1v8qrBwIPd6iL58e
oJCeyC8Z/Ii7P6Xckdvrb56XA5OAGyUBKJBVeqzPQ02EhjeBF5x6geemtPcR66Kqa+D2zz3iRIRp
FC+wpFsAafQOrUXK/0eRSdzMbxVFEEqeRthoVpwjfDZwL8BnIwMePk+/vcbDimVU18AXOBoO+Nfp
J6CESy+OVQkKh8XX+DyZftFpZPNwp+Q6Thyi23XHg8zRilsHjEFskBHkBRDQ8XrkOF0CSLxsEt9t
mzOdIk95RpYp8NazBgPRBsTpEY3xWLLeHIeMz8vEPO7vxtDwMHGTGaHTflc8SI12walSR/4QtmJI
cUiQkciBVXmKu5UzlDuABLztTY1xAXPlXesWvD4g/4LtP3Sqc1yC0b3Ww1c1f6YVLVFwI68zIf7B
Zu3eUOkkDpPnVll6gw3XrVCY04Ar8EHEX8dJLRJeZL9Rmgi99dtNdhDTES8ktrHaoTP5S1N3cjuo
wJqec25rbIAfAXAMP7TFEJLi8hshbIsknYdvLo5x8yhbX94bvAg/3nwy9YRemoHowahYuk0i5mJc
n7IuR5aqHf0IOw63nPS/EOHPk9QmI06aza0fejo6Bhv/+r+FAf8ABiUteij+9DLUTVG6g9OJY9H1
5zuLUGWwUmo4WaEpcSxuMrC+PpMwFrxLHaViVfV9EbRX4ytMaA80LDyGYsmkfhImkSAFmJ8Z+vMt
quU2HxOKQ9UP7Fb+PBo+QTA8EI5WktjjTVH4+45dd5JK+egzqCdXGk5TycwnHIRc+7ASg4c7xukK
tGfES6OSasuu3OqeHZJdQ29THSN58InFIvcqLR26W2pJGbgWgaltaK6ziku8Vtj/7yl5miam1NHG
5VLNwi/HhVLQa44+nNNHbgt9ZqMp9Ln7hjY93y7VcI4ccfeZqmaH2BrQN/M7IvEvTmcAm0x6pZEq
ERBiVT6KPqBUAN5EDX/nowSBRQoCcYX7Z1uS7XguB+LrwzYo/md4Hf55zGPJ85lLTl1SYNy7Z+Nu
nHE1psAboeYrxkJIW9cFSWkxfcoM+Bz19fnEWiXcUyF4+/VwdhCzTw7ezDfEnR/amc91PqRPcx8q
+08PnLSsbxX88X6SORETir/CMMvPGQWUJDBSabrMa0f/D2p7JQGtc5UJqodRbxYm789dECtWWRW8
+djN3gVfWl25N7lWCPhdzsj55zcU8tSVQSGH3BHVFjt5MkRqW6k6OB6HOyYp7Rbd/wtX//n5ras8
Ws6QOGjuyhKy/4Hhbx1u9ZbND+BmTUTygNenrnpWOyTAjsuVucVHP9Mnx64l8oxotwf9RylKkWJG
7zhZeU6i32DQm3sXPP7z/FOywe+aJwZCjKaAB6cRuvDVBK2iSWswaxyqDqMGr9tWE293bQgFx6Z5
PB/qmgx4iWEDO9WHTC5+N26yAGYV4ogYfTbprh0V/Eu4RrnoHaFi5gaoVplwwbPTSV+56aPcw5bN
ebH3aLwzO6COUP+dgPB0ClFbbtYyTKc+89qX0Y79x0bAVyhX0xAeDskPArYqr6/tNDaWCBHHJeUs
5KLPS9o7vDkYHdaDkjMQHSNldrhGIAlC7UHI5fANUeGkEuxkb7ughQczNMR+sduqiO503dtsok9J
IwuY/jce4+f34hOijHQkaouKZNDU0eGFy/LwFXnqFWEA0SrFb6U/8iFo/SECfTtr3HYS62B8C2Xb
MkGhfgRXftqURA8051s9e3suYtoCK6aOcezWjJi1yg5n0w08robzV5yB107mYfLUL3gfleANFjNl
W5iOrzaWT8NjN2bNwbeIPHlz9CBJCKujUr9DjSG10T/bUYNJFPRat6OtX6XOra2F0iDFEoHL3np9
NPHRoEuMGo7GykXa9uw8P91SNs7/zA12Qagw099W9miNW4cjEVObb1sH68AfgS5BdLxRgTkOSzit
78HDsCV/hNeMZJ6VBURmBpxqnTou+UzvO2NbDucVxezvno48lG8znK17Y4OjV8DEWvik52RphhPL
vFbNbQ1WtWEftIqxba7WRJgzBoMWTPm2iOaj6zBZUvWAUwrWuljzgqRVUnLQP7iI9T3cmpWeh4oS
VoihyyDRy1Mf/+n+iEb+Rh/b2tcaD7dSvP+DBPxImHQgwPWRgo5kzsj/NfFAfmC/w6qDom77U++4
Qkb2Fsy+GEp27qC+1N0ppa3Ok94NwQhmiqkkVkiSf4lOmisu6D1nhav91ymq0AlL8GvgJpKw54y1
p5stPUNnh7wp6FYrLUfTydYjQrRBefjSiLwI9ITWbVp3V4hXL1LLrB6OuEaeNOzRGG0J90vkOchi
Sb6dU6eJvS+f/CMFWjHhnzTs5gsSvHMCs9OhE/eh7GI4t8zzESDLzom98P3Z5RFuLgizCsUYmb+L
D/YhuN9bZEuUldO/DBaKzXaw+Q1QvdJ+aLpueHSlUUosMEP/1ZXSO7BMSqK0F2SI0MPnJHVNFkWj
vsvow7LdXI85SE2HDqpZnNlRQZMGlnMDQH/cMJ4PAN1QHa9ACx58yrZAhx2VQETJKW1klsRYxcBo
D1JVyS+TK3vC+mg6Q2sVlm1i+VTzPvuJQPZ+Ybn0j5L6Ab0Xyqr5jTzDNQ/5zU2XUi8aH3ktXcs/
mXcwI93iw3UY0Qzbtm5rgm9zasgcbs6f4F3Kpze3I7WqepjG298WxCTGWCOzUpFb4YN64yBV8V5E
lV+IsGKhlUYd5OM1dVpDPpb9j6QPJCet5TaqQhFZ5n/G7rmD18qZsIOrDsL3O3Zou3tsaNZMNDMB
1e9NIP3UyjqDBMHtucB1aTnT6Nwa3roP+R7zU32HvNbWmV4yVEYjgSCs7trsjzrchtiCGX0clD/W
gBPUK58HGcOaoL+k4dkQ7pjctn5hsPy5ty0eDdT31nyB8JQgRTDXY1NFsVkGGHdJtpe3zO5Ln0Gf
fLQod/3VbIrFCxep4gCT9pfJIDhABky8xSlUcpaXmEXEmhCkv4G1s8pdj5qEM2vL3pAlX3r8Wbrp
pjuh7reCeXB6ZKlxi3F0ng5B33D73014SoHxc7QkhR2pKNtFWpzWq3vKUofOQ5ZlraX8YF6/CHaS
2F+gD1BfBSnPSDcTh7vqcrEjQTw9qCuWPBIscbqULdpe1Hqz6t+nqtPGiQHeFYol/KJk0cEqYSn9
1qiP4QtG6W3cbTsKE6WrDNRs8toi9ZYyRtbcOMuNuQ7SSmzwRWpnhNbNkzsaefk697g+pItKc4u6
crDhgkPP+v9cyo/Qy4MfOewbAsDQcCmh8xwgamEnk7MWJXgwYQhAM4dqpQTot82La33PFWqkX+c6
pP6BN6nf787aLCq+HM8exTKAdVPXPAZvpR7X/F73WeVtRJCzLb4YRWSWHQ7IvD1JKWNl8h3Jf9Q8
qSduGjyZ82mPyoP4A7GOWrRkKKUgWf7DLbTO1KN77s7W3LHIS+Z+XdkqduiqBpzeOhLXFB/5+ZKE
4MfCMXXYnDFgLyLzF4GwNC02QvNQHaPMOG9ZWc9UmFEQ3KsIg4idum5f00xSKDS6wF9JhB5l2zhU
o1WJQJ0M49N9ciObEACrERaom4IlJT+4TgBKMJQkXclbk6lbF1WPcVhV81g0M+mICriBLsV0puvW
Uv74OoHlNPSnYyI3fw4mZx3sqdV7djp/ADG4vVGBzglySWOeJMSluctd+IJb2IP2TKO13RMHL+ag
5AjyhQDp62gvO8Vz5A7a4Vl69op4oSLsL5KZybacyFdnxFCBhOdSxtB7LnbfBJKHyYD4ftiJSi5p
8h6lbjHx+eQF+HROCxpQWoD/HG3N+Y7O0mrCb4z8N6qeuQihMB37KNcsDWCmlY1Y7fxwtm0iiWtA
ncnyXbqdsyGcTE2hgeKdoYIRf1rbilMmXYww8GWYHBj6oUldt2IIayKS/hRvZY+9aaxLq8z86fuD
wTEM7nmil2uuG1m7YEUXAYEf/aCAittahtgkpFRngS3SNw6ii37NOu/teBZH+Kln5Q2HBsE1UgPc
8swId9K3MzXNyb16Vs0F65cdVhVqrz625CjuA9ZEgoRkfxLA97yqTp5Bgf/ZhuoLdoK+izgpk0S4
A4n6hWy7IgvuCLyXt0M8HfuMf4dTiuGo+/461pOX3FgAgsVV1v+OBwJcAAYKJv+nF5QHpQO9m7nt
pfm/LsJ97Vmt6vOD8lg1vRxaKP45cnMToH2b+I26MC1DUM5URUkjYA4MAZvYijwqE2JMli+puBYI
4qw+KuD+seg/qAqBR3dGhJoogLCCKSqy/TqAJdVRKQ91htq2mrzIcWITcFUExucFxL6msnsQnzjv
g7hOUNOkHqjkFgFINvryJJB+np+FOXNUL/IwjZfjfZ5FZUD1exgbLUf67cWuUgvd2hhrbZ2AOgrj
m8ub9zi3ldB0CaemXwt1xWiTerRWqrqanIawTRS2GbmaJb5nPdRicSfrRP4SQDfcT4GwW3l7bj1P
mElRauMorO7s3dRg3jErlvcus9ryc+ep6LHjEXGIiktWiPqguKKp2BIlP2QAIVvos8VqorqQhEgK
z6W3grJMYahNo+Yk6RdyludDtAUNaOIPLxEtPYC5uiFxHjI33g/5FP3zOllRapB8G1j3onynf/UN
W1UNi6n1ThqQJkZYzkf7qIkh/vYFktceXWJi1MdSJjepmawD0yAl7Lgyk8IMVga8ujt7bz4MTX9R
n4lRbasFcv8EMU5RF8GRl2biUT1bi8WQYS367JpNYAzVDSmTAJ68hnuHQbwAYvz7/kklsG1PYK2V
JmQrEAE3vicVW2lJAEdglfG7sHD06MvSgQha+Ani0/PWwZnrZr8JiqAuWkzQ4RPs5hpBBCln6LOS
HtTxQYVsRedPJ+GHujZNKsg61C3LfGeXTaaBM/JglkspXM570jM108ET35pfCjiXQ9xPUhNiOtsj
2rc4vCzYcIKFa+wDMqGZiqEMaJjk0U5lpPjYo5PtsEIpvpkVfGszjGgbGHMk8fpCQbNSNIKBgKbS
BF/Oa9O4s12yRVFXuKDKD2ptBL6cyNwaeJekNJnOF8+g6BNx4g+SGqlVtCgrYlllH6vlDpv6Zq5Q
sGG1Aa76q4hEDbSjUwOhTtre8H1Lw6KD0Y0e/jyQCC5efLRVOYEOhR6SrxrUy6Sb2uMUtS1epths
aZWJpIKvR7G2tRlmBlA6oQjXreE1J/GiqTUPXdVC2A0N1+uIYLd5wvuXxp7m/6I/CAxdTFBiMOf8
TmsCau30XKp9d1gEqnf7MpWE1TO40uGN027qsNT+YtpO7wSye8fN5x4NLjqsfIEL4aCbultJCDd0
qRmkFCz14wjAzLmwoRrviBrwq7UT+AnPnqVxB9zetMwjuhK2APZdO11zV/Lt55jB5/et2zEkMkh+
YyzP8bab2mZjSn0AaStGnWOmN3uZmItpdMDA52YFLtCSkITMmeSVswpALD0SJtmrQez3eK7amQze
KIci134J3UbhnP5KWczczw5nosUbsrai46cp+K48oZpza5hAa3wxC9OvHpGID2rZ0g2W4f9+EvW/
95sMg3j9GoXYkrnSzL26p8HV5NIBt55kqgVVpb9G00e6B6gSoViTpmhGpE033yADFzzEMJg7Xnya
sv6T9CZFHdx/KJSgB20thIxHO1rER0v+PByTUnLtMKEpnuWVzTW+GWBN3Go5ocwx1a9mDrFR5vkF
L01xzghMv0X0O8ZuIc49JHTmVHba6L/UZB/kj/NHxAvBCdmNwidM48xjon2PdzpkvpnKcJp2gLns
Dl54O4Gsx5ucFxumiLLASdZviTWaVlm00xEMWs6rEOec+2YNUD+iKXv2QUCFExbUzstTCEfG3pqK
I1udb8vSk4iVEx1SqL4WoNrqYr43USw7/3fsfuS7y1ElAsCBqb9bHzgpxzez8LWacMv69XLvKPCr
qp0Uap+nRWN7tkx8deG4iffW3vuGntAYapfVnw7uyccwHY5AyfcG7iCrqP9JRJAfqyqQBIOZ+6ty
3XrTtnedQxUcxVeD4+voaQbcDKynQty980PZVxiwrgWCf7oxFsmOveLmsWNGrcDqcpQVOaG46Y3N
fkoKfSXMYvJXJ2YNMYV9u3M5PU1oSagr5ik6SMyA7Hh5gWrzDI/kpee+wu7wrgcm60+NjudmXfzy
szHLSlXg2rjKockF4d5jjfBUFzOI+6Ivyp69ml93odWF+zmaX6aKUPOeYkAOKy3FnV5tG/nsy+vN
wGptnn/9unZ+UFf84/EjVKfhRBNaxGAToGS3LrjbBG0lAz+sq5r3A+EFuG7kW8cTw7ijzI3Yvmyj
N9HzUzjSNqej+Aog1jTfkQIx0KNLBrvajF1RCr/mz3OjE8DUYdNc18NxGZKLBdqxSE3BU4uMNIhb
mcVJl8slQ7uGcAUT1XybD0KG7lffgVBJCxdhzDkvmrN7RXZ+25LeQEoOhnUCF2IqLGoyx1xnQJOX
8pkNbU0PB9ve/l5bw8esJayZTdzAfgVOuuUn+GUeFi/1hSoXzaYCN0WGVPqo6HMX8zz3B2aTmwdd
j+FfjHXe2jAalGOnZNS5f08TMwvDyC8vOyjAjuzHTFZFMrkZaPgcGm1S+BOuGCrLTQueo8gO5Psa
YxEtZJ04YKrBH+cBiCGo64qWIWl9ln/q7keIGb+YUrahu7ZnSgJazBX5fuMOhC3fBPgG6EgmQcZ1
I+neJp/dehLkW/dAHe7DgYMv3rrAEQT+m9uOsBSKDtXrthM0PziQeLUVWiEAz5gOpgqkPxvdGP2W
VSQ1FH943XZRYxOIyh6if9FyO9kmqEayh3kHrtL3fOW4IbaH9PW7EfZLdCPIVP8bwO74lUoavEfA
0s/3gsNrCfqXlBA7A6fw7rcjwZC9z+8hlomVve8ime14jvT6FpUPk2Yg9YRGk9CDmhPMkgh9fknn
v0UCla5Q9/ngf8mbi1VtEzdCGdK+7Sj/jH+z194VPIdpf9KHs22EK84uR1JSoBE1jowVZT2+Ync7
6y+DfoIVEoLnuTDmKDjtX39Eizp+z9fBYALfbh1mFF3DfvoQssd5LxCKKLS5tZwE5nASXVNYqKFT
gV8VCXgd6hz6MKluDVfONXN1AvZ3m6B9a22i9zkZHoKa1X8/xF17JTJ270zwPnPjEr/zlj1jRELZ
3iGQBpGE2dhAcO/2z5GPQC6PmBwcW5+pd7sVVDqIBNgnqGKz4e3FfyNV5KaRG0cjuluIimid3rlW
V0luiKSKSYkAthHNLntmsfhMH38ZlA+Uv7MlLd5xTfQLc7tNX3yKY8V8fUwFbhL+Ndubs4mu2pNh
c8sHrQ4EOBzFbaSVKxQAQrh2FbaxJeVNlojqLiSsK9Hx1t9XruVU7smzCLkSeTFXQo7+KirwLfKB
lDwYZ4vBDUq16yDV55pp8WfOZeEiem9X9Z/fjdPBYMvtDrpo1P+4rPufunpBKoKhUph7JMvxyg/K
zyy7JDIEn/7Xp65CkljxIhiPyE182Ke/mLXFNGEJMbNzyoYM8EbHstKS2uzG6PmiOpJDyp50vMgx
EPJDKRf2G/z8aF84+48TbJPsre2LUqsYidi0Noq2U01ZlWU6xcy01Mwqg+jFSkWUcG2SX2XbLiBp
Qnd5zUishAe0w+7oBhbhNl0e3HI60epFDO+tBhSET60BA3qr0Ylh3nV4K7kjxTPOQVtuIo+ort+m
VYiZmWhyfwXAt1aas0jqRwTX3smvqgpQfkGd2p7rHr+nXJtXL4d3T40QbEz6PcJnqKjHdWe+XPxU
AbVOzJPWrwaIFVl4heF3sUeUcNY3fE9CXeR1ZNA1KCKAtMcfneVeCZkc6OydGmiWop/sxNnCSumC
LNzegr3Tx1zzX3us87q9qY6T6/g9VfWhx0q/SoT0HazAezafjEkex5oXVemiis+8ZNatHJ20gs/X
AYyF7FFodn4XsmdwItfTpYUjxG1gtLqqRvB9TMYyhQvkTNEPciKIOUV/t/Whglqtvvyu91sH2Yji
lxOgM1ANtrs9MG21Uv/A6m3xkJfLiw0kMdZmTjPWnlwZporClS6T83Dd0+UceqjkwoEngW/KMlLN
y1Wcm+JW/hBxjqEzJjMM142v5PZ6j/5pu1NWrn18g7Y3lr+14ho2YyeWzmIvsq4WJi0VgHPvRn4i
qE08H8XcfLFcOx57OAZqFfpaXtD4m742VZFbNI8XQwJ2sLxGZk5bkJAEe6Hhyffd/g8UH+1rLy+3
F7HkjXaVhMidrVf2Zx2IVi8RFMRBRA6LWig8/Xx/3YCvkGnw94IpEud6jKNBUAD9OV2FincV9gPt
vu1ovVbkJ0AY7J2TgMrr/jtOuphr/eeFM3e5IH1njCZCKlkMg/28RD257EEBrgupUMez/MviBDFY
OwAlW63J4Ln4DT4PnrVyGU9auNu0oAoSDge9znjEwRjL0k7Y03fWOrlJ+jyALgq9Jmh23f+GoCFN
qwSiIO3K9UTGr8ycYnnWACngqdSd5vPS7YfJSJuThwqsHpPA35ZSQZX6SsCfc5nuV1iOv5vj2JAI
3jo9CEOaE/zXTL5KOF/5EMcX3mkh/JzdPzJH972Ef/eNmSGAKk3txNrEu1MsJ0fTB1nKzsQlTAPB
grA9DXNJcfaETBKPpLbVwVIQu+QPtFcDlVdRGpiQfVMjdBbA+zUd5CzgYhvAibLIpXlLKfYXl5vY
2eIXVqKC1hfEXAxjrHMWBv3ElCfP3aXuE4UxpA4XRTwv1tWgeOOzKg7il00zcgYvWQA7Cm31MMvp
9B101sBCgbHPEp3VcwYP1r6/a+WIE6E3ZFiuktwKZ/ZJSBwGmTgvEC07NuD/+Y7oS4QOpUJmR+Gx
Y+hc/3a3KzEvCbsMkbxsN+yhqoycNWGSZXOta7FY0ksGsEUVqyiegVf7csQCr+r2jcKBmJk3Yifs
UYoMmD6mhMFX4nG+ujGu5ZU6RsMWOpnL8WSmwjdyuXJYvmhmYlmPqM1hQm7uNzOnBK/XKggK84W9
MFNauOLsQARC0p/LaRWfL5wPSsuAOL9owcpEAJjkiePwQ1hQKuPqNx7hd/la+amIE+27CwHjq/rH
8QqtJz/zNRflZPu1/aW4ysaUQy45ZmcmBmQNfJBAZHfnAL0qCrFn0KjFc9kB6eRf7zrJXwuw7gK9
L7eB+e2ogHlDnHjON+7YZqiPeCAy8fcnOkrIflN+MD0eeNpMcD/j3cjyQVjsDdhVbNHHObld3L7L
n1xK62mTIZJJhazMji8d/rtkV/tJ+RfkBaWcSLsMSmhZMESh1p+5hEHe+ZdC9R80vspjoOoeU5uP
AnZDzRt8mzEC/Tu4hUaZm+PGhOlJlSyUoi58cEGbCxS+GW2lXzG4ypshOZORplXCTtR8jQys+U34
bGR4qNnvTe6tkxOjaTobf8+VjdTR3x+3FDX0ZG7CHCDz7HlcLNCRDyvRK1s7ax7EfyXwp0/fngxB
7dmHhtPvJdXDd1TCb00KmG4Cm9um+0Rpi1pOMuyCNk9WP+GLNv6BvJVOkfPMfYco/kvDUN2wcc5I
m5C4wBVYaF4S8uCVSpZhEt375WoMi7AkzPIWAt1ELA/WUMLb1CcSYhcMLLVkbPannSogh5ijmyxy
QJFifyAPgDe8iijiXjr1AUcB37sex5K8MlEZUa1dRoIXavd9deMZtzSZpithgGMstTaSc2LMRw1t
omd0zROOsIbuJsMMVbtq+9asQDoWrAXQjlGPj6CuBCBhI+mMDDJBfAPZ2ZZIIdbjjeVHjBs8jxJK
E0axNOEqxZ6jsT+li7PYs5LXMV4S5+j42EvZiBOrHro14faz1tRLJWqeYIJrv3lt6/0g9Gk8ccGp
066E4zRiq/rJeemoWibWF7ZJdJGu8pQSj6r06x9i8Yb5OuHIDFQZECP9FRoIBro2e5ugY9rj2nWm
TpkB3HKnGcIXYzunHhNBrl245SHyOWDqBFKD98Y8VUSA2zkS9zgAXMHNPLpYX39ZpW4l1VHpCp+U
pszhmDHIz6dpvvAPtqN01Bp67lMemUoOAYynCkriC+m+ZJ1h3e89Vdyo5g48MnJYAdaqhvSaHSRY
VxovgW5093mkL8RLzyBBgh+XlyRRVkDl+AdYRFjCYQq36PK8Ocdx8EHHIR8kl8arUu29E3JJItml
QQ5O1Eh/L+Y/a7g1cuyn0mMhMoQXaZWr5U6LDv//Nqgd+zJSsbdMkMoiSpWUIhz8ZXJTh3tl33LU
gS1amCY5kGyO5ZYuiswaq+8gnVAf0RXPrFtx7KcoRvoLdqrxYKJulrVNLUeL6i3vhP9JhGVTscFd
RAwcw9EvKhEdNt47CVSej6E3TcbAbi2yy8XuCMniI13u2WgUBviPlQW8nPkvT59MUiGe03Dj0cUs
OF/doh6kyaONqIOAKy31FpGCjHUGCUmVcVYOFVirUKhUOE9xe45SfJ74i7hHsEQ5V/wVAHEmhVFy
41e71ln5aPLl03ZWmAx3jQHILfPlcDINWq0FQBIFb8dL8pcGVC7zH854GVruE/SnHFg8Sq4/wicV
MlzMvHfwfTzi7Nrmgzn4FjGwPfLEUYAJ2cAPiSsaWQSch08Z2egz0XhnfupOp9Y4RZCpHF3sq0sV
o9Wc6uI0NIURczVMkQ9IyiRjnvHYRVXo3/OFWSgqkH5ArnoqKrDJZo3ZykVR4pYd6KgwC13lHmxI
efaNgM1A5d3yMpyyHO9B13a4R0M6Tlg7KGjjKg1Pr/s5pEikndN7fUCKpS1e7t8uFA+DvzTDwlUc
KO1tXm9oaJEswF4vIHHJmY1xsycOFkwg5b3um0SygVaNhXYyihpaEhJdZljtoOZp+qpp0Ve4IfF+
FrNgSiCKVCici9MPAnzA6jTxtDXn8Twcy864DS2KzrYimN3v6En82QBXcx9UZee9mYCTd7r9F3IY
a0Oj7FQLxsNFLelw/zZVikuh+9QkI/I+ZOR3hV4ExmDPlXN/2bTKkVmdr0YCVP3MfYKD0EFyHUoG
SWrJUB5cdYj9kWsKoUzJx+lQILGCzVNY6WeQjeLM7pcb9gWV8y5gmUGg+aVR9YpS6r8bprTy0Sht
hPvHhTKV5IiSKU0n8np3bbELGClp6kXFy+gDbMK4cZpXG9AaqZYj8e2nbzocqTwjEJ0R1hoJOSGe
U02mfn9mMxhcK2Jz6ZFQmXfykUG8ir/WJZvrcUvmEhYgZ4A/S9+pCybbj3MFfJLdml3jCF4HPNrj
TyMewzwOl2nFKDZmdoWNDDr1Bt9ACiBrTUlUloEVQ2j0ibeKxCgX8fjfOPMdqb3WM/dMkBxt95C8
6Exa2e7QJVo4+EsUQfvbE2i30E2jMbZRPuCi1kTeQk92YkNlU+K94Cq1Isa1JY2bMZYHF9BInKpY
vQydFhH+A2+vmb08mxhplFNMX7jKE7avkycxopu9HfbFX/t4aPxjSUiR+FtytZnJInLbXxHGHplW
+yXz8WXPCeJEpKZyvG+GPzL89wYklnHdvhEqwoYQ7bV2XpsfL+zZdQhNIi9iXp2xoZ3/xW28lio3
hdsAUUakXpqu7HuPhzyLhbHbqdRuAIL1C3k5gnWbTk4wsn/VFpeog62gn1WnyyzHtIkQjuY4UXKt
74BQekboM9zTSIoGDaTExFsxu1slllzj6n22NH6EwS+DIycqsP8gB15DN6f7wTColWFIjRRTNQaJ
iZZ002ZjI5DUQCRB672PmLF8tbPMl5QztY8NlrbHGeWAlPa/mNEuAVMI/2j3vMDtjFJZ6yYoYkXJ
14P5MweUDR7TRuD52JrVnIuvTEOX9u772mxfBQqUUGVcYHXXnEh86Lf3JHRxcGky4VXiQeFh/HrM
IjePrwor+ips/WMyHrWbC+2RGU3UYmccRVLHGtZi2AMmXswbuUDVFsViAmVpu/evN0rlfwGwzUjl
O4WDg9WKS/iN1MyCeLPaCVUxPAq7DRfPfujmvOuPnnLIhY1KnzT+ECsGW1ZqLc0R6Vo1HvlyvArP
gXaYCA8YuUKohUH4pIVR3mceXubc5vpdBsghT5N93qWq6oYRXIyh4qZIYIh0Mgcg/44cUCgL1ya3
PiGH3dPJ9Rp/MFvIN0uuV1VOVM2JubQmBQAQKgcpADY7FwQ1RS277Fk1waxv6a6BQwTPAME29kyz
Ke75ppbcRusHOSGG7GJD/Jl7MIRHvRgLUNoRC0eCUeCnPUFI4Y6zegpGvN2F2bF2JbIA14W1T5LT
XY1EAGIT3ruuWvMc2ZvNll4b/XwQe3u2Yt53ipQBvhAU0anM9UDujxLJx7k3xG3UdVREOFzIJ5+Q
rWvHCv1LqX/a5sZ1kE60DTGplD+56xSH2Psk9/1vRXRzZ6sCSRJWHTwVcdUhRd4RcKltl5cTJAzc
DwJXDalv9Mbzp6zxkZ/oTLGLuxBtlHYhtmTvtH5jFY6TqqADFiotPNqntwP7wDjAkxvbqA5JwXen
xD37Fx89KVv1VDHiPwXVSkLdhXxY7qWUr2I023xVh7i7wV5t8wucYSPOq1xoHb0ddtVRuvvsdj2E
3qKNx2FAZf5kLLl6xhxjt3kIGPCzTAuDtKYhXoN1ZUkgGsPVw2iqnn6wvjksvTdp5rbchBZpielK
ipfdtNMu2ZIXLhcC8EUJS8mr9yCVwNlwN+xPp3maz1t40Up1gwmQRP7Js7UzEHKuOdwAFMam3DBO
xoZKSCmpZ9w5yCeLlaRe3MyLGtT1Qkj0bu3Env9McJfZIxse6vD/5u3lsmx64mpxSOkFOimYaYDy
n63fO9UP4Hkb5beg7HRs+mF4aReSlE1W0hwHJUVZuVXLo6xT+uuQalShlWmepDxKQP+RDGZMGqhh
6m7sIFFuODOPPUI42ve/L9DkO3oFqhvYfwoC3JsQm8/T2FtqKN79iPHWXo0geAfYrsd3YXOsLyTM
/hnjosNIIfnXXRYZ/UKUUQ1HMUj+ztR410RiKTdTIlxclRGcSvwyjUbbwsGVbLzKZxUmsTEiXq5b
qm2Z67pNufWHdKq8NTDj1KU7hLPOoYEkTSw82fJCb0eVRxmDlD7hKezZ4bBJ+z5vm/ifTZtp3Wt1
tSPX79Osi6TB9YZggthqs1Et2K6ADzAdeVsZRJYg3Whm5L2tc+/ESnBKG0ox0qANwa6D91R309Vf
mB0vDjfWC7rmz2IZlQjPMWcOAWW29vbMsnTazJO+8VGXNkXAhjnEH80S/pgs5QNGOVpvk7lo9OSK
2YZ+bitGzj3gL8FhXWfcyIkkQAhLqB7KeEXyMpczJ72UKEmaGK69BWwg84JNXyHBTbP5Y0ydSYV/
ZunRf+JYGGK9yOfIVyRl5BHXLimhzyNSIofz1Ed/kS/YnOHJhufS7AsRrQ6FYowlNdZbcpYeQDhs
pnQFDv/TLcZgw8IK9tpGrCgUnVhyF81/eWrx39mdeZCJM47How1R2IjfXCVVT3X2t16boXzmPuTx
Ab2QXHJrYofN6peSH88jZ97PMrMCwVUXq8QE6dqxe+HHEuSWp0BnXSybuiEx7Yo6mMFAXUwadp3/
xu+4F0fGXc+/Ot3PjRSjEKnIGmv6/yozHi+2CfSAeX02ldffLZPFf7XEH6yLicjisSGXmujGRdtV
d7pBENTXainYQOAJDXb0Ua7uYo2XvmhiLV0pL/6txrvhdpHOT5S9JP3O8MFCa38mmjGDs2997z00
G91viZJP+PtpTg0K8LxJ98kcVvlmzKeqH9WexUCFlM/zNLOfyOrDHPRLzX+wxtBMgpqRfcYLz+cR
NEIzuA+K2FmtgrDbVMvf0krdW9RWv5gdzvURsVMXCpKuskOXCuJYNIMrwIe7LvYdumjEhLuok72g
LgeRigAPSG3MtGNG6LnYp8rezLCHwOxiwqvenhcTS0CoyzQigb8U1KvHVNgFHTNQqkGYPh0/hq/j
tSNJ9c22mKGkV8KnrXXf7SqZK+6FdHE2RpYk63ro6qiH+0XX9AkHflHV0fxe2+RYclvtVEiyIPSh
j7Ksl5OYTg/L3IcQPdyjNlCLRuR8XXloNUJg6jO5L/liUn8MNHZpD9qIneuINbr2V4wCAk6Z44jV
q7SZkOpiUHIGzN9EtKd/1PLZ81dpbNzUK2x5bkK1s1YA3mmo6r84YDSnB/pq9Ypry3yHQknISBMc
u8jji1xfig7OwI6eb/YgbEGT/Y8eOA+euj7CRY1Qs4CmqUJTr1Q3gvsWZTtisve9AzqNrnWQrL51
VOa1rbJpvxx4hdVvjRRUXKM5pz7YcXJp7I6T9H8QzsFo1OOJkI/FsVHKT7rzovjVxnIdKzmcsaWp
VLVJwIkUuJW/2CucUznLb89oUVAIpjNqKS+cx4QNETKQE/lo50vZA9Sd7DJmyOf8C9T7/7YuQbVW
fiHh8wDlT/SuGRl5sCWf+7bxwomDmFaN3lCFDiBFD8aN29qBl4piMsKK3s9+9UWVk2nKPmzm4tO/
L78xoHVdRae62yxndfcgi5YjMocEO5YE7MyOrXGs6s0751+JA0foVuVRCwQLIOBJRUMfCHv6pGk6
S0BYy6IihJhIADaIL/Y/Q3wJDB7tWqQkqQHkIyaAXBQIfX1MJco9WQFe9Et9NnTXMMJYpPyHnmcW
cI2lNE/WB1E9erwmXkuOg2leMi4pFXiza4buo9MqiQ6ZzJZkp1GrnerHV5Ik7Ah3Tni0xdz02VD2
UrcuX0FnNMpbthtnixT+ADO+mORgLZLbJQsX2ecB9lHtm1L+k1P5rpkLoUYOVi4Zjh62LENzT+Uv
ssv8PxzMqaYqJgxNno53zQUaNElJEd+g5xXmeDsah/gzxZfCmZ8fseSipPE1/cvJMBxDRCsMNuLM
hJd5s5StCzhVXFD/MZp8WOPQG5fXrI4bNE+p5oXn2ISfaGF7SHujQkjMkMJyJn2IMxmjrwt6F4Y0
AxaQDd4W/6dUyqnqXQFmCm6tVB/mcmfqTD42DgNa0SiuZR+07XVbJifDbEPvkcmk1Sp0k//rLH7Q
Z34/upEEDTvCuec0Z5yRo6wfrhWP1/EElmDpptDX+GAiVAwegFPo1wwVDzNZya1iv0mCVFOYv0bj
PhmJm2SXA9f3LYb6lkx4c+9sZ5e6SXLvnJjjVzrpg0Ljqbi5dp8L6VirxiiF3uoKftIqLyGfsiTd
pC9hEjNE1vO4/oEjeduNwzoLssCo/VF/c2eJahogMt8b3e3WTmUdTtDKPjCaERdtwTWkn7JBC4/h
n2xw7kJp6jJDclrTEnBZtPCOMTKTWNhDFg6PD9qOhU5LiaJAF3K1eYet45/iS7Ahlh0LJjkyJ2V2
rshwxCOPKoQ54ch+JbIVfL+5h4T2JaDCj19EY/kDjDAAS+pqzmfv8N05zhn++a3Y9sjrNYv7bU5J
5Qrtq/mhZG0/yq4O2TIoglVgAxI/BR3I+5M8LuerDHokwLdNonDmpSCBIJO0N+hnNVROfeUVbLur
I5e4kCGij3vbB2YlvTtWubQI0/gzs1G22n8OaYV3SL+tGLIRveCrKxbnsaazMIPG1onRjuDXTcWe
Sup4qHEPpaLW4VqGciL7ULvZ4aBKQfe6CZqYRbomukikd+UwnS0EC13be04cJ64GxKslRjRGJANW
eqpG+cZeMmagh4TgnLKXSfiaAQ2snagHAkLf0j36ch3PBr5NZl5ejVDXp1j+GdHBQx1pG155KM+n
M46eoMO7lc+vmIGe1G8QW+2d9IeHb50imYB1xrhMmlQjypboEhkzBVvZrBBiQaP6tdIo7clsmN9R
laLsj6yF9SGnpja5+hTl7oorVNemlhY+Busl1hVn31Oaky0yXoKonc1xRHvG3G7EirjUxKW9fyL5
NK9/Z2GLakw36SaVahyfMlco7yxv5gBa3zrZHuOlQ2Vx6eQbdOqxo564N6GrGaYRDA5NAUTtobi6
jpX5rSQc7jUTa3BTxzdj0vuTsU82f8fpy0LnJ4GmkikLdL+URrM4gVp9c68LUHtKtWcGv+xohAlq
nRBRGICctXQMv71fDlpWqgktHQ1mXT3cHg/r05d7FoYVbPs8tIhSozbeCz6x/Oa+gGX0/PYCKuSN
26Ni+Pitezmi+qqlt/HC7FMasqXH1XHiuEwwM71ggEQUiCUZzOJbo5w2zZoCV5Nd6CUdmL20Uloa
fbufPLcvbecjlfP68a6cSCS230PcQS96g5jqp+ItG9TERJzBCVyTSTNw59eLxYU1MMf7msV/dcGu
poME1py5Kvt6YVV0H6HVKdAlzRRPyO5x+TtHNIhTWoWPYc9IgLxuVl00j2vIL3UObwNDEih3jkUV
LZCrsb9FL71Wn3oa75FFqNTONrw4A2koT8ydt+aSO11xq0JRqW0HgBQ8QVwhiBZh6rYKlSRMctwd
9EZyaBzqXPh8TW1pF2HPom54z5X3SxKzYmYkIwrTWKSt4H6gN8k5CPG6auiCxfSatEks/cQ+gvII
UjD4S5OBEM3N9qkAobdOL9oXBS4HhkoA+dYwIiewCQ94arNPDEef+tLlIxHcLbIwmxT33tyEe5Ti
xi/Nod6BhwwJIV8qmUYXQft/e8rdXnsVFCjn4NGZTN41u67CdlSnfrG6BkhaM+IpwnWrlKMKrtNH
HOR3BdhVDkrBwspK+A+0hbELejoHCoMtdyIThk1nR4o1yOXo5pV3ozSQfSqfm5hzCLjpCRNChK/Q
6XdocZgcNyX0Eimp3Z1fHN+AC9cyAlKEm67767eeJuphr8GvQsnwcLsa8mhJvyKkyCrWBf5rJuDf
0yTWE8+M4F7b0qUZhDaNnWEULlsnHhuJ+Gh59ey6VBSYqgxKhtemgn6Pz4bXOadUxZpo8mRMacfP
XgdaFPq5KfkRYj5HqFnYA8Yw4wHkV0takE7TxPJmOyyp974YZThI3ZUe2rsHRdpGoWZq3sablJJZ
Wrc54DqDq+0TZ1KllRlibmPkyLzE/qwWlsFUlAcf4Atcy5S1oXImvLL9WADZSFB2Srh1Pmt/Phk2
Qj0qhIHhG0z/qK4IhnFkhBDwHJqHweZADFosAxLtKPBNeLIzvX9ELdkTL8Kd3hQa/ZYUkBCDxRuI
DTWfuc+AtE37Bz5vg0+p7gHNuc87aY34o2vCrNulia6XIYSKg9Yzgth3SbIe92hI5pzLX9EQ84v8
CpQWDdQwIP8BK0se8jMcfcDK1zHO0xwR6+naiLlYfq10WE/hbWzK7kNj6Ieql488OJShNb09BJeO
4Wak1/dnNfQwjmCGHR/+zrbaiiM+70su/3zrZdhdUDS5+tzuRvspOZH5SRm7qxKz/fDffzzOJd6E
03zIfhgyGX4iyIeCXxVUSIXeI3E28RyQZz1OFTLKUvnF1KRMMYnxWW0tac2MPraw0HfUfsZJ8re1
bm4WjAaF0kXBHzWRcxoFTpuUKnqSYRLMmXNwalSZG1qsAGfKmIJaEo7EwPISpVXdjv7BvUbo66XY
04ylOErUC5HJtvIH7BZvy+8Vf2DbjRAcFZ4u7FyreGUBLKmN0lYGtFJSK+EeKcfJfWB4zqRJGgbE
MIxc9OsrnYUoGVWgZFE7PI+3R4aGLPfIQ3xyGR8AqqOangZDxtqAu2BJ/vVxmKMlIVFizpyerAr5
IYKqt7dAYrKLNqAUuHCE8hGD8bt54POo7DIq7NGz6X/O5vhGXorjvDCKAtVlYlvgnk45IqcztrNu
441pNun81eN4B6okSTz23FsFd7yucDMePXYu7x//x1Pb+QojUk8i1A9Ieb7q3OV6gFqWCEC/9LEj
133XdrzpBrT6BLny77mfFTlFoSRcXHXpTsB3OWy5LBq1+VnbCJMQEYq1WuGZGxmZoTW2SqriaIrm
Ka+pjCQ1vplhi4HD0grSAnJNoJo0GJB+y5Y397jDf+k0UZzSzrvIGlsKobV6uH3qxGpWJ5DeyMMW
nM4hH+fTdLkEwN8WjdaLl6xavqaaqABrKzbYgnrp7WyAkrAS2kkiEpiXunDNlXPhoZmnHIFjokkw
lnYzCpmm1DNdS9FAcaIRlI4WwAijeRYMJ8TwKzMZV5s9KQHZ056vxeE4zinugHJIDjYkiYbnTqw0
Y1itVrkvrCKWVrXWL8Kkct72bE3g4lGn7sfN5c9xSCLCQiwHz7EeneJyE93Fm+bSs1RDB2Bw73sI
EYM1UlN77TbQ6M5UXxVvETeJc9Jy5c75pGTqr5yfeOcG6qwOCYuMTlrjYpjhVLdPNQiENjR29N5p
4VL0hoTNF+1dfkZ6rqvITFm17HiYL1vtOzS4rfnww1HZLihUT8lE31tmJBg/kfTAwc+Nt/tiaOUY
cI9zEuxr/hystuPikcS2xGe8yJ/WUbSAdkwjU61PHK50odwlYpovydDx0ja/gT5so+ay+1drfcIO
0pJvWZU07eDYpA4ZhY1JaKJtzp+Z3VfovEQSzFH6Mklv9LMMOzp7aAFxd8+UDcHNMVUPQbl84I6q
/hDtM6nf7Zol3UDLlM86SS25bTcvx8wPy1xw0VyWRrl03Wv7PZd2PI4B3ll1wut8CIENOvNiQYqC
1spCTXkyyDaFNUmt1Hi7R4V14O9/ALRoioSOWWLjdHwyuehg6t5WWuPs1wCu7onmXDq86WKROhnh
fZqltCFnT+Ihx6zb0sbLX54qQxhuMyFY8AYDn4Qfp66AvgJdQFyJOvTZkZrwUKGzDFZ2gpyP2C9R
C+80o97thUVs8jiBPTfsiYPfOJjzB8yA0Q6FN9PCfAQIeIYG8n8Cl556KDvjWSER+lsUOVTcWBKR
Vdlb3qxgY8ccZ581/hgPGvks3ahQhLBzi2hvApAmVPsJocO8G/trDE5DE/NDtcZPCTIifRKXYIzB
ilUrOp6PoVolx3nCAOQw8BWcuyGMxxfecRTz/WlyK0Y8EpQUERQIWrnZD1fYMe+7QHznXJqe8VTs
kZVbNpGmKH8vdfOVK5UddK9SVyblSs81WpsBSq6+VUKOg9BqmRkN3KaL2BPooxW7d1wYoStj7UJR
x8D4g7b4kRj5pnoaKBnAGhUjFtpJeHtVQjL7BmGyZywYRHn5efh3lA8m1YHKWLB7Kc/kw+KYFCGc
IjpVEjTeb/fMjGthCIJqCTcAa97X7esAf7cA0vNotA8U6/o7cjp0EASbCDVA/sajLZN+GgVP8Smn
1TRmTagizr5vC1HfRhlmB53jd+lU4wDlklaTTfhuLcJaA0cTIWrqlwJ8lfCAuII17ZadHWUpBNot
1ETZQqAGJpYoa/mK1Alz4mvDzduoWuAutzYWsJCL3ISvPXqDgPe1KJlxb097lnv73OHGVp+MiM4X
Fjp8FoVdGV1mS3agTXnviR/5Up2+4te5vYHSxKU2pfo7gk6XezGuH6L/ct5VOmBMgoJwyVppRa8H
g739bNJuu9iXz43XkwLAf2/DmvJMUWGYX+suV+dOpBpCY4sFTl6mf7ske2ctgdsWnWusrnZt4ULj
l/nFWV3kbW3UAVHJorTGGfgxrtmsuaazzMX8VZJxWdfRY2Kv6uqUMv3yuD85x5nFV8beDpRLBWeN
AVCBbBVbw1cfrmkRptS3h2vh9hVzRe5HGrnbb3XtPqcAR2mOKfaXYnuvci3a8BGGupv3pUEf+0iH
JeYZz7kSmhcLBCV6peBK0cz2Tr5MU8DK5Td5AoRvAxTcwDHitaXNFviQVhRnD0GwUGp17Mg9lJ3n
sCiAIDbk10kIgE8T5XgG6q51V5j9giU/ljbIHR6/p7I6RxkSAnSD8e3OKobv7R3CRmkZW4H9vNHV
NG5FxaMiRc+6VLZB+QcLM1fyoU1efjl4PtoyyS6KsPcs1b5WUd4Nq76gBf2uzoojo7DHClVmLOTi
xf/6XirJJcGI4SPuWsswgIATJDEyRXx2/Dt7heTQqXdtdT+2L2TXKhvkbwMbss/zRqa624u6cejJ
qt53ZGBMLFEjCjEpv7NKQDG9z2UfmrcJt9JSKLN2VzybYBsM+2rgeUNgVjPcU9j0uaZPqvufiLTa
dcJszqOc6TSUaYqEWgvGsFNDOeXjwMHuay7cyKh7ggaRbRGlEOQ/3a3p4JqlxidFPKdDUbwn5gAl
KkGtTrlQM0UjT5GFVi3apu3pang1MQWYbwAkYE/PLdAbWAX2LagACksRSqdQKAVrNjsykJXhwnLP
QWYBi4cJmaMutcMza5DGZEO66p/63hZtLg9pmCmhbm0klzZnR4ZlcQnEZAW/H8d2JlZxSUf8VYYH
KWth/8mGwjzz4Limd9VdXVCwEzhHsf9637eerndZZfMF19JX0ZWzsEAEgvy+5rfTHktvlIEE708n
2+puOuLqdxpeMUaqbo1a8dtnG9EdTotYzdkzq9pMeQ5jUwCGUto68HPw4f47kD9clOL6U+cTm78d
vec5MyItLf4rXMDl718d6AUi92DoiX+VsULJwh8zcBnzT7KfaG1VrsMOCezGYCbWd94ehTDj7jb/
cJ8K1LyKXCIzq9ok8x0ybPR5D7LSqeU302xsaAKMNlrmmCiNubVAaJqCi9fLAnsYh3ULi60sfP+t
t+l4DLPV7qA0IaLDQ5q9kviIYHFDtmIPqYxwBD0Y26SSESMO3oalvKRAVLGLMmKi4D360aZETyq5
GjmdP3Dkrn+B1J3HF5niZ8XXxrAiMhb1TiZP/mxy18WoX7qcc0da1zc+kQ1M5p8Ixvv2XFOIMTN3
5pxzaUyeddjnw2r+nKyTBqo+BbxoMtpgWxYbmqRgrN8sNMDmaM7gcBkToONmuLNmSRuiR0FBuKjN
hcnLSqFI5j1DfYTCF2m6IHA/zR4oCsgT0F+KxyBZH//8VWq5wJKIMvLwOQak7DlPZopO+kzNJ3Wa
f6V37ox9cMNtHYstmxri5q2kO5TfzirqF+omD1YnXg0iL/3k6nn9JgMQnGZGuxESTb4/lM97d1X8
PxUOuSKmxcRKmpusxZSvma6IH9pLKLWF552xG8BGIOKFYqDuXgS0nwQ2pAC/kMxy+bcOKkFA3ucc
Zxj5x8WAoZLGmwYZSouoyda71Wl6FcpALszbszUIF52q5QNAaEGkE+AWhrENMUTOnHsOzSouDSY/
C4dbn2hP5qUqOa4U1vY+f2A06tFETil94/3Zq01eI5ElX7wh8UCmsdy8dNiEbYkmceZqm9PDTDZ5
IZ5QXoAsnPSQkLTw0ULv/D8mZOaNrohF8XATwNz0pp9KxNEErswD8cFheQ0Tf6UImxCK9bkmmcT9
95CqrSZaIqlOiqY8YWyy3zVhCC8xietEGBWFLm0zolnkobkvza5AC9vohP248g8ALTWKIhtDIzcm
QHQjmy4K/zHvfrjjMyr3IVxjs5YKlQ8BMJN5W9SbES4txJ+EITXDT9archhY35zEReBTQXzsEMTP
bEMN/rgI1XQmsCmq6qu8puEIAERMsK3wZkm+9Gbbs0XCJI3hYv5pkFUJRxaTiwEjdfUt/RxLZOut
TR8FRSv4+IZs6fbRd/Wth26a1SNYQ7vMTxwpSULC5zd7hNf3tWpG8aa6OgwcaJyw9GWl92ESLuvE
mDUY4YtYx7SIGJyMmCP45JAV3V1/1LQI+em+uu4o8iF1o76mGUdLZmDP2DDRRCLYK8gtarayzcmM
8ps7d9YvsFkp9VDqwr3skPtukIMxLNETEnDweejBlg1/oaQMcwGr3VQybXmgKu4lhI+nwGtcPLlu
gKWre0nFtGsoiuZsC/zC6X67ghRjK6BYHdalSWjHVuFf++/5p4MFCfnNYvK8m5xpfCFPi2FW4SWy
kKo+8zco+EyZ6up7ymKw7MGnWnFMVIj3AdwzhApTKrYZnsBQlzOjrYI26OboHuNi9ZwEzN04R4IB
pV3m/Gp+4v0UU23PXwGyRwzIqKNrkY3V68lGY+raE7yqDpnQ5YsC/2LqU9FFL/dBrbfE4oRSLXGJ
LEwzdDYCENaKPquyjr7Xzb/pw2sbRCqfZtTIqVvdyn8cQtzydgbBRMSpo17S+RMWlYR9tFZBEZqI
8vFyM2AAuxQtjadBK0xOmCg/3jVkvdOANTZPMvGGh6GHt09OYff5iE+4WtxJ2Ds10QdojZOUw2ir
Jgs53UdGjeoM4gfooIBdHpZX0ImVh8sDWHOo4GT8pG35Rzqwg1GjRbi+VmwcsarSoBGZv3fw8/3Q
ZV8tZu6PdpYchEh0dS6p40UWYpo+x2MkFIwc8d2Rl+KGbfJAOUHmyS5vL+EIdHCK9EUfZ636P1/Z
Z3x0JqFFY/agQdhEJVY8BWHQBx/jd5Kary2bqpH6U8378p4u9MUR/98GXBfz2VeXnREI3gOUbc10
YlcRFTBbGWpj73pJL6A2OhmyngbQwHNkHgd00lYN6AvERfzJA1VGbhLSKx27J/CKM+iUG6iNVSed
WXVgG90mAqL81CTeMBjtDQdDEmjMIIsI9lrpKNuR5f8Z7gvrw5SDvHAH8M2ljMDxa2G8nFRXK5bz
rAuC52cFg4Ih3F6jBOyY9V2K9ApVe5uXZknAHh/s5D4BC1+ED+Huk7FHccPnYmzUqWWazkI1vyDD
NAu9LBXlSDhNViONUwJCyVFTvP2aTKHqcgyrxJfcHKZh+UcL52JRPKHmn6KmDrCO1XFKbGVvBi48
jxWnaco69br2L4lBLV1Z9B12pu+nhc37jocHxEcmeGgZL8V3gXJXrUfVHz1Xatdo45W+DEfxGcZi
irreNMtUO/fgRzO7mRT5pPbbJteGn0ZSZm/VgF0K5Fz105KosGx2zZC/Fp7vg8jMTXtCDTXLLzOm
lR/xf1rql6C4pSIOiwZ5eNKAN1WSSqyGO+XDxMPSc+GdUahw8xPX+EjNChczCllXoDey/hoG8eRg
CrNAOtkGPfpJYVs7ViEEvLpyXrKqWxhgesRFOm/9q9xGS9zr5uEcGdIXEdpA0fFjYpxwmun51eOw
EDi65KCE/1FrUg1fpOm0AI/sh1URSgk6P5XSGHemapHKcRhh3t1JxjXzW2Qjg8iae22kn0JMWl7N
lWVt4GBzqVGn+rROJRpcq5pOiiMp/WvYuBxVTZeihhGp9sTuVziEwZ7cqRuPmAyLRDsCMTtlsmYX
F81WaZ6k6RbdAzsGbdVl/ONFeRQpawS3A83tH5WVY4ISKFiPGgfUB+GBnB6OoxTW6A6GoYtyo0eV
nRu8peHyYBl5ZKU0dBpdZDcM3AyDe3bEl9K0CTY21jXVOVrxLJv9EuUrg1Wvk0uUF+ez7aPnNNjm
oQc/ZCYkGtdD0XVGjbE5lfHbgS0s/MzWU3ifftVenWo4YU7gNF0i08L79yOobW/MQMnIHHjdQM1A
yPlsAb5ix81ay6I8xJTxQw+0YaPsjiK+izwwOHLmcHoTcE1yu3xt2rD/o/OEKaGReg+rNuXS+ppO
tUPIJpJgE/UovPNSwyWpns2M4Zo7v/5iGbd8p4pKT4EY5Esnn3y92BQXvX2fWzolfYYCb5zxC7uc
Xqhha58EOqiQjxpnkesDlNVrXQnCB7iPTbUvZAN1FjN+KOsipj001NArFmL6vdPcMKP+8lnA18Pn
/erMxXXbYyot6sfqMuy+6Mx+f72FrdAxDdlT66CE8sJ+BBGApthrp/I/Ds+LJy04Mw7AEU0h6LKV
Rdx1ET9IlCMJnSFqaSm922AqKsUNBSNG4HfJvsYhHRX89LoOjUndkcxahX4vJjmTPnrQqnOuZ2s+
/26iABYVgUJ3PstKUuvjcbwuPMPsoDWHo4qNyIVPaZtxukulpQQ4q9pABTUCu+IQddE6m4GXWrvg
L4oMcWZxgmedqR4LUsroMxFl//c5nzZIiiQyRLEOeRNnzK8LHUWr9/5Ve3jP4OeGEPHPfCS5xiI7
TEMoxskk0Dn6sBpmbe9AYwS98Ih/uhiJ3RrRl13RHaWgRgAyR3TMwMz0by4INAbiBH85ZxmQ7JhX
0uYJyGqWhSt2sS8RHOzfW/nd0Kk9EIRLFfX4UvZKypXRGZYDW6TyltxMHYdOkxK2XNm1AABnamyf
0lDBRYbpt0VO/Yaus+P9+jlec+uuHIUgAxCBA8iBJVHi70bwL2KhalCxqmWlZMJO0EacdlziAqeZ
++Ue0YALlY6VbL9YqjhWRXfc42v8uaBl1xnS7jIh31B25aupk7JRDuLqK2/hQl4gvwQ1KYeZE1qi
vaxHXBSXKXDsjLf0W4BFwFrXW8DL13alCgBRK2P9pMyZRYi/K07HF+q5pRgHyLmfsaIS+dO2maq5
VnuTmsUtdPi0IWwqmuhBjD2YU8QueNYgM+QIZUew8f+qVUoXwdw+rzPsQ57oe2vqJ9dIgzYv3cXy
m5+PSBfb+YdAj3m7KWYdzKM5fcB0XOLoeYf9CeC8vcSVY0ol2fUP/r8Zdcx8JjbBcdVkvjyxv0ew
84C+9yGivaGhQgMwYSJIvTEoPIYKXbb4eZo0e1TTPWIiakngsVJiBq10rkB1jK4ga2Ln7Ahi2LTK
3Z9ctgMu91FF9Xjz24VVQC8Dxya0h7U5tjVfkyqNo0amDxwLxuWd9+3p1GMZbPFGlnIIvkOwpK0P
SDQsvheH2yDoKfnufMBTfSjOUR4LCYtzoNFFianMV8gcTXUiNvEjidWYEOc/N3mXZqo9KbyWf5+r
nGsgV9qfaz+MDqEYOo7kChh3xY7CiFEGrtuaFeL2Jn5NFr2novGx2mkbHnp4PeVbJpVEvb2rK+kF
0+CLYOEp7yGLMzd2wRN/9AZIzzYttsbjJ3d+3/uEoeRhz+tqgQt23hGG9GTQhaVoiNHvTp93NEpm
2RcXAlrou2p2Sthyugbipt17a5HhqcECKIb2McGLCLgMyyxQIf28uqN4ntVVrNDOXvMjRtReZqbk
vZEbD3dBeklwJ7lG6rT+/efPv5H/tKvy/4W8O7S7Y/ds+ezABlxQR4+xz4AQQnaB1bzCG/PDWPtT
dsU8dKz4JuhaCk9qcV6dG+M2dAnoNsLqbwkPKX+sVq5OwzmlLdZmE1IhC7w/VQB7yT6zt+bOmh4a
WOGzg7VGtMLNHlCS9LUaEYrp5xl+LUl3MZkiwvGMioK0nH/IvIcQUXia4dSHrr2BUwamxD29+hrF
DqOmZQz13kpWvKEXFPTpwjDWIoZyD92jkumv1sT4WxBZlIcYkymx2by7hl8NRXJ004pAhAIpUqIo
4j1YOuKSP7Bl0ix9LXxHraKYtcZEYREs0lEXAMlLtBpmwj9gFLAu4jGUd9T2ygMGN7dxcyJt8sdY
TVoFEp6PyzkPYmWU/rgV2aHO88aeghXvjjRfzV40N8QnREK+w3/AARbAjPGNOjTPVXaEj9P//AC5
T9ai7rrCWsjlsJHz4xQNKN/W7DsAHbtNp3EhjGXc2JuNSZecGlJVglXRRevfj4l29oe6MFdYvfOD
03ldpbSEhPHHseZ7dHxRPjAo1jwoyAaSSJJxjL/Hxbt8KZDCCAuq67LTRRmwSRPFx7rPMk8iJi7Q
wNq9Oi9Jp83h9U8/NXzudnmnRz5fW4XLT/d4Oq/iMHUiQdFJi2FFRE4X92UXWjdwpokoSDdaoFP4
IyPc+X+EM/ylSIjm7cdaqiqW4eLnVnfMSyW0riQQoUqEsRjnqts4Hj944EV2D4OHJLn1cqBJgq2f
R3ZMbYA8YEEdEzlrpmKUWdn+Ma+AUjJjlZPGFwkLShVxB9QbpJJbj1k+5qxhsZhbF/jR/YzpPMhu
PBSseK+coBFb+wi0Yfo36620ommDcrfZ3avBE4GgVhXreMNVhcZ873SJTgRsvPk/sgCBfj4DjdyP
/gd5mK9zXaAMacyzPFy3SmN447qplTw2cwI1y+q6EDgRMJkB762uSuyJ92nOkGcnX/EtN3djFdAe
2bGgLEbSogBIfZf/Ds65rw+OpdtFtzcqBTD2Z24pCTp8K0gJ53dR5hDQD1K78Mj4vMg2kTcsj2xn
LWw5tH53QetaqhKAgaxQLfE6j6aDK8Uc1MAPegPpGIeYntIW+b74DlM5JvstE9V3PZF2pUPoTc6p
QekNqT7E8uw6z1zyIWK2TWLOSrecdrsIzOtlvjL8GBJf54+77eNHEkKJZYA3LwHb3oHci+LaYH4B
NUCei4ag77kUw/PH8vM4zXdcnqiIAjOf3qUYA1fS6WEqVIKGKgHJYB6ZEf5IB8abQUKWcaTQQnyk
7wGpI157mqkkpx+5cFq/VOWnfetMc2iQyFSOluaH/PtsP9f9zHcTVZ7LzleuqKHYkldzcggeFt+j
TCoZlWNNMwyae3EKD6BGfpUVOhugiDnv4oY6itxtzs8Z824bja2eGzg5sQIscpEhKkOICpsNxmNv
CyVi52ABlbhDoEmT++VrCn9pcimRJ2xfl+S9/8n0KVUuhsDjdHlKNW/Sup5GgxkSdXBiXz01hVxa
sQsqVhnsk5Ze+H/JMtyjsH3mDez9NqmO6/jBgnqKaDV9EchFdvGBFOTwGdjBGCrfr5aopvki2bSR
o9oBJ2W3y4cXou9lIRGl2z5EWCUJEyWUwldhCknxI1JxFG0Mh2w/X93TdL8Ym1si5S4dmj2gU2p9
DurMeOZnfcUMq1AN+i0Vc8Mf0iDA2Y9i6pgK8egxs3688X6v3tWNUrcKs/Pig+qyim8auQYnznvj
dOPCnLrDAubeYQVrDx70g++xPOxZ7t0uloPSn6PMEE3RtprW0FhfCjWiQvJjyivprt0gYrJxcH1n
8suVjYi0ckLcc4TpQUrjkUgq3LTO9fl20h4uQFvBLcYzD5B8JWmGGs3tpczawWgUSgR36zwin9QY
anMVO+fJJLHl5LKBuEgXrt9VY8rqXmP6seOYgdjIlx2nzXxyIR5HsuLqDFkZP+TtnYji1WujdBW4
zET2BKEXZEbrDqh1gfvZ64q+GHbBW/cG/LSIsJbuhxCjGYjNAjos/NDAj6veZpW9q7yZ3gcd4THx
7Xm6INP76Gw1+rCmtIFiwR21mjI90oM8eGGrZQGMWYlnP7y807E+5JZKA1JazdemmQHpMHi7O/la
n/x6JX80c9mbB6qz1wqKtVcBmyYgONulZuniU2263ZQ737Lm9NLfGBfpLCi+gVJORP1cxhl4r9bT
Lpxmgj/MGhMCcoZ8nA1JxbG6t00rY/AieHFQyLQCGwd9jzRkoq0JFUiEelCahjumz2rOfgYS8Y/K
BonHM9lrMidzQi2kjzyTtYxCxKG7+VlMpC5MbNibIrnPhD/K8JMNGatrpcduF/3ofDuBHj7caPsT
1rH3F3DG03ySMKQWVlV4PPvRaGLr8ZqqL5lOeZi72d0AYnBwIbo8IG/5yVxZuJQVK9jFDOqhpYOI
1XmHp1XhYvOtgZItrjV5m/M43L8T/voRCaPjrXaNRo45VApw+Qtaa2aTEdb+VUbxlkPCgknepwLw
NaXEa/7LrhIlX/8UA2MTbVEbnDyiH3i9uAon6hJ5FKeRrao1vNweka97AXOw+emVa9mc6MYw8xy5
kaxhwGS4yfWv9lYnYsCuaysoA+NIGgV+ZacCy61OO6tki4fZ0H8bQLvqt9JRjkIlPZ4wGxTC7lmy
hfHsBruy6FrEV056l07gybcCg2JuTeAKNQcvOoxL11yxohS8kV0aZ0L7jQgKGqL94Zy2pYxWlzFh
DS+ZEJEFErjmz8GH/2g9BmSyZU8teLyKPPIB1+64HMlQgB1N+bcnv0tSNtp7+P/5S1Xx6UvtYhJv
cl+d1Cg8kVoQvZrnOV95sjUCpUd3OBFCW1gNHjgbsVokusfzAQxmbqah9272SAjkNvTcFF8hmzu6
yG/8u5XZqHxAcfk9dW13NwETqJkTx+UYx+TU4NfqXpLrJx6Oznw4iyU6Nq+vzseJ+NDJXK4CYiLy
6hmEYPkp+q51/hwUH27rHZIgqtmCii/EqDmEKNZDoAOdixdo8ID1RL3kQOYuWnzlwchO0/2QLp7+
j6TZcp83Rl1LuIGqA1xHFhGZ2MYhWUDxF/P9iccyp/xryf/YKRsMUqh6aYwjx1HpVIB6Srm8IfOJ
GwVm1uGQqiYCK+EWAhACOcH53tEMSdYzllxvD4lbnLLgm7KowQLETFy9ZJSa0RUodcGGvTEnKAHJ
smoAzWCiiMAvO5TI0pxr19goCUen60Wd/e0vyCxGEK4vrBx42MexGW70oT+U3umtqbVr7LTRhmj5
XE9hMVp02ntG1+8yN7GCydZEQi9GViK/cH9sow/n+yP8i7MT0DsL3LCrMWPlsd/Y7Yv3G6rLI1m3
b8g+/OunxaO0ofbyYQmhxKzqeiHLUNkJQqGcu4+2sgYyBwYU0G1xMTnGK9DPZMSYdLeMB1ICfzXS
/TTL/McaLXAM1yyGPVPAAC1AIEdIxGVTLLDY2U20CGamLB8Hclly0RI4X0IyaH5Ic0efYYn1RfhG
rRAz6K90EfWqacm1QYkt1emgK6j2LHeDUKHr0zYCoo2EsmQqP81FRV6q4OSA9G+W5AsJj65VGtFX
qvzBW/upB5Bm5P12kuqJF3as4lNsbSlgr9ax1MLY2LFrue39UviDPJu8x1PvSY20WpQa2kO87gmT
kho1SciUhMXRQFMWzyalvZDjQgasGCk4SYOWLD/52r5Ssv3jiRBz4M0S0tpSMQ6qM5tgWsd5rOYs
LrL9jzU4HCw6doYVJll14/yFuDboBdaVfa1Er6j4BCIeJ4GcHSLF/WBY9Yi2U393YwGQRs6vtvFU
3P9ddwaPewA57z1sEHE/QJKU4qb/zbGVZOwzERs0js1GcUTswK6XStjUDgP7jXNEWnUb167vCdPM
rqgqKXK9xwZ7DByZvpg2ZA6X1Dqq++Fj/hlqIvjJHgbG/qUoW0WehIBqQZrgAMvcyrFyZkGzkp9T
hJ2lEttNd7f/t7tdeddAiijki+xgh6tDBWfzXGNb+ugkhW8688VeWfEbja69W8sATsF3wFRRGJJX
Lgx0aZlyGgQxC6nSQRLX0D85KuNXNsI2Dx5UYy/O5AlThEVHC+Ud7rM3zIwt1jve0Pn2HBANY4qC
yz2nYcg27KqSgDJsxD6CwCWS8vUlm3+9/VW6R5zJbZAE7hjbfpujEU1ICkYjFwADPTiNuxq3v66Q
AriIGnlUWzjoi6IdugjumTf6rnlZF/J+mlDnxwvF03lQ4QLixtADpi0EemG4RHWsZhTNnhrkAOuf
BENqrAhwO+ksNj6w6XHQdQnm4D1j0PmszkqwXKwr7vCRAKQf2tetz74BnijkZZazbY3AExRDVET9
WQ04vOu7ITKm8oYMkGjTNj5YpG2eGKRbOBl/lp2NvjrI9gMXbbYfcEASPjzVf07Ia6pb/beV0hkl
76L3K+pltUB9OQpXCrtPmwwHA0MZfjIvmLovjXeehbHP/xTRWMseHU+Hnm3rpp+bXvpwTf9+WYQi
1DUqpKoztXgUkBeeidflUU0RxjiXMVTLitKdwQMX0TYJcFzGx+0nPFrdfTef6PBseGCl0qeVuU+O
kVzFZRMc+y3+wS4VqArcxLY6m7KMK4C33eMZUoTH2qJMz7IeK4uBABRKtcswpJiP7RPKqrqrY3Z7
X5sUaQLaVhHZDPNoZeFX5lcesNorbjF+iLG6vDxxjBbVAfNONl29qapx6XU2xNwrVyFSf2fYlVJ2
WEY5eCo7UaCFDhif9Vkr3QjTVRbZ9+fJs4usT8tPUDIp2JSENNVuBl/9D7d2Z++u6oHqwRubvI2n
r30eE7RahDHh6TCxvpFZtcm3UgE/ATNiA7PzEJfIRzu0UajtquFOQyWwKF6199W3Q1NN5tYTTgFi
oef3ZiL56DXXOZuEyTl9CKTPiSpTU2FLh80pDW/gO1Bu8LnfFyLzl7TXxKAXAQW61PS0kQAM9EI3
eHSy0Kpv3SFsgUKvns2CzZT9/eATM2Xl3qKGtWEpht+4AyFBNkPBNrhUD+cCYGMH53NlsDnNsN20
Eq4G3mb3NOYO0KF3js+A6+mdJJuw8b0LknfYI8br/UmR5TAIM6bvpmwPwOGcA+1iCMXaSHQ5jTS+
7vHr/0BPN4lJ6W6J1S/8t9i7QjsLMU43UZ2qs+11Rsy4ePuM3He6Q5k1rcF3fz/AwMk8IQzMp9Bt
HOl5qvFa1dmL/ECuC6azh92LuVe0eMMI6Mj2OlJ4IIWqdoefKQ8TStxOO8Ku43cYoghr69DHvrfD
DwmQPgK4xQuwefITckj7jhil05BRC9fUyglwdyonpW099r9m12eC1uElFaoTKBEE5+gwwxwFr2Jf
1NMgXeOGT92C64dJH9SaawFoxvS5Jia5EVp0zykWj7fLnxAxaMKWpz2FNs1EZj2DfrQD+tJQEmu0
JaMqhTP8/YF3pwWPiZpNf22Y2mQB7zlDEsrxjuRjeXokOY2GKmpNqNkwhZ508E90NhWWY4gjsRT4
rXuxuy9U/4gsMtS/zWX3DO+0luF3P7nMybz/o1rn86aRkd/5NJ87DOVnsDSQ0ALyE1dA00/Kza09
6PY1wFUBreT4HjnsCeAcHnxykncZF25RF689xo/kRavfA2EH3kPqxZqFXrrnT6yqa4y1p4OUvC8/
kz2wt+wstVV5nDSU5SnVxxMVWuymwPZ5c0oRN2p7qozlqwg1la+D75pt/9X7+AdYib9nmjHq+a5c
59oiHnsLOw6ZqY9jyR4B4oLvpE/eco/+h6mEsKdc8Patp4Q48rrtSYiQZ0+CCVzBZThs90CJ+IJK
plyAjECfMqCSPPsLoOnmun9fFphxtEancJEk0njNXo1gayASiaMw3Fr91AJd7miO7AoKn1YoOdQs
wm4M5siVgJZaTi/Al29rAXGkf4Y5BYWlW70vqU6puAWnP1CnTvnPrRxMLuNlsTWY3hx6bTvbCnXZ
zBZU9gwP8m4c+dWnYRP52rHiKGvOY5D6dTtu/XhIJaTt1zBxLoFoxMyay3mXxiefC3O/WMOEDSVx
ZKYWXs7+DCXFMGnIk5VgP5fZhH2GZOnvyCeumaTJolbb6ql0hi0WA+wZkqGGZjCjuHCyfV+TaUFK
JIg6VOZkHKdSinUDrbX/2/F/ps50rsVLhg1QE8Nq1mR2wmM3lLhTyiIlmwRDNqT5/v8HtIF751xL
ohs6lR7ZpnJerJrYoBxVdpCwLxNDDymni+PUK3NSCrWa/wFdj6129olNDMcAhcyHqoGOXAsoeMEj
0rurpuLBil0V6VshzdyPcexY4fvQdkmR2rY9diGyk8wVFeUcAtJcBpB8+AQ0tm/vekS5Gp6AXyAV
8dpwFICXrGhCne+1I2BTufYHUG1mTRG02hU8hdz2sXzXK3geiuJNb8FYm27b19/UBwOIRmr2PKIu
L3u32YaHJsKsRyZ6RrQXVrIIGTrRg3DxGSS5XNfEaktuyOsZ+5so38bxXPRrVZ5eDE7k8pG01Kh3
q7rcbVbz4gsmoKtjWhGj4g3c6KHe5WqixNFNmH9vSGzeRDpZAVj38iwKhCGWUBtllcCYeijOqwC6
HmGbFyWSTAkCQvmDOWUhFzog9w1w8ZeIxKaBiv4+zG97Zv0jT9GvoijYgPCDVsIXl+xPNmcvPFwC
cuI6Emm6mA/ch5yk/J3qYavrHqowd8eb2EVwb5R1JI5s4kVPfv/3vAal3BEPBTtdIEMy3yg+EDrj
E0e7yTTCZcyst1VYtzieAepFlnn/MPG+6t4GjSgStkLJW76QVMsgY7PZNCsWwO+0o62OFd9Sc2a+
WDD9vbXKkHJ5sICnXbqZjDeNo5ecQdWm6Cd+1xoHMqIdBCtfKpxXgsH6KbP3ZiSrRO/iR98PBDLU
+iow9qvSpLSTz7LPBP41ahGtSrhrzfuJ4ljpOb8gFOXsCNZpB5zTYg7CR0ztg8q1waBCWsouKMQG
NGiEqEbrAXQdpwDXosAEFo3Y1Xjz0Sk3MAmZ8iuLN6wiNZabrsWgy7d1lOhtOA2AAgROLbphXXMd
iXIFEqLehmpgiDJz9EPCnpjH5NflMM3dYmHynDD3O72m6N++ibTa6X4TmrXFhmJj+TWoQ7lB9QJc
ezaAPg5bAVlYUFfEzaCawKj1OSJXU4bi0jrV4eIMGy/Ro7dv0qXMmmGoyw/WzJuZwZ//m8xL5KYV
r1td4WX/YAuBymPTzZQQ6hox/znLRGB+jkfS6kSAgC/B0+HcTN0uikJt0NpcRIbkTAWHVznkrlFZ
eGtkZSQFWew0uxR8YGeL66NaGIdzSfrf9N3ZreppOUTHkBI1/wRnTUfxHuWqJtogFFusF5VpmGKT
bq+yhA0C5FmgUtNaShSzBBI33giAbHXXQqoIx6Zz9HaALblo/qK1qn9B/YgpIZB5H9IYVwM3glou
y12Fil5ZDS/NjjAmVB+h271Gak4jC2aKlVlGSuWfzjP+/q6MXxgD4+VEGFJXK3vOD4YnC55sIGoU
+jL4doM+G+jmxErsW1q6K+xwuCGUW24cPfEWrZiepThQNw8fHMhBlxQn1YVfTAOLq9dZnEPNIr1z
Rn1H1re/gP1UbBiEMuN6pdhK/qZWMHsG0LxRkajC5w0vY20s0gf5+gYwtR10cGOvmwIaWtly5QlQ
K21jMVQ6D9YXN9Zy4DyqnKHHkeetscJk0qp7EwsB4tW1mgDbwzthvyrv5ZcZu9aL4hilJkoH4t9V
2k6jbW5n9Zm0mpxM0TcQ2b8vshgWFEmNamiehJHzVrQSd4OevVF+IjaxQ42PjOOW9Cf9yJ2bJZJU
VdSvWyXL1AfW5fg1krjODtQjx4jvONYMub7pVKnobtNgBqWEDuuDXzqTdy5R2Z0GfqLzxhvjLSv9
opZbDE3OOS7y0P/FciodFDn+iFoB5P133RgxhyGt8Msuk8iInvdGkeVGkIfAWKRw3U6vCnOop76W
r1PEDQgwRzmY0eyAFR2ck/eTcCastD5ri1nBFY29pSOzEqAJa3i7TrYmzOpv7m3UYNonuwlFcyms
BAgDJUBwBRak6yUnUyyIgH/GViaOZpgylkbRs7fm/fN4V0ZEfx1ZYBNgi2qP/bEe5nxBJoHkBR5n
Y37dWNTZ7FwNYO34MHmhfRcGM8VzjGcot+bvqdyRFRaumkIQuefi/xJlR9AEuiC+bLXNroALr8QV
kT4mRxjXEnGiwgVwh0PqV0XWi1/ziTtDlRdeARQhNMUDHm2TWci9X1gh416OKthNYkuLBWS8qaVJ
CQ0GMaDUTg+2w+QM9470bq4rch398cm/Upv9J4MkTACGPrnJrrOz9SQ9yG9ZkS1m6YVvWt9xxvIb
f0CcbcibWRmOL82st+QT/EU8ydglNuuL79sp9Gh5vsndud5S9MAGjHW7aFo6THBExaLewbhvSNrv
KIQmX5WhsTXnV1DJ0gLmLbNoRo9r6e5JzXUCA258xgpbKwVhNeSfT44FhodFkLmQfUL/gCWc6G4v
CaiKTjpX79JOWVIplT0sit1/mx+phgwJjmnkQVVxypiAzurm1roXJ5VLXB7AeKXcx/NFLjYUNole
kC5Y9U1FfFxyh2sxJg8T1aCVKw5y8cRwBWSoBHwZc8YskdD8B7uDtcx0cEvIiSck/aTFaUfOhmWy
+OND5UhKB/XQYWXAvw240MN5r5u4C4/HT/7FcSKeEy4oHih5ILDVrnnJc37DI9pmKXZX9e1X6ulY
FgFjUh00j1P+4D0JoR4dteCg8PAdNpiIsDhQ6EdwNGtmPdGf5tL1Z9I7YxdWFKDmou9QPqvxZVqc
7ocOeRlqYMpBRLhe81qD9BUunyK2HS04G0/h3cghEm3oJxnjpoVsGb+QDqEcYctB8wvsU+aeyHbY
iTHxLjntXGEXS8pTcdnW3QcFZariaig3c2aucOG6vvrkd/r2RnTDIfeNynu8pYH3JZ+W0uzR+WRu
Kr0VkTuql83rfZslomJLPDVjizY2dYzULq/2Fl+1eqBS4wAMXAw2JeS07tLhnWU/rij7FCq7k2cV
/QCEiYx/7rZCh/rrXMJHseovL7c4Q0opFpELO08sos9/NbDiCg5BMB9zrKaHvnAgB9XWHj3qS1l5
uPXjQtgkJMsZrYUjalAWuX/eWXKQuZVzK/gLLaGfejYaLiB6Oluqq7ZHwpzTyijWSzm0H7maPTeB
Hg/eFw40ZirBDeMq3Utvu8VX6Ev0l+bvpIN7cq207pyRnKocDM+lpM5Nyh01WsDDmT7Y6hHdvakY
RiE83RU/uXo4GXC8i33a/kEVUriZRTPhAfPfnrgv70rs32TQXoHItsRGn1oiSwIxFtdKhG65yWQm
OWU4YHjQlise1F8rGoQzWgbevNKUEkC3ANhEEsdvdVeAA+f9sDofpthgCOTK585rs/nLj/eDokTv
H/mrIVTxTxoXmYzpD76pf3oCbjKLkxjMMg14a7nF+VPjkpcZfOYBMK3624Q6ZJ2hV4YzqTSs2N/b
9/dG6XrzUS+gj8qOH8CGeJcXrGwjCGzLGx7YobkOcqdRlM9KTN9MhPj4kGN//EKg2oaJ14NOaOQw
4J+n7Q3pCdR1wqMEjorr/22ZWcWLpfrF2qKPYS4bT9nqVdUdxmUn4giW4UbAy/DSNKv1UBvMbgCR
rbUdlgIaMGVNOj7mWL2XoA2+q7V1XLBbM0hgib4ZuND81W7BjiOq8SwHXQJpIcKqatvC9qdNWb9V
S5GJE6DRRxZVLQ1ODDDFx3YHTUy0y6tkYizfig/4nHRrItZKmlbJ1V3ejsggk6ThOYMbNy8QaH3j
iL6GIhABucpvLs2su1BN6kXmkNcFct/S96k2OJ+q7rvkt0qlA9zMlronHRcxvsguBOzMJX6LHgTG
dcbbA73DdmzYsqy7FyGOmZFa/gJacoJNeHzX+r8zogr0B14tyWjMJaSn3w7KqEFACa6zG6AjsB00
eiD4XKonUhARRWtVLSAhLv6h+j8tqWy85ZVrHQ3UOSSYlRj5REL5jWx8QcPc0TPCFY2iyoXWNTpM
xz6QYvpGVxkbTQPv6T2iB9PUxbPjxjD/xWODjPxwp3mW3UBW0qzNFTbPkZoO7/GV0JWVds8bPq9K
0eH+GQMmqPTrVq3GtC3v6z//mEVpb0FT1n481HaIztIo+FmzgM8cG55Y7cnowPev4jU+G/e/lmBn
ERKU3BqmzQDpQxH23tSI/fRI+/H4rM+TfgDaWrxY1cNMYnyqIPtkw4PHTP55b8oIWWfct+jLbwNJ
x0XZeJz+vj2urXAHARtLWvCvw9cjZ9WGSk5wndOFwTKud8W8VwsZ9smRvbmrOj1nUqIBt5BXkoVn
ghM3kieq1UhfwtYJ0Q6iN4wcYYBty7BzLqJMEKm2x7NVvYPh03B67I71scVWMTGXSV0L4Z/UNzpH
LYIvVHwzBcwsSp6yksPcvz36gTeJwAhQDsa12/oPEAaAmRXNBeTv+2HYVSX7E2GzI08WZvj1UC4V
NjGTSJGDNcu20pNQ+MokHBABT9nPEtLWRy1BYtaNsSIWjW/17mCh2Ph2pbV2wHSQYK7N6yXsQP4R
9xYPqm90ZMnS9ziPH5tpkA8aNYzO33DFnr6gEq1tEtwwyS90JR3fLHvzcaukcZ4h8xwtF3G7V8oy
t2jnV+sVE8GVO6i3xGppMJYrv7kkGhDcXG/+QVR+2QZ7DQjJ0dCh7xUpRH+i1cba7E4cqSl5MNJM
4n049LS7dNzccp2hhWX5aYNswdTO9k//pCmTrV3Iu9Q6d+WSkhXI+HjWJU20dlERb6n6G5hTRFmR
tUJN39QRWBwjdYTMvuKRTetr2QyuHKJjnKwJW3ds/bcZhGSWcJkk2NRece6aYgxG1w036wIQICiv
aKjds6dVOTJjOCrZBhI60qwej0+23TXzPHzeDL2zu7xKvk9VrENapiZJUftzX9HjmoYZetgQgyWS
iq42/xEcpi5InDtoa47oHSqZXap3jQx1MqMHqEORgHiX5JYOvl+lB0LSc0kSZHYah5kA0n/c8Lnf
42FUVmVBwlCsCwQoE5BYu1qsW460AuVxq+xAvIZMxlDPtdvR9F5Vqr19HYre1e2MtUCw5yohkl6s
C7AiXblfmW9IFQHXwNSr1UjUlBa2JtDFJJVnl2L/BZmyWl+uHx4xri3kLejbvau+x7oWC1lE21oc
iPOF/dHnr7WoCwlP/IpSohtv1/X/MSWLuI5CgdgZjNFP4mSIR/Qbv4S1iix2Vv8u1ohVYmc1rFOK
LQdES0h8acPID5KB9EaZAquJeeAY2T2HjNOIaryzWVJ2PjbGWf0jbtTQWlhrG4DfTpCFQFo3YRTL
/dij3RCiRQLrMvO8Z9vQYS1N/fbrnRfvS3XVwZi7p/5ZOqotlcjws0QTs5D1kztWRjqNdH5HODjh
zzD6jShddu8XNyOlo4KBREHoU9FYGrA5/AlhE3Vth+D8oYM3DaE0lfkml9v8rgVdsqpEki426M9L
5gPtd8if5C/Rorj4VFXtxKqGQVyenawkySgYVXhe7Avd/OE3RNRQwsbg1hPTh/h6+bXd0S8dhgMh
HQC2JIWNCJbfLq/PsTQjuUBBijaZfKX6QtS3sQ+h/Q3EuBKT5/14kh0S4TyARJvgEa9Po7LCaCNF
BYAzggKvY4/acB4f3S2a5urhyH//s+Jd6SqKU/Dht9/ukk9mwWF0vlk6TdbNIlC9/9QWINGssFKo
kYh0G5S06ltvfWHwHRMaATVTg6YpLFhLZBCRCVgvZxX8/rustlJmpA9+5xzI4k7WB4aq1xgAZ3cP
cLN7XX8WZMslS901ZxXw/V9Wm1cn0VYt6tsR7XyqyeiMopwxcZQs9ICoJiO34xvu/4fvsIFmDsQL
IRwr7v5McpMSQR8LJASi+kr7a+Y8JuEJLx9Dcf5op+UE9tjq1m7SN6NPwd/w2wO91USsp0/c4fyF
vCLT67sdCXVZ2avqV2IawWn726iUubhbZqAd6zl0QTiqWsqfy9ADD0PoJhx+FNNy0wkIaRACEVpv
8GCUHO71iaBDx53RZDJnhzMVTz70MYWAI1VAoPxDPk+/Ttv8xmL2DNg9Fnky1G0Tvl4yQDZHE8H9
s7yAVZkOcX3GzqfG5b9cScQszBUpA+93CmIhF8tpdS7bW5t5Xt+H7vYWoVb+TW4cBHiQaHt93sal
1LVB7uZ/vkhLgGl6IlQ0f1p19VpwR+MP9tfjLfAMblJFqpV9D798DtxMfDQKwvYRQk11RcF8tjkk
gB4wyAdXM87pbo1Bmjkp8lbC8GYoKe3PU9Qsr3Jl0uJW9chvSEhojMS13gga4TqSUYtPrWti3+du
rUZpFpl2zdj6MFzNlZk0a6MZRQiKO54BjAu3pc4r9EvkFclp7cxB4pNOXlH+J4JXPMSPvUJkeeXd
IOBLmIQ9Lm3aqDc4HTtkubFJwYsIwwIq0OZS6VFyANf4ILI2JZyXwrHhpOdG4BWPi5MvcC857WTP
RDLQK+zfS4iUtOtrLywPyrfk3yK/TPzuV2lsToLrrl7w4FvquNNfrOwf7xMxNiaOcKdsBX7N3m++
S9C9+U0wmyvrnjGLruRo3I7VwwvpcaN0Tu1w9DqpVldg97Yjpl10qWzUnU9nN+ca6TpzMIRIGnLl
XESMM9y5YY8XrveuyaX7/JAwy0qy+WznQxa9SY9vjV+ealfnZhOn3rrArtk8x3W/YzPTJdM2WJuI
4WNFEu9I/ZRbbM/k75QXIVAz3SNH53j76Xujg4tpiXLx0jf7iHKMFV5Z03+rupQ4IsjRp6TN3wTY
bDoXHdh2ra6Ym5D5roNeHSBu44XzDvuRvhAqxVTTt7blT28N/+pnFJrBAV/Rj9P573meoIEw+q46
4tpGZvnitjTueFC0DqgYeIBrCDbX15xaSK56q5rLvbVdPWaE0GkFklM5vvb5SccSCh9rkq4MBPEZ
7is7lRdKggTGglv1/VlxqfJlCxI1V9zkR/4ffzY1tk10hkXnLwrYa3VN2a7DM5O56MACyFqZG7ii
q1Ol1RA8hoRrHElXcfQIut/PoQ7wdSe7zI33Uob8/g8p+pojWxwVouqVqDpsBAVuxkS5Il0oHBXG
j3MO/4VrgTHnoRqWUZC8LuveeO37L0zmDCSx2Q7WntbDCtOVez8fnWoSsDpEc90df7wyJUe/l/X3
sIfOsXeWFjOGm79PMorMk/YBVF/XVwXH/7sRDvVW+OhOUOKzysAHD+H9TR5TFPY0nauawZP85Po4
+PwJ636DATRvAVC4Udl2QOcQmIQEQsmDvnhGeDaCcRpyZNhynrqt4xTrQzcD+WTQiY8r4VeaFHsX
KfJ1F5LZZXneIae5zpSMABIJDI1LuYyFOJyeUfGJfRRpAZfOoWKyX7B4JG+Q8gsz9YQ6Vd28hRa4
0MhllNGPmRc5wBxYb3v8/zfx6Zet4uT4wUXF8jRGWLOPupWIadOnOFlIX07qzfeHvKXLqXjqQEbP
kpysegFVVdJ6mb33buaFtsvDoy8rt6QwveEABPYSfutcPv21Jh1gVdi+6t5rShpgVlgKXCqCNsTL
ohf/MZ/noQ0/nY1qsgScei1RNJp7tCX2zQAqpHbDtyKjecXbIEcyEj0DYiMPbul+fU9UM3u7Wzow
QRH4YO9uWjYfmTVBg0u3nbLo+AJRWYOFrTkcloGwJIYIoRSs+und5l3+AxgfRrAzVll8FVjZuJ3y
0T5uBXvyxTt7E1KK1LWnr3peOws9NWcVKjJ2CDeISiEbTHORM7p+b8wyaXpaCDHarSTYzhptkymg
gcZoDBUYaHX9bWEyX9Hk216mylOba0kA57Ko5HPLGFq4syYSXdkFB2IAoLI/DJgq9smyTHbGw9PS
AWY0esO9t/Q0TtwrLdKXXJqUBpH1eT4Wp27W4w/+7o6TlmfhE52Gu5tBhvmKWq8uQ3biHzGMeAT5
0UhmX3kTXEDta+s3GLThXMBHJa9pClv4iTscSPiLB+n5CGJAknbI0pTxsLzd50fz823cbLSwcylZ
e1wkISceZ9F6V1FwhFvvEiyecoYBPvIK/xH6wQgDLpcr1WiGqBO4Zk+iBTidJ6hqrZ4Bgx06VifL
VEG5byfkuSzjHQX69nuY47OBtp9TmDrf7EyADovwdfdqM2KkdRE+g7yvaPfbi2israQZzOGpJGhZ
UsVOWTgPNfgPSW6aT7INwBYkuMLqlmVdniFr4vryIZQFgrlQuVPoVqPqN7m4ivC9trBHGQ+K/xeK
K+s1fW5SW/JywWMH5BF5IfmfWLU9z09zTN7IcjOM1l9mJ2crSPMNdts1TUQGVPqPXxtgmV+SiIi3
qEwTJg5vh8vII7A9QUFJNIlf01HjQcuJQU4+HDeR9rsSDe2/ApGixYrDic6F/LtpbFX+zstEUyz2
fG5hJw4xTnsj20gkgLQy/dofUI4f315LWmmGxjXtf/d2KLa0JoR5uBZmEXjN+8YlmttDDX6DMIkX
ATyx8550NLPOnMlDTUYxo6elZW2cqCxV9I7WYkBVkMZDWtC55Q9iSKZO13ghz/Zv5hGG6jTU5wC+
wpefQXmNev6cLUWtzMfVEOBefQOn3iaMO5d7glZRm8KBgEoNW3jucNP243zrriVuck4UmDnXsy73
SUun3P4neI81oEhvUKI6qAKBH0Bs9pBPFo6RfbGD8elcr/ikkUfHi4zmIDSkDu/88kMK1jt1E/oV
EjlAd9FFkTMz6Xsmj9RTKCMEsS2gMR2Vk/3JD97UkPE459XnAClnsryWQ8mNU1TFr55X6GPtlP3Q
oLNDNdlaODvzRIg5a/f14a1KDg29Dc3KgFW45l6TG/O9DPwJIZf4Kn84KtebXyWsdDi1dc/Ui+/E
cOp1MPREE+DRpPF7zGVQtbhQLmO6eH0aEiL5QMmP31HMSFgFr/xRvL31ClsKqy7+fgNjqePMA8ov
w+FrmCPyjsWUfUYlusAKgYoCMXer7v88cGDyi+X3f56nG8XeGoFFMEXefcBm4xlpv9qO7Jhk7mm/
vsJ5+anmWLV2/Dw4gg1tPp8asb7eSimKm2oLtavz70A+aJYf0w97afTDVfDEZoQl9j/F/ivFKB1p
Rn55nLTLK8vjNITUPXIdLhRsBYXaLUTPtnIJLWIfwmMes14fml41wT7wK06qa2HF45VrSedj9iQu
46Th/Vwxvibi0wMRZJ2ztO9XcSruTmPH4YQVbWKokpafmhI0+ZWBYgFLcdhyIEGp0tKy6SjlSQd1
pl7mh0iYfYTBb/6KYy8DUQA96BninvH9PBCJubJnPmZaisy8bVuTK0vTBQEqcL65lEKCsPQNuchG
bdvgZE/LwQOMEXigJ73lM68tWyWh3VpmLF5oIGZR4b7eBnWQY6lp8d+qQDhPSysZwj7xEAyhq16P
+KR4vADn/4wmKUegEh9kdPKo7+ZMfpEgfepkxGe+eqAfSeqYeYh/nvR2fcxCuoD0MO32zfleMSkN
KFDXoTEhZS18hNlJAIQ1pyxs4bO/B9IpMSa8QJim0t8y1ipfIJm2roGWL6LQu2W0e5mUiXA16YTV
PLyi8vgrBJH78JnJLZ2wSLvDny+jp6jVCEBJR+NIHJKhLyDL7+6UAcmC4Xg5mMaylim2EvnkYFFE
6v1KICGnEL2niAQ5Y1Z6tiyJWYF0u5IszAIfAeieZHeHJUBpMByHjMQSYRN9H8q8bfKqJ0BqqjxQ
XgiCm3jwGGh3V33aIuPRyVa7OSHaPIMdgE6K9NowrMtTUuipEnghcsvHuLmd1aMVi1ohdwr93IH0
foq7+uMvVgUzMIWDoRjrUIwAqoi+M54K5aE/TNkr6gEYVvXuqCFe61YXf1xtWAYI1ZV8n8RWzDrD
2Drz4E74Io+He04yiaehK1yB8muwkYJenOPdQ2y9/KGYj/N+eYZdBUX+9E8Wp6Hj0kfE8jasTCGI
3AP3xoLiL25vCsokX2SANjq/J4hadkTWe9NchRU2VAR1sSUQmScFzfDghhbu+BJAdDfeGBMtfaHC
SPzKFLwf/7NZYEnPEUTGQBRfyYDA32H0v812g7G/Kc549FI9oPuMVDWJPGMEdPli3FDYaM39bxZw
8MhuRREdL/ZPVjg7PUPZ8azSnXOX9q/yMqDNvS3EQTdgKQHMrG1b9pf5yENvDytyCcIy0nDMrORO
sSAGODed9jJVrlutlRfm0btK9gr9suX0q/25Q+b55PDU3kEt09uI2/MO+39R1qdRJLCz5Iw0iFKJ
F3TqniNammwKWyskvDYqjz0ztSGLn2aimm03ZJS8A7a2OHgcQWW9uTjuvDd6XFx2nbZEHhql1ADg
oRSriSwe+SnxvGbcQogtbUH/hBOzRkqq6dJUyex9BiI8kySo7opaAlBiSsTd/MNLBVOE2XlGx4L3
HJwu6aGWCeaSg0QCGN0eo1D+Z14F3QphxVNcEmrIBq9RbyezI9CnDxdFnhmA6++txR1tARCnC5dR
25qHnJ984jsZhQwDWyFAaI3DdrK7YU/URiS6tsedOG5PdX3lh0LWcplr7pGHpopxrweYTXxdh3si
odjACvLSnJH3kzup7lXh5RsB9GH6VVjhA+gfeRDSLGxiKhkhK477NqTF0M6vIB1UdseoMDfOWnCQ
Npjs+i9bHEwWH4n6s6m4FZkp1hmerw29pceAFl/F4r8BEs/JrQ8PDFihAuIciLTpk6Z90iLzSjPK
Tg8wnByEdhQhQteGXVHircGule+O1AFudvDSpKzZdgzmskUSFRsDfJs4+GImqcuDpjq8A5asm45b
Q8L0eQny572RtLteEmrQsDJOBVhVmAseNxkP0k60ZyxMQ0RsahFNGFu2/m0mk1GySnaW4r0rCSG9
lcGrRVJ7QtDu11pnX4sf3gsCa2bhekb5oQGG+padEfKt2Axx/RPeBdR8DGDDBnn0MUOejoByPl5v
JkAUHqxCGKq9VnQMEWL2ky+vJgRgOHT9CAiqnXfQlo3fkzSnN3nmBkZzd5AwLmuiRx5UZqGoMOwU
x8h18pvopwqDU4v2gGJaHRvRdZZlMQ/aZigmYpdbFDv1Mx+EUEvfwrLCfrGCXB2b4Ddepo/YAoGW
n0mri33Ydcu5sxj3ze3WVogDzyHwWthjFJ8OQuf/YDumKEFG9gx8SUijMb4outcSwqSuCY17KwRm
CDMeQs5HyGBvCdy4fzd+bXaTIOqudUXhfFqF7yTVqKMGrEY+7rENKsPO5S6FO1vwHjKMSlND0DoK
WlTGLbzvUDUbe+4Pdcvsx4ZR4XVENq1E5YX2qkbXOWDhdcXoO/vKDmWjFtOh88Ms6k8ZuWRLNgjt
KSR3j68T14w7jSYwSAt7n3P41dLmqoVZmIW/uqO0Zim6MlsCo+OJr5AyM4F8uRTrX+IpRizcLrc8
mzYpunbFQxXHBRAoOyUcRq3BLQnFPf4SlevMq54MmeVvfxVW+sSVhm1+A47vK7v9oZFt6rfdBWRb
zA8q12OgV7kLGuj2LFz4Rjg4kV75v3tawsDwsLJolpF9yrbAGdG/8E+qwx3DwQQ1g57EO1Yjveud
GHrypi+qqzTZzbYJ0gIOUZYSvx9bLVL2Ub1dP9PSEkdbyhQY2ufF/eLd81iOaHMwHSyIlhjnOfbx
HwEifhA0u4mnriTrCUJ4uIQ/u40U+tI6HHVew1UxLfTO7vzijoObLz0ogvXdZxccjt/67+wEKBTR
E7aiVulXrdP6x3xBaqI5rfpsAAorn7UwNJgqZhCH18iLaSuihSqltSTq1rFDqaEwfZ8J5LtOB0JU
60xjzjAkAXt0FVOYuPAe5sEFldVZb0ciln0ZVy0WAnkz3mknUYY4LYitPDnNtZioClDLMTgPOzSn
JoIfxaVBe7KPyWT9CI/VllRxhiodRJDIeqUklytMOuB879yZvcuBNJbALn8hwSHEferXyZxDUiDO
ATuKG9C3JVxuw3cSDPOhtBpg7QKVB9eRoIWd/LIexNbQuxkhDn4L2LbWumMka4kr86HsKEnXpj+L
LUp74qN7aWmvZLgVO6/sjee+iknvUGY/cV2CR6lwttdZZlP4PF2krnxn0rhGCQwBXlT2adX9MgRB
kaj2pUJj2sA5Cl0jqsyAm5oUfkBL0FgSfV5g/4PkM2DLigdJeyJuyPDiXfFGBOZ8tKKxx3iGxBFK
1h/UpDjnh3RCv+yHQo6XAc3ZhY1+arw4+Q/YP7KRJ4yva0AgJKvOdFaPmgoiSWMGNvsHn7d8ukYe
ghYe48YY6x9wW4MPl9sweE0i9ykomHOF0YCuSWyfRpxTCPbj+f2VIFFRmn7fnmj7L9EDeS54yzk1
2kB1K52GkrwQdIbEZ1UqqWE5uVfDyWOR1OM3NQH0uXL5WzR4VgdIYmtqYzI52CfO7n5Tj9KaFyon
1jxh8uQw5kONHONSsWLpxMevqxPTQwNGvXnzmlLEr8Kfw74ayIjEWoCeKcr2GhMENXUIC2LdisGX
HvyRBl76vXueFo7p62uJA0YYStpeMxuzOdmbh299tUmf8b8i/wLNgAof2WcG1Pw5aqX8QBWI4f1A
xxsAW7gkVRGSHOkcS8zgD7TEXvHBesSkladkm1+nmL9GhPC5iAlRSWXuG46LMQPs9fAJcK8UJWeX
a6Ry4kkGcvY3veJ8pjBs+fVl4UVzbnPnOcAy8TFLdOfx4HdSP/YAVPbXxjlxjppwbZJcw8d3rxR9
ynG7Sfk89SMMSC/qsI6QcdIPZLj0OHNqw4b1h2MVG5xkhMDGcbLfki+gOK0YgkpYgRMsOM7dYlyJ
FpH4RTWgVefU9/nuchZIGGCvUo+fKlEH6zv4/SwlmWUqVE2NdKXiLI0IJ5v+LFXr49/V/JKq6kLA
iyxQjxRUhZTUopWZljnsPCOVGpNsyx0iWm0kEhbS69TUDFdA/BJ5OwE8GLsdODcsTy1rNs6odcRH
n8zEPxFupv96c9aOKP4ZrxAalU/d0zBid0YnKOSp61P4xmsPzymXiIlFqNUyerKQRmV/QZ1CX2ut
efSuNN21uhgGXLt0+udEsVsUwmR/yKNi3OujwO7ptU5V4Z1L1/99Mf4+Wq4Q+328Mq44hVDad/qV
+kagrIvw8wMxkiio8WeIeDIbrN3HARpRb9WQxeDujQldj8FDgjpJktUVBc3E3Bj6jjFQ3jY+mwcQ
W/Bx2SMnq1RdTNsh9uIwfyLdIBGkb5bL+HYmmQc+u2GpcfH02Ur9WZZCRzy1vzIASOzK9kUkF8ua
tRZ5W8ij6Pu2Pv9T/U4z3sQiSsrTc4CwJz481e7BT7AMfKK/z60SU5XfE5I7MIZqZMFOqBAwFpG5
63g55ARtiBXotCYVnZyqP2QjuwBtECjH+oixDqueCYwQ8ifVXHOjuIUNBAuR5sPQIRery8XBJSFm
mHxv1F5r0qwOXP/WXaxoZkWT/9aoB5x+Iw9FwvyvX7TouFhVLmxkgWZ9+HWlHUez/nCjQU/IpGAx
rLcPHl9B0p09wGuhpJ25DBqNam2n/SNJXLYo2cLdSnsfCC8+yLIN0vu/7weEFlzVA+KilG/xn4Rl
dFGYOang0OJeobWtw54kxZ9bIvcaVibYYmtMm1YEAK+kQWIGx58SauT/zlcGCeFTu6wsxdgdF72k
mooIDGm7gG+4MZYjpWd1mxi2iKAbo2vd+u1wdyifOSka1jZX/Hxf6FE52vx0Vc17LSs1ArCossta
l8EuU3JR57uqJKG6r86DYd7ZLqGuhKmgRC1awaogNgS6G+sjEw/o0FXjct0p3yKPFq18T6/LXl8l
MMQE4g55X3OuYgtBjYNfUvgjJ9t6jYd5MX92MVaz2MBZleUmMo/w4GtiupbKqew0mYx7zZY7bE8A
1uP/hG+15NL0tA7dddIm/IacTefRkKFuxUsVXGmREIWQWfR3EWxIBeBf0hIc1N0TNvzMtxFtkKpT
tGQEXZ4Z95P6CM2pzCIjcpTON5T1PYEOO2x6o+/F9FI87P9qZaDp2Ugp/QT8whXhIsKFmReGmjZC
gTRizkPH2UbQ6i8J0AF6amQNnF3Fbd8MlNfsb73LO1gbAuElepgFP7FsaQ61kN1hImnq/XKl9C5J
mUEAKHOrCx4DK41pFArBxJcq4nNzM8TAIZME0XiZh5k35K/ko5WCzql5OSJI7EQmuzXq9PEWkc3w
idSL+AAWLZqMhaST/B+/W7QyrX2v3LYEBRoy8jWUeTAGw2c77z551V4usePbOzTGuz3tzXNKbU4S
IlP6MJ0np3Y+Jy1jijOT92lMD9908v8tx8wB8WfxR2uBU/b364d3/mjNvEFmyjHNihB9VDMyLNLy
+0jmGO8OBcWXtXJLDxcuSAZnQDer3ylZGtg+u0FbO+WmCL6ccdlC2eFKnO9GZg4br1lCJqSxIYLD
OdDapG1NUwSXmVvpdJJytgJionEBabYCYI0la1EMeg5Qjkt4y4Gp7F3QYZ1PtNUvspy63LRZOmOR
lHMf7KSUZRHOD1QzHEpAamXG74ZBJ+CzuzMuXKF8eahEA1wSkWKvMo3v88fa3ve39dFiOcdJJIN/
7gBcMHsn26lLx/nwg64bibOTJZMDcFZgJbCRAYtsfNxSuPz571SFUZ2JhEVtlJ8hAk7zGz/1JdQ1
J3/yNEY/LF4uRCyNgf3fPFjQp7HLpfwCiMOxKETpi8H5tJgkQiPCn32XYtaMyaB3TYYGR7li0C6i
ZJ15pCzUcwDhUsL19RQ0McMlqOUHeiWCYtyVBOW2Z2qJPIS/TyVbmRql6w7BkD3qAkrNhC9f67M+
dG82LkmNOXQewtTMnbx7ZdPnzKxNrJaJMFCRCdF6tMAbNjC6bYST/aE36Qmgj8kuYg/K0obeVr9B
CLyFPIfVXW+tiDNC5OlIUiS/iJKxfRHrg3QCKxnTSnNDoXA1ESvPPY2Uua7kaMxSCG+S4qmrLIYi
vg78sZwja0gyxw33rPWfIUcqhA4eypVK3Jsd6ecakPlE8x1JBfyCvB7VgGMLofM6cKGknVY+9Orm
ZocwdmFOB8RAyv6QnwZxiP1S31KPIlKievi3qGsyoYwnCN2SQtFTqlmqZPvXAMnQvTEJNxdSrxVc
sBhFPUFpJL05voNCqb1CE9Zz84/ncvHgaOHaPWzpBsI3Q0LF7WhElH8ff5znlyvQVQRLTvz5t16m
aSK9hfFGdeyPeBKFr4EEcMUmWbvdnPbq7T2MAlXpY/ykUvvtx+Z8QiyjJpDV+rZoFauyMrBT6+n6
wpQQ1oj1iRR3cC5u6q12ijq3mwzOY4frGkSOvlP+wALtzqjSR/ysmPp5V31//XPqhTOKD5w5vEgy
hOMH9dv3Z8M2fZMfXx1qY1ltVTjGh7X2pIBNzLfrUSw56wRQPxbeF3ATzAFXnkEIe30qLpdk9NdL
98oD6EISpa0DpKwW6opLNg6k1H1StBXd4e8QTcd+GBLKj7mqAEWxllxLCoUvBvVjlBpE/6dvmps+
mSz9aEYPECXa/b4xFjJISxyvy+gO8O/Uv9d5EyBJAHfCjXiPWdG04YKy+q2jLwIjKu3LcB6f5M5d
hbNPdF+kqLWu8+5m1Cpd0B0vKyj0hCjAzFS21pMPba360WKVFnct/BUNwGLP4ozmyvT9GGT5qm7k
tdeL9pSIS76fU/f7E6nHIH23lRYU//huSHTKH8VYu/2ZgTI+8UuXcWRMd6HTiPo1d/LOZ2PMcAIh
uFBxlDz89jVgDBTrQIyY7m5d+bpRMzwdQ6t3o+wIXyRNOQBcq6RuJVAkQHKOBniSZ1aEHf5iesCr
Z8vewFBR3VAsNDQfqP+x6eG5igunwLufX7WK2/BhusjJ5v8N6jTyEYA89/6TUjU2BIljQsGuIF/K
8VjIYqgPOFQMTdYyt5IEb7nWCf4296lQfWld9SiSUUU6uAYqvKlSCvenpIle6MqvlGM2YTDfzTGY
/XwU/vMHpnNPfE4YEnCkh9DQ5wbjCaKJMfdZkcZDGD5IrwA0Fb4MNfesHvvc9+8yS6ay0XlCvWU1
tLCSqQv+9fuW7X7WBLCZqzx1Sep/3CAt3r+HjeB6/e4L2BtH126A1aRQWxa6ueVTGNXWKRJSKQIv
yzuk9gNsjIOgChcfCOjPqLI7Aq8CEssm/eIu5vDbUdMMdXsmM1/ZcEs4/xIAliStsl6CJ3vYaF6o
vgoBWiEU5j7rp8/B4i7RLToMMqRMwUTsNo6n3zU4cfblGEAsS5hwgFSSpZy2RK4z1z91JvI4l0nh
VptqQ7N8Q96ofP59zS68hmcQ/ZHkrWtdFmHo2CIXOBFDPj3fb0V8pbmAWzq5Q1OnKKg5XqEFilCB
saeoY6xTaTro2SFnMj+zEzlLU1YlVSDaAxGmHjfz2iZCe2pNvMMMlTf23LIhX/W50RmG2jSHj3Uk
HmY/cM0CqAotJk6vRK52LrQeFKOvoTAdIFzGR1nlR7cJ4c8/PL6iGnT6tyjq6+Wmyx92xN1HS7I3
4iIU613QaV9unBrnzH6CbGxvunEUv3cNVM6LHhD9/Z/9QPrLtF97tdBpWKBTzr5nEItAklzGga9D
BAeVNJZvcQ3GNHmfgzt59+kNgKWOQlUhqkstVNXvWRDFRI6eZZhNYz00VCpev4d5YgoiiiOtaabs
i7CX1GM9HBupFWjcJ/QZN7VZCj6qjj5+kMUIuuM9BOYuruGie61/yj4fMD+xKQ+zNMYSTBO+LUEH
PPW21kLpBkmnq9otAPB5+rtVzVc0W17NJ5jgGvJ7zyWCcw9yEIB2TPqlTK+buqQhstKsdj0WRBGa
Us9djXWJRfILNsLW2cz9Ua4IcKTvnQVmf6bT4wJBj82N/cSlv+n7sc2idYevaeXuhzLX+mgW61g8
kSE6gY2EV2txHGxcexigV+h5cPGpNpEWqjPL5QFDSmCyA5msgygxPOEQX3gVCRtjnEaDtL/lFUcM
JpiaBqGRckl7fC5iVQP8x+ROji8bVbyt4C1HHGqu/icDuDTZ6t8qBWBclTyA+P52rBLrIeknJGLK
ctBvjEInbadQH0undJqaDlRwTc6ffxdugFJOX2v+X6/tHc5u6BewAE3l9GiMlkw+bVs/ag42nhLL
XJUzI9r8QxDz1F3yB4qIVct7WAHExBPgorJ9JpBBxmQUiwpA/fTpzrBBlGjHEi41AW/OV2M65Ji3
qL3ArKYlSmhDt2/3ZY8II+7vgxqUEBuxfhJIgW+mDFaZ39XnVuCWytKRbQZ+b2Fo4c/viZMU82qc
IVqyZVhroUdEZJTpDdweeJcfWAOxCTRrTS3gpYCHIyRGZaR8ikHaMGEppJ36PiXF2Up6xUVyVHwi
gIFlm9yTt/37Z759G2bo3nWRqvIq7ijfybxYjoL3wSYS0XIceSEgbo+saYnEB4+Sf+iV8t4I6slU
4uf62VhqJ90qqGZyk0LjSF8IN57icaJKOkrhvUW/NGih9DSySWG1wzMmiDycrajlfSrP/TJhu0zl
gZFIiXM7iaUyEoJC4olrqDSdPYnmKr8ziXmGxk5KVlegGrIBpmbprbUbhQ4uJWPUoZ+wAQ4jkUzX
qd8qdXYYUk9FeHeThLSLqNxQcJ9bJn4WWHTRu0+vGlrhakk48Xz4S/29nJOVfa4SDgTzG//YqbpC
qyj+YnTtPI0L+03LRyCCzuzqZsS6edauWowuUn9sK1M6ALgI+oBAIVznmCzxyI8zZHqBWwvrRJ9U
+0YId4B8e+aPGPVaB4BYBinRVYLF9o15zWzt6jVDl5q48fJoF3VYtYBwQXL6SE1F9xbsPKHpdP5T
wRkmM/ES8vGTz6DWQebKDho7LQi59LZ/W8jmCTSDyWKKWpWqy/9TJzh404J1M38FC0CyQCbxZYvR
B8GiJ8LaXPYGt9nqrkYH5YVdV6ltHY/njnCXiWE7ykg+QSLVeuJ1fVI+HmnUO0gFniVTyONxZdxq
tQsHe+EzZRNgtR1/PLGXwDe5iW6YRzxrpydlIpE3vyu1nAGk2LZFQgJVQJjuaa7hWItqZ+cJ9kUE
Zz53ld4wMIi3B1E9BfpdvhExcZbkS7DBM131wg3G+31yDLVji+1AtpxFyS6j5RBH0ITS1+j6WlOA
rL7EdUieLWeG3wqrAPEQEDPO3AjfNKeqIFFLmmspKAs7q4qfU4018GJKcKsDbFRxj0199rtFPo7n
6+Kn0g2QcxqNrOV6MatTWX9fc0cbSvG3T13ntLXPBLKhoJ4R0aB0lWBec309n4nYi6DE1dpCl1G1
mboinRrG5ss8xnRyILmmsDw/4mdDmRpa0FiEA7Wp2I4E/Z3W/W/IHAwwEu2+AFkYqG/i9UvGFkt7
pswbOWzLs8BVAEw5kKIUFPneBjmwaaJubJTiaQHyVTpG2L7SCwsq/dEkh8zUxLYR7nUdmzuPRSeQ
82D5TMBUBJrZ7/e8xMVvLBq2HN14UcczPoWXR038dJgcRZY8Ufo2j0v7U50XCQxh2s3NJXxJacCY
7JyGUxNJAlGr5r24b1yZfjih5AwU52diG1rNn37CdRL8C84JbB91AfsHo00J8EjP5834v/6H0Z2/
m9Jh5oyi7iiKOCal5mzHyZTQUiWoRYhEMLxgyMAaP3bnB2wDe/urDY+159wQ+OY7VnuIxHGhmJ2B
7GPxdcdBKcYzOf/rfJ3x+uBwpfpWmsQ2V15/CWpf/wSFz5f800dapCItZ6v4HuXlctUftIv6vn/7
nThPldhrARkhj/XG02lX/B+fE18zDuiMH3T+rDzHci4eOCHHK4i9GoussD48wPqMUPsyJ6oZcDVY
aZUPq54E5lh8yfd8qaU61Om2C3NRFtuZx3SY1re2ioTBUX0bdt/5jDFCFJI9I/BXFd1xkzevZlLN
u8rLD2WQFq9MPH01Eyl/SuUk8nslwGJlrLytt3ib9HolPmOWxDKLm8XVt/qhPGIwbY2OvvgUmJyv
JtCmsOFaDhzz6HO7vpj/l4cBsK/6MaT9AoUCpvjgx99+o8V8L/yxghXicLT/aXZJPdOuq0BiZCJ5
1mbek9T6Xa4AgKsVTPEDZTxsO+oN0QRUVdLI5KeYIChCxYuPlcz/OpLp3bmkYQjK8h7kFTn5Jg6j
xtlSIsQrIBQ5YzZ1Vtu/jAdY5mzWlVfHUH6/4rjQozfd9Txn3ACG/C/OC31aswiC4k5wuObiJYPC
FuwYRwiwR07uAB0VQ0R8QTgh/HS0QDFpwJqTNqcSl9WPrGMXDBYWl87A202k4g1EQXn5zZ3FUzhJ
BO2/74mQd98x/Jsqw5ai2YNYglnLzJyd2mx6WCxYZcBmRldwI93O9wl+7U+11RszaH6WBxCQWZFg
WtlRORM3bfY9Q2zPYPWpI62m5rngsZCpjo9CywWYupFSPSOMFPRGNYeijki8n7oPoQeZffx2U3QA
eFE4xiXE2Ash6/lKQQ6hQdBxqnaHvNa1RfnyQHcUXEYQH2pp6MKzEQ3yVWJNShBtckM6xBbl3p2c
D5gUS24fCbVf2+YWY41Fb2Z9tuu902fuFI1XRyGXfFYn+6Ffqa2iCgRVzJBhynF2RJdmaukneNF0
ziGF0Wqhs8ANz5q/vJ8SuUM/iGCYR5CKJQZS+K4M+kf+Nn3tKxucfTjiqXbDwrwlhQ+5XO69wAA7
84zxh0QQuBf/JWEcbWwjPSRCpRnDzq009yyGT55qv+bslwwocFxFjhFsbh1u+H2IA1pdBFWjjmPo
jO0yIK8sZWy1iw4AWTVmwMQhlGCN2tHr0HNW3Ke+u2uT9yIWX8+KJFgPnJklcxYQLWpbyxIhpLL4
n7wd6p7MCAPF6ALvZTJjDcaArUnYGwFRBtjhZRfvquznfwy7HlbQhxcwYHvPDh23I7m86JdBVNqq
PCKrOLWr816JVR07bdFqtK+DTpKYeq5VFwB+wgUrZDfot0Jq5GLmXPnLeJ/lUwgnnlzxBq6pfVTN
j70vEtyD3sRn0a+2wrnDh9zZDZuy/JKbFVoGSMA26AOfu/9wLJ7XAToVGPElwSbZ6US6dfnCrmZy
18z4PiPNMWWPFLFQnE8ERYemYAf+/e4hx3kSexZ8MvZz1cy37tFrSzukf+DLtcSSxcs7zd1vZxbp
KxXMToMuy0iMLAEwAMFB+/TCQZ+ut9ilwjzutGJ+Yi8JnH7OLagnLADHNe+MRiSge4nVLyHrxapM
sPrwDejZAEN3ZZvVGC5mAZCDqNm9JyVteGlYp1uRm0DueAkIHXAk3bdDum7YZ+J8LfvAOuVzQKZn
wO1c2u1SAsYMFnJ2ij5b4yX4U5KD2tOwd3TBSSD+zYF84cTU2tfFTeIskJw8f9a2PemZO2PeYlFq
ZXcFoFX6TRhVlwU9DHRuAwKwCKZ16GYavZpsfdN8L2+b2Ld5xGk6jSeYrqg+4yjl//FB8PSy/5mR
TGUb15WYokBwZRHX5h6kem94I+u5LKuBbkLYhnfX5EskrRYaw1FEigJivUBW703rJAASJ+ah0enl
M1+uqFjw8/HkgEAg5CENVMGLpWXvaa0vVOYzXjtSFLENteZ6k3U3I+5uOXUaQpTXwl9c63ucHIMm
KcmLEHgO32Q7AXJg792/OYkr63b6SqoHmod9hQzpS07db+guatcUhfEWRIfBMRAsu28RpJosnf8v
uz7FtvisVFJuBmoqRN4RTdVM9UFb6AMYJcjpzDfAO89IfJM+DwpydrmAD5Zlwg8KmW23FMMP0rlE
KW29AhjODe4Vzpjzoku1+KyteVJ+G8btrCNLCiR96PbQ7NU41bZxcc4pyR9KPD7PFitjQWBwORHv
EZZatMTR3yYUxsZfKAkYF4UZGTxbl5PvJR6B5W35CSCZb3pa4eas1tmleI0s01Sm8J6afiRRjSbw
FOs3nF76I9AZmD0vmL5As4DJoDNXO6WPL5NH+avi1r5zL911XJnYb2RDZgwrDqcquddGyz7FDJvT
cvtjfMELkhlujWqByFbbcjlXwQJ6RVRh/R3J9AY7DZUa1d2uIfE3eQ4wVg9DD0O7RyXPP9ufhK/R
qmwJ3oMmBqO5gXf1TLXYwNcqc2eiMrfuM5KCAbfes6DxL+kCdo4lsXIYwoDwIcukGDg2MOe7y7pW
+r21UcYkUNCvr0pdD6Bz544tP5t+ZamQBChKfp21pgxuZHubWM9OcC905F8f2+eoPdVQVremXv99
PuJTQihanS7KQLu39bDf2wU9sgFRaIv7D2wNbbu6nhpbuTXEUVxPio4/BxImGteSVOno2g0Gt3OR
3bsF1uZu83GdlBOBl3aBXH8Hl2KxacswnB3Roe0OoyKqZjIMh28P76rPtPkfXLK0dO+xmwcKPwoA
Ss3zY1BFRBrO/yG+8x/SAxexJnC/OrjOItBckcUFlrN2gm/lIQLM6r8pYTrDpkTGv2fC0UvccJAc
fRYLhr7q+Ska2xjSTg4OtgLOlvJzEeXp2YqzEFJsGROdAjmhw4/KwwhK3e9pgXhHQAmuZqF61IjO
TXcQU9wDhpQLkRqzVFaYZB6GJZwuQHBFPgyer93tkyrt401+Wt/dM2EDbD7NEtHAE5PZkKYDjbBQ
BVb/LtkjSfzkXPvseWTLhAuDTJoiK/+hCThL4WY6uhQI+OraEqpNY0zgzKy3efqUkOTkzQp6R+Zn
hWhgMrOn/2PB14/7jCGwPJlD6d/Hp9FMpNSxs9aeHWrPJ3hSeo/9sUnowt7Qr0ZBHmBNfsvkEKHP
n4gRnD5OBrQcYWg4ZL29p7Qj3VwF0faWdVLx/CVANQRYGv9k39isHCf/zCweegQjTvLQOSMbuGPX
OnUAGQotW/3up/uDl82+zktzVMK9iYlSlq4oGDqT3aadbRshTBpOTL9qxvq330P0NJ4hyEX0Xcio
VoIPQ2DqGNQG+k1RyTnBf/rHGhTjwHc9hMiaNgsNBqBbhlsKIzSw+xO/HMunlsr4x0BfwIEkrSGP
93TnaUcFEp2fihlao4pNX8zTh3i9TOknYWrJZS8szI2z89QBvyVUfPayJA9qhUBv+kxAIi3mZhxQ
OlJTxr34DQrDbeJ56AMpsjjz10GJzfaMGYAMkyjGbJ3XA6S12AFZuaQWod+jRcecE1VRfYHAkyUh
DVEMnFvMJQO+EEfs6NJ6cRrcVBFn7e3WDv4fuoXZ7rebyu4qB3AyLoTTlQ1vBqNTMEzqdy4Y4bkN
V792cMQg28+7WpEj81/YZc0higYyChjafhgFqxSogCXEzfveKYzLaiVkGoflIO5R9HlsjmNqeYYf
wAWdU8KxCEV2M/AjhSuMRUSVuS7kxb1VoXhGUMfsVnWUJVjzRmPSPL+rwoTYNkNTSN7ZzF5r05Fp
EpgXsp8odQTi7Mt0keJr6huMujbbgTtpA2CBVXFLfYr3rRT/32A1c1HzXMxFddhQ9ldPhzaFUZ59
iXYMg9dozdY7YGg7qtwMOQ4cT1JshOzU3IUgB8T/mfXCWUSY2d5kZoenhLKiiKfBaCVdiR6vNaoO
1XHYcZt28LmMkF64GUQsLLn0dEDsi1i19tzd7Lrlk8994HwoCb2SSbjJTHTF5OM4kKtRlZ44RM3A
8dT2LP6DtS98nyik2pC7JplNWomT/ek3+4k5UVQ55qU/2yFKpNPHGd/A8WtIVLMCzwGsZWbYZm0G
zvBeWM5IgsUcZnsOc9iWwTfX78dV4IiXSOUOe3k8wXl//mpqH4KIjV1pPGespvumSOAD0WoM4L08
N2ebVTm2ONg7CjfJSoVIKDsLtoxF/+ySI8OHtiyK2Ovspei5n0KEQQE4KmiX+hAhYx33vpWzN3C5
T0777g91vVxJmlyLtUZLJje1BxUOAc+mVzD5zJr+r13rkw9SG1yBk3NqVQIXl/4Fv+hLeSDw2s0O
BHSrHRvgYAaSDJS/sgjYTIq046ReJ6Vv0rg7h8yctLB51QlnFRv/Os0Jiv299CxnsXMG0q1MOJVx
vflgKz2mN/8Z6JbI6DLwvIk6QDIPQFBugXgf5otw0YKej26yJ0NFmn5j7R5pLT6+J3pQPEZK3qds
M/URP6FnhnQZ/8BYDcnlQj9O62c9R6QMUwF3juBzRCKLzHoweEszpzrdCg38USy9IG5WDwT2LD4d
xV2pLpUqQWxUXAU2bE8ZcSkCHMjeG51vbSXPKcPs1Kt6DqAhXKcUVfDE4736lDJz/GbsoY2nPM7y
Uy7oPOze3j/6GwSE87DqzlMxGBLQjJsHYOgW32oLt8yE6fWA0yp030v2USyd0zkl224EU4fezICV
xgrx6XuNJ4EyPgNz9KoLxURlxzTFLFZ45pcXlbiLzws8Lux0xNWXK8TjhUVx9yAEJQ47zBZ5iBTw
LyM56jVKJPcyaEGc0D9U1B8WGFS3j3TF9rscmw+N0NkWv48Ae80Lq8EAz6bQ3RSS9YFmBggdyGFL
AT85LUd0JNuwsKxpSeUy928n7E/utH/b4/zyl8S6prENV7Qx8MKA0jXh6dMkN6nPcLR8C6okWPio
JDOyR5tDzEJTIqMXu9dC3NzL+HA0eM5NLW5ENZxa2jsmYakGGFrDOvzDgmzHe4ctJYcgacLCnL9g
hehMLk6imK/dgDyx5R5cUC2B2e2JiGyXwDaEUidGLMhCZ2SJwJEAlMPyrkwKv/3WqOX4siIqfnti
gQ29PtOL5/K58tzGmL5K3xlQ+VZcU1jqn6zcAIgAyLCqG87k7xk5aEQ8xj4Sr8/Ka/QhBfOzd75V
qpK3egdej1Z98NbtgyRdchgTo2QYodaPMJqkOtfuCVxqk5GWOcmZ+lWblOk/x8UDID7E9IC0hasi
MimJ748LMhu1YGKsqcM2AP8lFMfttnCK3l/nLwdBkXjgIDR4AETdHUAyr9FIDuZVYZ5BDSEchE4+
NQchyxGdpE6RgSOBgjXRbNlXbWfFRMGQc9czMFIEBd+SlwjxInJq3PyJsGXAqV7ZMsYSy7ERzMsg
cvBXt+v91TLCjF+7C7NNxuDu8tVak54+0RKUSxRoZT4IZ4POIqFKJO2mSjaxBLw/qAUA+XubTwnS
dHIz7DXXwD/6zVW4QlYl+04UzulKfYBeA6Hc90lERpoAlWjLxYrQ90mx1JtbrEwOPCb3GMuxPtxq
mA0hXlKotvR9BrSsTdDnht/Kkuc6yL8ai23ugNolJjLjoN3BLliNiDBvsBYHL1fQHPgD61rN5yiK
6z5WE/dCZfYn6BXQUqZeONfijn+LUAcA9dRSHkmYrpdd+EY6qP3EoHqD0fj0Vl66wyniPrnSJii3
DacORsc7VrRt/mOQTNBrkrqbFTBz5uEhIXrCA4PXujy1uVbAiPgYmofK459Lvx+rAaeKbNRVdiUb
FYtWyAwZm4RFI2Mnu8amXcPIamb2RkEN5fBsMONHbXIyvxNhVlwh5IMAJrKN21pk0MNtWaxdSRX7
oK5gSilnv0/iCiWKV0b7VmO0UmYf/zzM7Osx8iRM4livk/TJ6HigpkELQR+lbPk+O/uQGIXJZhSV
427xIWqK6Bs0d5YRXZt4VydMoMbOu6W07QX5eqcFX7qk6DXhACstKtgfx5bJAYhkjZIdWWjOyCI1
OS17EWLwpHE2W7WJH1AZ5bPvvwcXQ+r/eEd9nh+NjQKgsvhcm7B4PsdLR1HwzzVCSANZoh4uo3gT
urdbaUNyAxPVwwrTRDHzgva5f+gS2wFLdndoc/m8VJYorON5LRXm2UZ9uqxZNAfD3rPpFRcRcXlj
8sl/py6WYhgUP2dv8MfOmqgM9Lo1O+TcrzQs9VFMBIobrhHVjwoFavHO4f6CjgoxwLnvN/4owp7S
HKmEc8LaBuYxt5g74hoisQ+M+bwx62XxOaeJeaVB9TbGvQc/nYXK9BsxX/K+33E8FeVw/1kN9jeG
CkZqArsyc/XXPG7r3VkcAPRiZ+v4hTtyVE7u6mCATNaX3lQaKvp+HYutgd2167YX0asX0jIuOvsW
InyQH9LWxix+gIX1y2jObZxvdKekVSYUJJa/m7AL3kMhbJNNQ/blgGghBThfQ9jkWkd1Kihh1QDP
s1tj/SmqC1rE2FIIoFcizH/JBAqNwQYcExw2zAT8Ra7qUWYlnejOqJwWmsYAjMrXsZWnAvHKtxPO
fCWpHMQy242uzk0Ut3y05c0R9oXPrnM8ZR+4jg+0mAcTn4zxyTi6Ulk+NCgwlYfzfRIcgRLlBDYY
BGJC4H68tM/yP94jPWqnMNg53TD9k59bVJ0hbDTogSJd1IhpTAGTjqKPEsysW+zSOB8GnUVj837E
YWaZZmd1zootxzBIB/QQzzb6C9otoJA0A9F21/NNlRxQorscwiVt2ahZiPq2Q1mMjFvITuFKcLnQ
lwqes62AB6q8KPyrtLA8lRQSw5cW/7GoGGba6MM4cxP3gQFIbrRWSBhxrxykyjotOvMIz5OKkYXF
tNL7bvtugcyFpxXYMdwEXgtNh7faIWpKJDfNht+dKvs4LCLThiFq5lvN8VTPZgTMC5K83m0aLSv3
TajF4qCOvJkecvXhlRVhMnT6ktHB90bmtzfoN6BvJUbfe6PEV5p5zhJ9ykmkLB2Hk9Q6GSBzmcbW
kGNaxPkIEFhufz43/IlHoPeHL6BtN8zuqIdKFwrFFS5rXAUjxmK7v9elSHRMGFUuz98F9b+M3vkF
R800sr+lx/GsHMJsPHpptq9iGlZ+69HkrwM8c/DNMR5zn3cF7aXxeX8xDqKCEEMfkE4dSACz90aO
ORsHC9Cio3Yt1F/E/uD5+IL+tD83Fu8mKUvA8uZWmu8E0jRB5miJdn9C8mh5bYrw3EatsiwJGHRn
VWZZgAjY8zy470pG/m1/kLfK2X54qsceFxKstyeLQzOlCe0DP9WrxL36C90LUXtXXsBtC/sEjG9Y
Hgx9BULiN7CrRUIAGHuuOPe/Dp0NBbWaK2aH+ZVSm4QZs2r2S3nKrp9HqUmpRxLXL9bQXXfGOLpr
9BPtD2Z9yCD1kby3Mn19pLMI3mEzrCL8Y1ub3h3S0qWwW2H4v7Z2g9YiLj4PxjyY5BH3PBrqDX/k
KxxkaXcFOlrtxFN3bGJ5msZyObE3+lEeSo2iUdekNswQ/rEKIkvwCkhhGnOTASEmAd09+DJEvyL6
PB2sBZaEpX/i78ET03nnyBftrMADyJ9wRfQ1tfwbxcRE3jyHMiej/MMPnvA3kM9iaPiXSH1JSM7G
99hq9GGI7OZ6o04L/M/n7dk8wPQdID2plOh82VT9bTk5MkwsdVDBwOla9m52TusoKjMnLBoqqNGG
x3FUJNskVUp8ktcCwd+D6yhAcUnURuAfhvuJnmazeW/0E9vGLRjaWjzKOdmX+QTXTn3OqjI0w/a0
fc1lSazR0PMjCnV9HTCYBSC2t+iA8wdnWpdqu8gMniLFw4UzhTtIo3IcyirdK2lQ0JD3JcjtP3CA
2VMXGlzkFUMx/nL7hrXEZ8aEug0ZXRb0Llm4lIhMmp4zk8r4O11enQ0kJgjGwgXWhp+0x6JuofGM
Ztztg6nDu7lyF1r0zvv3b5WepuwEF0KNZ+V4+8cBmai4LZSKjnzeV1pQIiThKq0DFcjWDo5hqkGm
fjPyN6IEV49iPyAgOzluaY9F9V/jJuILbxp10bEBN496URreseaB/XdberH4urBgcM0UVtU/oo6R
6wDUWdO6BawhNNUwneb8lJ4N0PrYmsVZkUuYOIV/6vf4EhsXalP8hwN+Gl6u093gCmfR3C592zHP
cboRh63O2rMvkQJy4rnkZhlvMxs4BIZ0aqmRaUKggDzXsl0RVAeQsfali2sJg42GklOwaeBLQZ8W
NyfKD8O0v5OH3FEey0C7aqWb4pn+l9Rs4uLxOPXQv1FObalX9GiJ+Hj0lJ7/hXhlTJyECywoN2bw
cyjSg86FZVh1Y4j03QJhSUYKsb3xuddCw5oeitafYxULjZye8trSnJPnhkjNm2K114JaaGSOMIz1
zdobWOI1a8W21r/prRmv7HvKE+sIBPsGkc2ZRButLjq31AnOICTIxNoZQii8+C/yayJh5tDHEuTA
B56y0xAhCFXxqwx8+ARgM8buAFhHfATavqAjEw0j1JyHW12YIgJbzRONlgWVKp6TT1h0WpBp4TEQ
dl6RFJ6attKV2EbCGM5TNV516aM9xk68tuLvy73BLpxCGonZwgc1XSygfKr8gGyAfPnc5HcehXY5
GO2ZmeSDiqKc+V/8Akj3JQj9uibO7S6wWF3fzIXeRwRBsZIFhvuz5G/eK0e1qrG8U4yUSQRYyRcO
MOwmJu+zHpx1cR9Trdt28vtXTolu7XiQAzYxL2sdmSm52L+BU7W8xzCJOY6+Ti0IMYhGLcodwTnL
Y11q9QMtJ4IYJiD+FMpmVvrc5XljjSEhZ6K3xj1g9A1RfgeIyo2T3dnATbgCn9Rk2K0NG7jOkMvH
+dzlQ5NZBqp689I+TLnGb9FuU8HqUlAV+MdghZwFLJtO8JMWpKWhg6uOZW/tCP2N9xCHDhEb0azg
O8Aivs6SHt9vh/z2D8x1q+ZPR9ZCre1o8HIYRIvMTWJnyhPZ7BU3OsSLXW2ftKjVbUyLUsxQ++tp
PMFqifSs3MbDCc16wiFviNU/5UlPVTdFCvdR+U9NK3WLmHCpIgt+W5+bIhyuH2PElZWl8bLlpmFU
2ih2Ecaneb2VYs/Zp0PXmP/k9jCRTbJyS4SIqpBoAeXq3+lF8ZyfTuQd2C7dfq614E4j3BBENzji
HEbDI4BSbuayKn6wmnpYhxV6WuPCGp/6uegOGvhtK3sqU1M6qHAWRXQKXBFoyBfxhAzbDrNoqGVI
YFgBwkRY1B/1wEjKwNg6/URoPy5h/aggIYDx0BkYDXyUjc4uNXUMlhUJed6LFR4rD2lTn3NFTXga
KHmjQHQIkSrBFlY/3tpXdt3jLzqqW+8alzzAmgy7vZlkZVQM1/JoQqTPz5d9GoR+dvcjtamIzr51
sAnznanzdekmPxD2rSweWDOSqvcwEO0e6DG8HX0MPTnwlywEUpV+rjK5LCS/EFbTW+sXRMzAyR0E
+B+lVBEHaPlUiGVzhoKWJCVy4wzyh0vvUmN3Sneuhm0Wo8ZjWMUPHFtoZ19H9kUd5udnAZeNgoD3
iq0yn8gmMi64YWbJzpBkHvYzEU/rLzg7UUrCbRr2vbMHdxztvnIKu9AeP1KCdn5Vjf0IqJQ9kTjO
zxIHW4lZvgV+yypFr3ArPihhfdgnPUmliMnm7DeIsJOkto9Or2AlTAegq+vCNJdYCL3OjrzLlAVJ
Sk5MdSVk7G87BPrWQM4Pe7F63J2xf+5lDjkYkZWkAv5zEhLV0FcQwK0s1+491TbtzcOlx+AqSnor
ovjv7vbZejAfRxKYLQKpFenn5YSxBDjUY5d1/9vp/MrKii+uOyM0hxmWhCZHryH0mVXLSockDzS7
AcimPgdvqZDMhlBIrxbOXv70PoKI0lx7pqo68V0PGdffttIzXx7rOjqaGqVnRixdLmGXIqwNFsZS
ez8FdUSLU2uuNHAWfrjz5XNSvh2/BBaoRPAkl9ZXL+uV5VYARYnv1f5oMjw8pRvFSfvZz8B/xxwN
8zP6tWSWwrGeO6N1DO6rLGTFp2Rf2duKrgAsZtDjszCocm05HNCSs7Yn4do3aJrPoWg6cSRJsn2c
cv+BovwyCXTx0mLqcaA6TUrqOcrI5tzTjSwBqpyLhB0LCvsDYlmzUqOwEbk/I0P47lKarwLz5Pmp
i3EMDehnLKCM1qrfa9JK1ycvVbvqyiMRtlY0OTzNYqNKewZiFHbic/EtDfUoRdwxCrsNy1gh2Psa
2e1YMcdxQMrELsvRT0QE8Ry0NOOY82tRARettNeaH3mcQ1Xo9cywBn+xCR7coN7Asu6GfpPMobc8
p/s7CLV2e5PHAsGqWeB9NMW5235jBNhCzMFTiWbA1BED81RlZadBPBUkixFgkHuXoaE9aDM+oL+3
Asq/s2LKyB3ig1j8KgoosLz3ubk1y3vuTbYrrp5lwtwKiPSoLaxUZMsrmqatMAWm4jJtKvH0RI+J
sx0PxRLkYJLikyoulTiLh4hXINiMACJrWG3jsCOAxMvvq5Xv0jww0zenF5eXuu/OXwUD+C485u1e
/g+ZyRKOuBLqqgexnoJvp9MmrYFs+g1X/TaIK3auLxNcU+rVILaxHx9o7NNopAH7me0P7sOVDYm5
RaDkQXso3r5y0zlfzbz05I2/W+CXUHS889XS0cQSONHGKRk+PamzQnJoCtgnyQ6Hy2hbORbCFc7x
Y4o6t2wyP7C4AKxLu4Ku+GgqcGllzgRxN0Wec9SnUSnj6KRI+wYJeuOhCxkzjqEA+Rq0Z8zvh5wk
/XogaXYXY1FigXuJrcoJbvLm1OloTDQNHh+TbZVk6I/1pL4ByvH4X+vuvE2d9DeBwlyHQO5c/2K4
Z3yMTSrRlJtoo8l62+Dxwk1/OjHrZJ1Kg8N/X4ztjLeYyVnf5SBF4aMB67kvtYmC0fNm4gOsX7Ze
rTqowsHI1367yUx2tISHsKc7DoOlwo/aeSd1FBjF2THlT5UyLuusAG1D/E08LWa73+KNgEkfZVyS
8E9LaXVLJM6pOBlQf3cWNqCz91AQCWK9+LY/2jPcqU5bFHYd8iDGA3KVAv8J5l412w3d5UTDfDY9
0XXiPFIYHaEI0XKUEJ9Bv6CiJ0I1X/b02dF7Cd5cHt+uk6nobMz9Au0ogiYXrO1z0PzCtlUoeRH7
cy+NyepCPtneQLPeShUWm6ESJEtGTsXYGtJ2DpsUfwW70DLBcrlonUFLiWRtwqsWm6JuJ70xz29K
KDsML18Y9sA7QEIOuumgIoIDRatJ8lejoxOWUWUrcqY0JHMr5fG176U5yImmR8KZKFUYytOi4gXr
ilKagbTahXFpt2olZHXUOukOYqyZwBksnOGmwJoBEqN6SBk3nmR3p8TaG2esxX44jhzZbqSMEcIt
BfPg3bCXiudTfRqGzs5liE49WFYIBropxXIrLVfkIoWyG5HQ+ojplOnBfoQK1dH55aur4ULjQVVV
CNBBmnlry1t00wMrLB/uSkZwsBK2T2KggvhhsJQ+GdjZxC0mlmCtC8O7x489bhkbJNCy21xWGDjo
t8rQSsSa2mZxcxDRFGTLl0KsKNuPB64jwCHgb39dKsy6zbMU0JTOFXXkuIYF3K5tkxdZwBYmH50Z
ejVsPoAJ5wIaEfJymxluTlVynIR3oTuWa8D0fECMJ4OPUWPKFyhkst1V74elQm6qcsXuRJRjf2il
dvQ2we4c4kaG3aV4ZSyZycdka7NVUZ/2NzUYlzchOwEEo4g3MtDgCU4AMdbi2E+GB8VHTKH9OnXt
0D/l55RFnubbC4eIc7D1ecr7L3TSeCd5zFlff+UEyUi/hdWiAvCJpcdx95Ttk6gzgnDFL3LD27Kw
Rn0MAJwh+4oxFHGWgqwqlKbi4N5zC+TZ7c+Q/EQ8svYFQys2zenEmxGucMRdZ0PhNU1Mij54+Hj4
y56Hot/JKSkSuBinWJXy72uhCtZA8cpa8zRIjK+lT3IfaT0aU9SfSmMQKhKQcaWWiCPQNzRSrHmk
wW+DhhSiPR19OocqtUC+nSKDxgQr4FK9aM9b+jSkKgf/hevlGMoCuQqXvJHr36Ti6U2JHrgpqQi5
uUTJMNxXaPEihtptMbMCpSCkLJBaJmoYp1eMEd9XitTBP1ob3T0T9vjymKnNh1SlOAE0bT6OiyK6
+H4za1rRG31yxpmbVfokF8AVnHk5wlJKdLbIB5I3jbS2qnpTbsEKj9rhEgU/HG7cHbTwmZNv0E/A
v7sKdqtHfO3NoEv/qwoGL6WkaRE/YwX45VjOJPExiH7NcgaEZulHh8JYWZOdEUShV30GiNFUeWdX
kSr1llElhT3Liibl0jzsA140bYIYFfEQ9KJyOqJRLNhymoHT0WaPeEC/moFXQSem78om+PdGLerx
UmTdnm8tiMkE+UhlRuF1rbDfuZV+IB+E78oxFEgjAGOGQz/dFzyT5K3uUZ/1mufgvIRhkGohP5Uz
C6BYT9TFIpoJaDDE1AA3t0fIN0MFyawh2af5IW7AILEu4YPPOsJUHSovrH+lAyMvPfVyW77SV29G
7mqiGyhkzJO5vOpkwksKMSWovlAwMVVHZh67ManIUZJs5vmepAMQjiKOIPLdLXCxhfnZbn+zicI7
Awt9Ttv1ZPA2BSSGWFt1ifXIscYRp2KLqOba0kHd5Y1Ind0qrZgclYdmgu/3k5k0P3mfNsOUIIEG
jSgqAApU8io3AZ4ja2pP482PDSpjYfShidsaWcwaKklKe2NAbTmyMzob4uwKEvpJ51S9mk6nZdHR
ZT4acPEIVA5Ci3MFd1Q+4nEz63khlAgH31qYvw0LwhZo9NKo/sRrWjwkZg32+40YyPbNb03P3bMu
TPrVf9KadrGplQpe6Pj1bZksDamq1oc+Z6aN/seotWQrQSazrCuemgG8KTpwBW1m0su78ykA+T5e
TyTSgsypu6GcaeEuN0N1q6l3TNMOySCB4slGk5702CrVZI8FMgAWgXIn+s7+zX/gX4FOo5ZnqvEu
T56MkYenkH5VrjlT5jhYLntcSpzz2UNCXx2AlEwK3U2jF9L1M04o79IDoMRS8/nds9QDcqJBgpUq
5IwAG1gYo4udmd64BqsGiepKbATf/OaLfiRHQydjbg215LPm6gjCA4IbHXv7fgf0Ifc1cPJrlpsU
4IQ5HDF47hw+V2meUGMHjzTzHPrTUaZVzngHl88R3XrUETzeejEd4bKP7l3fGcFjI/QxbBI9FoxD
PePPoJDTC7W4CmmTxUx+u451n7yVTxeHuo3kMr1pj31W4/TbbPGi73sKMkTMQnQxtB+d3ZpQhAuH
087XX9a3RIfUWtNxPOiv5fBAsu275EpUDuwT1i73g/1ZD5SOVunOMz5VHWVddswOCYdGjINT8Ygi
9pHq3M4ivvEafPngnotqW0Cvq6Sbwd53UVKCegeRXeSxVdwtBrFNA1mPKMq14JXDu9u8DNmuSjrT
NIqFLURAusAsJBrxKkfplw22PE23b6+HUSH6XxfiI5X9XemujsaBj9aWGxFielH9M7kveyrdIPCd
2elvrjHi5+rHP3JseJT2YZCr+FuHJjreYa2g85BHk8SHio4Kv0nJ6fGpiUXhHIOsci9ZEHmKldD5
v8n1I38hP9Ared2rea8XF7yztx/Wc5NpMXeKuzSNgziyj4/N6kn28Cd+pLW/3tMW7l+Hs/0VuXWZ
h30c7aNgRPmPEFEkGOwwfqH6lrqc0+l826W17REd2HX4XtQd2b0fE6OmrV2dAYjRW0BbiBs1sKW4
0KFIonrQ1jg4PUv0bsEVXjw34mIwAWhOlNZL2AU0y9s/d4EAW9lDIEjE84GakdE83BNLtlQgWj44
CFQztahFFiU2tjppTfm9UDXhHu/c/kjdzyED94TQLyqVaF1QFQ/s7Hzi0hgyHm8VJDafmbTEavMp
LiQA7hRhgqB1zso87KjKLipg67bo3c/f+DshIVJKArJ+TxDHMSZ1P8XXkGKc0SPur71wfCasvyQT
uw/z3GLFAiDdmJT365QeMVjMofW/wbLj9yRyhw6kPJCUodmMf6NTxpQy6kjV/MxEoHQLx2kb7b45
3GNezZhYbjp6JPQKbMDGX8unqWT4uNLritwww+dWzbyET6IRP206254Bi1eBplduIOSkK84ENrbK
8Iip6kCyZ+qyCO4O8iMeTtaM1dP7JpaO0P3wqign2zQOS/3RjjohddpEi5/+HX2c6bK4drICUX/Q
p0dpLDqHrmTAkEXbqY1kVvl5K1G0QQPUTdKd72TzM/IbIVmTnQtlPNy9Ck4sTDmnN8VQ9ilUeuJ1
Z4yEVcqdKEMEmeHtpeIpJxluKFGt0b+io3fPew0XLUUhMMUqbyZ5HMNuLB6aT4lkgdymJgIyko1z
/uLgHKkJzpgBvtfq6q05FZEe8IYWergX+aJCmNosCh58Dv3zehSFHVoPmjDnx1UD93KJZ53umyYW
oBjJ5EcWjAgif65kMSyyyaB+kM183zI8eCrm79iWrOp7Hfu4CHfJufQ5i1AOQVZld6P9k2hHT069
RjVIzR440B7BglMALnzR9RC7vco7/j2hvzESkQY3AJH+U0ys4hgU99wXA6N1lW6GE51eAYs5fEC6
YH7+oDAbiGcMuezqOOwSb4uOrqGtsbO1S7CId/PmN0UgV+OYPokpvH5UuuS7h4lT7ET5XNZQD88P
4pkxBhPEys8YMUpGQc5N038osiwsReFZBProIwUty6tIpM8K0/ZDwbniK/Vn7MUMyGuqmgV+Vrxt
ged0NF15CVbUwIVnDrjXFeeKkACKgaU0ZGgcArHxoJx8jhQJzJjwGhbY5ROCaBLewkQHy5gg2Rz4
RAa7vTqUUEV1Z59UFuwbx/xKCiP/OO5F6ggpOqfRd61RRrM2o7I4czD86fUdZG/i8HP1JA1w7Fq4
k6ROMZ8JTSXPKneclorCvfhauwiwsWZDV/0QireFFo1q/RuYF0G1lBinYH1bXz3W7om+M4fDILNY
NPr5CyLZ3AhhEpck/NZ4EB+QaRVxv8XOmja0d1XO8xB2MKwxU55KMJgXUxD7HtaKCDBUY2mS8ZyW
N6Ob0VbLB+BU6ZNvUQsq3ZUERFCg1n5cXA3TOpVhr1anyHo5tfNPpXY+0isvoo1EwXpMlKphuPT4
349w1hILt94VSsZHF5llk9njRfplPn0tNeQ+WCw73OGLWIRqfP1Ai2DXVJIEz0JdaUTRb+3/671d
e2IPftKsKHIWbnEwwQpjBavFCkfbn7hcGkZ5wacasQPkDm69egLhcIbIZHxszX2rtu1leoWDns04
bWmcdv+4s4XVHxPq04VnRbDKnCH89eo9Q7AUQQ6lo86vhdt9TpIiUlxXRQFWPjTKW+AKLeoTcbL5
P2Bjln+IzourVt4vnJSTXOt9RBb7p87rZmgx4njSNEAAFz/Cl+HrrH5xfJY5cS64TmhyuX+h376X
oRoiPPinvVhj2cIvNgw0SXWZ3IooyTOLEZjx9GzD/xpXW8nBqPzyVqO7XMOUu2iYqslS5LYWUZms
f32E35guMz2DpiSvafJwDjLLemXERpLxr/n5Xpo8hPa8jWE4GgS0Fn+zJ4mR+24P3Qnx1vGiLqrL
tnHDrHaaJ0EkpxoHg5tyqnzsel+nvvaXdo+XZX2mOmPX706jHmuQZvlpLjskBTgiz4Xyv0+EzOwV
twrIEIaXPSJmMV1MgCkxwjiJYfEV/4qXW6iZAkHQyFpQKvUVCIXObRRy/V6D4qGgexoGuE6Ato4p
qGOr2e2i+T5C81Xmn+MjWIeZDEhSyCve49gB/ELPKq44XNMAAbuXJc8pTw7hGqnzU5m43Y/eBPWJ
gm9vzWIp9puAIjWSoQ6ti/20Pr5z7RgAYQZULPdMmAe1vrXug8VleJ5xn5rDcNz6ubniJmiTUFDm
04SGoxT4Q7JhzWiCYeAo5XbRbJ6nmKvSXQeYLuA8DEC61hnbxyt2Ij2Sn/VCw4Ay05ryJX39rJgM
m4VcyTvuVimn6ISAn4irTC4ahMO4OLGP4M0PTFYW1xINK6G3Fgy1FOrvfd6csyOgBagXFwyMzu/2
h9OVMRme8Kq7j+ZtK3NbFIIAMP865aCBrGC++X8Gh3HXgkh68PkImvYIrnRxfmhtNvdmsq8l5HXz
aiQVozVz6KxSRcpnQM5SHma0Nu0j84K1cmadQjcWEmbkxnrK0y1EfAlNtuc4jCJ94DpOsCreT1r5
ayh9faBtWBV8ZT2eKa5WrT2mX4LmDRY1hB/p4pgAPEnwGEXx6qQnZD/dVeSlUX6yIE2S4ne9DRmJ
IpfRKyyizU2HYLxF3acYjnBaxUdb3mG3H85svTyLkMb/EoZn0+ONM7P7R40yciBwqhWWvGw91Wj0
aSVe4H0x1rcwEXz04bSsC6RjOjzdwB2yvgM4+7QBLRDq0bBHhtVldOofnlXiSDwXft7vIzTpGt+7
uVoyEy7Y7QASDmb3H7YfbqSrfUYCN3gq+7LEOZn/B2fjzG0jJHjPB7KCcZ4eDO06SMvYtvgeDjol
lWF+1SeOn8DDERhkdWgk2f8k5WJj/PGgZ3i6O/u84BtogUOBX8agrVOnmjICWkHZ9VNADJQe9jfY
64u1mAA7fWVlZV3Lmq1+Q6E7DtyC7JOsbn6RDoZiB1XRMjAM4gZ2Ttb+kl2ukPlKiUCnypZ6QoyJ
PlG1+1GCeUtNSqb1eLDi9liIPYACLu0loMkYWFb8hERGLHPgaeRt1AAlt5433hyxYk78HxOEkqfA
3rXI4IiXH+e9WBNU7L42t/6hXKcQqLCPFBdtYtqJb8bFaYEq2OQyM1r4b94ykPpa6QBXOYAwQw24
AfQPo69CEPmQSqHEXp41EyF7AVg8Xpyl2gbfUUPvW+Rz/Mawbfu3NmeOBQ8XGP6FvQjzvxE3ixrv
9JRSCgZjU1Q0EPvqCRlTl080LNwVGcyh/MEQHr43YjmmfjoWqvQ5+RdgoXmmzlFkpWTqerhaOI9b
rtheRGue6hdHcijLZ0xajb9s+bBfJEbJoDGIHIcUM52LSTaXAvRG07Etkui72S1wmtq2oemVdeA+
mFSdGvsCxoNYrn6QFmdtSx00AI7IUaCz0xkXPZ2+MXYHqszxQSXH8XVfAVoVCW/E0jU5s+J6iPSw
2YfWB/2j/szYUMGKs2zrWcBFhxONeTZ5yDhyb/3EPfyInTt8WxUzPlRzQSugbDqK+sD0wNz9krbl
zvVYKD3YURzJvRL+aVDhLCjOz3ADVunWvBoR6YaATyi+NRkL/nL0SyibRBE1sQLEljDthmnvwUOq
gSiQKAtbyWjJu+OX6BPWgTwRrmxCIGRBGFuRgWh3XU6XeKM4Ft8UhkirUBCwSTuj+ZTdVYr/OjQD
bV0WJdb2EEdfvFGAIGKKYRX6d0G5Mb23Si6lcwobTwAXOTU1bgzWryHhSlG/PecIfykXzJ0G5cpH
KXzbiko8rat86Oa3NOSakqpSpAEh2pWJHUcPJoPKN78EbBitkd63kL7+1M/A8hcAuL27P6eov4pJ
7kjTdoh9zQD264h8rq/E7wE252if2X4iyTGwstZPi0/pCjB/p/jxWYDqGgKtQReoQAIszqaohfz3
zvkW8ggYBNueAzeBYXV8bIuRnM+JWatkDEqmtQXo1BNGgfTROS1LueHxvJ/+l1ERwIFkxsRhnjV6
Yb3+N9H/BQBh4f3Jega8eRG9fl+Ml9ASBqeOUarxMWgNxAXlFLxY+Zxv5ATBfoJANCwsCT8QfiFV
VaCvzsuELJi/AlEkgnBGAnFEsFXww2swtRd3sfH48UWnLctQgK5yFM0mzBsvDYeA0sjWD8MYBdH3
VoZMBePGFpoioy7QvzMuHvra331PEUhpjcd8qQVDZuNLvf9xou+itXzzBThiWD9YLqlvVOCWC/1x
kA9eSrhxRQaV/l9LxheIsbRPfARjjEwIH41TGFtTXccUCBEGGrXiFwWJYizEP0U91Z9KWnIF2RLW
IlPzTQROUGzlNqHJhrSygLIFfYBNDXjwPhl/nu/seX/rS+Wnw/6si3cc8PKPSJ5Y0n0oc9pF7Neu
cDxAGj21mpd7Q5+FzJKberhMaKR7iEoLsFsyOhFMEYW3dogre9ZgNN4HqMRGhIFsBeWVaS6rUiXu
Jh7DxoGAvN9pa/veOCkaUdkDs4iWlnSspKuSX6BGov8wO2iBJShb2FPOKtlu5EN0fbm8m/VpS1KR
X7deqXAi3k9rwhOpIcR5h/9BWyEihTcjwKCrU6t9Y1L5OVtouBh59EAlNTnO455BBwWSK1X9U0b3
PwAOYnv7wDF2hDHwEacZM4du/9361fiC/jAGTw3RIkhDx/BUPJ/RDfW+BVue3vrigZu1x15tWcP7
R8EQw1RAF0u1Y9Sax8VR1xX3YPClQFpVhKSNCtMBy8o9mjNQRixY9lYqttDIRKuiSSLaEGsxAEgX
FV2a5oi0IMqIJUSb4eK0P9q/5XZY6yhpieU/U7atutNzH487+3VlWMAu3DmKRF7+K4mVAZmg+Trt
7994EpjloIqPE3p9YLwgEt8J1AYXC9Xz1jxKGCZbgYsDKnY7fm03+nqs5kac5lzfqyk3b24kNgvv
GT4VwioDA1ccPeXMppisDYq0BMwijTuZ8b/0WuXd2Ev6z6MKOGqAM58v1YI+SNH3MCZ1AcgrB4Ne
lw7Rr4A5BPlrpISC/lO89KulYyQWXooNVuhyhn2HWgWAxLG4iMubIbQlCZ/lHei0Ov3o1atB8mA3
z+G+eP/MMexkN5oiV3cfUgxoGVcB/BBDLbhWHg9T1r8HLevmNNJJOabkdK08tSwL5O4FKVlN9RUt
vjATzfAd9HCK9mOZGllvzfuWHVy2JcgKdBj2RXwOTPJT2qWhExFX8EPwNVAijiB3yzgmvBHyCS8A
I8K8iZ4rm4PLufUzpnGtHJmF70w4dNFyg2PKAs8gntvYwNDMiaamYCL00x9WOT0yZRPnDW9kjrb5
G0YkeUskRFCdFIIRCC9ioT7hFR4o8/QaKK8a8LvdbMp0omQinDHskLtTmftPwCI17KGl7F83bMGR
h26WQR95nKgYqk+FfurDspy+1wv8s8zAM3flyiu0v/MRdYDWFvJDAxFViS92Xjj6ihepuEEt2AOi
Cck8iDHhai1GeOJY1+MWEkhRuJSJ6jZSLI8QsSnqCLXMFtQ/Z22c+7ANN4fMY2tX2oiqpUk941vl
jtlLZHTaxGwFY5TrWVYceIJp3mFUKZBfM26wfZDa3BahNRUywnD2nPz4uSkWbv/k20K9hTmtpPac
FKzqW1d74c3aickcmsr/dF72rZG4bxqoFDSKltKjbTIdS96K4WGDm2DYsOOyVcSriV7NXqiBoNh9
orf8ECTE32+zqH0WpvzxXZLYA45CO5XapKKLt2ADDZSyjEdfiIWqf24cmTk6cyrMA5VLXIzUj8qe
Az4mwRWAkU2j/fp/lOegP3ZJZs1zqv59VzhvFxlJz3LqEZi5N2sQNSYCR8qNruSSgKTxIrwRo38r
DC7Nt//Pni+1oYx3aAVS9LF1TW28GBR3t0dXAQy03JAQazvrEmw4GQ7Xt6liM1eNQtfddlZdaYQN
MyvlTftM9hWd+ufVq4ORJ9ZDjVTewRQ6mOjL80ztb5hmn8O6qupTPtlxFcePFUZESHFFo87wMETl
En1PvNq2OsgUf61/fN8GeAxifEc+F/YPFO5bUYb63frWb8Wgn81a7K1qWhx+zFJ2cu6pI6Dw0iev
e72g5qEk49G2ZaYZ6lwENENbhiboRSayQbBzzUq+Il3eeiKexacIZSI6TOKZNlrvGHmbhkbW7K/R
pQ9xmEh5v8/mZGlAo8fy4VM0gULI6/EXecEmNebFuJXBkrthWqV5R0LDuRiKkLGgNpUFbwJnlM57
VkvTMimsbqj0abjW1WxOALIgW2U4FMozTAiKAGPCsrmef6melnw4lgOpVbkT3Wun/81oKZi5UAYJ
lidsDEIZyw8BUMUx8367rZN71njM/puZ2vwGPGdWpyppW/gf4pJt9k81QMv5cJy+dj2QjsUn50m3
UBLkMyZDJx69NF2B6VvTevi341lS3SsIBvzGc39RI9GTMOF00hHxvsRstZbX+bd2gxF2rNdUeVLY
xfk/VS0uACNrbD3BxYbi78sIKqE9PuWoGoiaVdSAxEe4rOu8jThTBc54izjlqoJJ/SoDIIniyXAq
Otxq6qQtsNyGuKSNT2cRqErvNBSHL48xrouOmpc7n/iFDUDGsVLYHiA8AvqbtRaNFxQdcOE4pVpf
6X1YibtEC0SqaOVfnA33zZSfYkmyqRVKcwLkeVP5TZtCn4W/D4qbTcQpSS9mbyKqkn2GcKScxmX6
+giiWopW8kwty3JejKbLLpYAsKKjK3+zuvr+FVdncHSbxCUip75YRv4jOS4V0NiwLLltv2tFqp63
owzieewyepS4tMzWiVzgOy/IgyIdHJFuWYXuGkiwQy0fpD883epQ/5uR0wLVKWP/3p1PfPFzrnFe
ZEbVjd+s5xi5S1PrqZjTLyuDfXP+EsEqkBO+dzP7MBfjbJUWlJ45gLf1Qy0TkwmHw335+tTxS7dW
MSj8eZT3PQe2fBekFZlsIf9iegehuyKPy0lf6D+CqIUE1ysSTA+pMkyY3IfS2/rWjgWztmi2JDvS
DXryaIvEy68Sob8bKJXMtNSKYp2XRucOiGEZTC8hTLzFuwQ5ItX+jN6MxRRRWwx0rIXNA8oH5ZIG
gfFk+QorxLmCEEWz2vX68+YzqDVk1y248i8OmZzX/iXXetpqTuLkgTGCkBHDIJ/Pig9Im9CpgBwS
itRMnz+zd1KnpVaPk78XzFllANWcaxSZ4zEDhsGyMs5cApTwBXzVoQB88pbQIqcpDEZAfe2Q6QNo
9dEP7am8H+4b+33gVhk5AJWoHtocT0cEBjiV0llgc8PxdVX/iQ9o1W6vb2Y1qD+bYpJTrZ0t/yKO
tI5VTAaNYpT3yLuYdW6hlin1uyJSTjjhLiCoVLfoWwISvSmcVLvTjW866uSO+y237dgW7EIFk6YH
qjrDB2+wD/Zk7EuYjFDQ8ZVww6S2j2YsUBtJxx0twk0N5sIt1LrQC8GWgpaFgHBKDL6tTX1f9BbD
01c6uHSAdcg68ysL1MsNEm+S+sbsZ/Tbdfsxj4q1T106hMtL/UBb3n1p99JbhmWQ/CQjKfFFzl7A
40t6R4uWQyO/rk/c+QEP/rgGLXoRYqnk60jylysuaTopeP947n4sb8lwbLyxVrU+V0ydGe8T8dnO
f2AGAEHpHm+ZMZ0YmG7Vgv77DV1yQlGqmFWmQgVrdPpYMz+8sqO6Q+fYgm4srbOkXsvOm52wreB7
WFVA6fmjFSTYOM+Ftou5eccu3lfSWg6Sq02K2y3ZMAuhFLu3ABhO3nX8CnB5V626AvtFY8kffG+L
qdK5gGy6D5ni/M2rX/xJpaaCKcxA6WjUlgFQFmG9TiDeKZy8g/96aYeX6yCQT28ELcP1GmCt4oqj
Vzfnc0Vp1nlGmZSk0sn92VA5BB5S7kYREwuIusrOF84Dj4X/rUfnfi8zZ/VYVJQjWNZonkpBTBad
e/URJ1AjP5DVy1MXHiuvZ2k6+aTkErfkAjyL0757fI588HuL9nRToML9M0Hsd+AKMULqiqjVdDi5
aissCIeEKH9srElreqD/aEu8rrMUVFMvFUv36R8lIlrE6IwJr5i3Q4EUAxk/S2fowm1Df6uLGdo1
Wuhe/o1srUuaZgIB0fZGFJAOA1cNUkUcCFtslD/+uIQJ8KXt6xHPaF1xzuGLSWSPkI1HZAq2lyir
miJgiGFO0hbZKr0vVnPnMiElWAhRb1UL5E/Nfie5b5EkF8dvzQO4hw38RWeK+V9/pG2yNKxTRmGa
c6qucqpX8Con49Y0KrttaS0yfIJpwVoENXv7wqe3Zawewegrv5i7B09EEa2HN3pgnqD4Ja8XP/oS
+oJ5ec/JoTBXYSNZpqEisYamyy9SD+LNQLktXxSSzfEWnw2yCsZJyFiBA6ZW6CUbGR2IXDaH87Uw
tnl3QyBE3siC+gBlh8cKhliB8h81eZeWvFKS9fK6QOHd2YBj7s3FI7RZ304OrbpJ1SMkGzYymP52
G6ksF3LWyt392EAtobPoVK4DRszbU0Ufghe4INGLLcdPShvfP97DUiotz30Pc+oTJ5RQyZ4uXRFs
1oHeuKqF0MTWgTYZuKMNBO72P7PRwkCUhZjCWOGQ3bH/z5zJbQQ3HThFwFDGn+23w5mjSgJKDm5s
YEcru0m4hZ7SmloRltw/4NVsUl0v2npqsS7whU972Zu4GE7xNXNfEqOsbcGR0ztrPfIeo9bW7MBu
RA+xzM2DKy+EWaxy8c6q1lsjEQcB8Bk1b8TQ9v76vHrcmuvh3vvuUcfZGcw1hJFRHMUKbb39EvZn
aY6uuMoTxn1Gx1CtVoihERd7hT5TI5tL15OCqNgRp30jl6G2E8ggs4a401Tw+ZR1lnLZsHbK3e5U
iMuI++C0RQeVg60Hym00bzZtd8AvxFax/LenCTUHmGCYLrTVwMKWaNV/a31gSUuN2jlL73TS96T6
kYE7X3ShIXHRIMyZRQSywdwZeQxdZShGMQx5bc65Ajnkf25luZIQa5zjbVk1UDywjp+H/eCbzXoF
0trSKGIGnm7UATsovjAomnZTEbGymf7UEN2KJY0qGoghYolTIClmHwL6fTRNMFkae8lcDi7sOyMv
5A3ec/2d79+QD/re2lejHwVY4enoe5mlo56K7wqfD8xq4dzK5XKgBlDSnvFrYwiQWRnnfaGMtN5R
Gxi12P8Q5TugHXtil+TqTuM/+wLJ8Obef1Q2ha5SS/bcoL2LFhwdy/0nSZX7N2sNgh43vYpEBXGk
P9R2yK+jNsuLrC+Wz4xfOmz1A/vaFfpP62FGuIBY5q+05lD/5XF4EXfc0yjbMNUg3Hod+uxi7VNB
PlMj/duklFHgpJVukwoW+kZPRcIWrpvHOHZUKadOIPsKDzVLSSoMqf/F7+SiChPBkdyrHOy/VCeM
IZ5UC3XH2B2YZes+jX+gcJI0DVqgIaq5RsxYG2oi1C8LgeqyTtXsTDrR0SXo2WHR2RDKRJ9dw8Yb
5QrIuvriTR76HovwKXTddWBe1wMIQVb3FuxTyFL5hp0nhSCWeS0+gj72Pwvw+QuJTOho+gi5eNvR
0lVxAYOKK5G/X5U18+07uY/FpUTT1nukYYujCkMajfTtBID8a6Tn8kGClE8vftfiUwbjusr2I2nu
U5fv1rnAazrWmjGCnD55NKA+VSZHXi+7Ri94edraRG3nW4GTnJK0PyywspIxDIBGtm4FkHKAapBa
igP/trEhtmYiLwlIqwOSJtd3OIXRciwjIgnnv634LrovuKWN0OYRIR4bx1wFXbzKarpWPFGwf61p
nNjKuFySqpLmfWY07LMKTq2yBKZgVRartdzjYolsZuJJ9rsCM8xARRtpo5FNBIProrSp0dUQ+HTv
t2KA27BnLr/hRhmDaOHgIqf7YHgJH9zx+Ors3wuZVMWQ2eWZPFQiHOZYTh3yhB1stT7egpGAzi3S
iyGPYV8zWFEhp5HK/AIIN3CtRlO4Es8gXeIRRRjtJ152HFZOS+CpDKcqUGVPZ/eEzIR0FJCfxYbp
NBaCj3cjihZoAFMmNxHv+AG2arG5wQMQHl2Kq+H1lFh3CNc/zw3RY4vOW0oh8saUm8xSBehQR/3M
npoMgg7HxlSvawah+vnlP7wxuyczmh2HU/2ZsLaeMLr8ib/fFvEXc3H25v+AOh6sFVi1hQYuBU6Y
Zzkttbni6NZUZBVHEZxZqKgcNsBwSlrx0nWiz4ebzgkpMoJCVZS7KcjPxwkllLX2eoIrCNONu0sK
ey4Sw76xPn5nAVPvbkqGqVv6djiROgP3EPBkS64ZRl7vmus270J1gZ79PVjPMd5whK1DX8tE8vzT
X2TBygNIBqgHNJ24det/AUhViJa/CFvd2IMknNDhaiR9jLy1x+6zsiAPFNQzrj5LjnzwPo+ubVn6
mGIXK2jaDAyXCwNm/eXm/KkOzK605/5aukwxJ4gObD7mm/WmfkVRScXX/PreAH8LKRlJcoBnrWBD
Lf6GlNPnt8hORWFJjNlcts7IbnpIv//pasgjSAnwGmxaZtcMfRjuuQTRDEsmANU9WSOD3DJ4hTdE
dvR4UQeIFoOkioPD/lz8sLWCIvRS7FirgycXmdiEbe54P821yvtX7xU/an/MG4Xsc9tRTEJri1HB
K8MReig758kdDmToDjYOAcjCyddab3SHZQNdl0kk3H04wCC1swv/nenxoUKdeUdwxg1Aa6MY6Tfl
NzMMgeCfu5SxyRND5RbXnfJlWDK+DQ86YS+yhirCB49e9XsSfTjz/8VlhtKaJsEN2nYianvz/+m3
9y/2i0OKw+Bn/E0TNX/phicmMaFvLUlwu/ItuM9ZHYV2VgqU7Jun1prhIqDMSyFz4VlIcxYbMBfG
QhSnOzibqpJZ9JRPETvX/016Zz5EdKvobqKu/ltA758qROelCZWIO1Exa19Eug0vQn2IDqseGEkW
Fg1/TbfRn9dh7rPE5zQFyfvdN3N1G2kZ2WGaADNm4WrOnsf7MLir2073EsYZApMxJAvBXEOljy5U
T1vYQVWOPXoc+b2RGwhMyNu8uOk/iFpfOC3Oho0Q82J9/o8NPHcehWdO/GY4JEfD9DW/Irp5Rnah
gWniR/p6jEBt25Tet6MySLry5ws78Mv6ZhN37TQvCJfunhju/kpofpabbUbeZADrujWo+aS97AF9
npw0OSfjDgbfsw7aUZJnZbhkBXXTU51RZTSVrb6qcfUFgFxLrBq/92go/NRzYdrnhyrTfs7lTAwH
q9d9EVJAL6UBOUBiJzv0EmboR8rG1ejjLscfay9zQnBNdpnbUn1+tMBAImtotUN5rKY3K+UuXlni
1PnMoLQrzvCZ3TrdV4BH+B2gT2EjZ2pQ6GIC4trc/Fx8YBtir8c3QlWkMnsE0Gs9PZrIpquiFuNF
/FMlwSWpw83y0sS99jQuQF2A2DhrCX+fS7FqHkaj9jWaQkBepv2dlzyZ0a+V0TEiwnuvggzXq3O0
eJTbAUEN4iFGiI4zalG7EuY1IIULWgqZh47CGykiBMjePWA5XfQRm3BjCKERaEyD2KY1Nvya6b0H
hDwJH6t2sIZD9fJjL1FEDpjgaw0Zld281jEhvb3TgJOTMMOCem/F9pg/91KYRrK+um7kRDtDnYXh
g1/8rmqMdWtDaa4ERTqfGInMS/sCKxrY4sei8D/cQvWv+8/eprTvIxhOnxmlsKpmusfDcKsVTfP9
qXROWwxa9vJc0lg3jzz9MgMGzLHF0FjuqckHKQn0VBiX87yojCqPBJtM8Of8Bh2J0GuzGAVu/wBG
F9qLMK6+RzoYCxddqIDKb270ccFTcXn6Kyb0+w8hod+X8JGC8UQoNhgKTqEo+J+LW4rBmaiCxVQf
LYMjwU3J2Y87DIPSOYA/4w35TTR45HG6KeJjCCrzJk1xhvU7oxXo8RwL5BvErwFTySp43ms4RjHB
Pw1n5vw0nO0+TTZtStlMCBeVNgDQ9pcTjqPSCkY9prj4NUePJu62kfmHaUFuogUTN316inS5zjZe
0bsrP1MAQW4ZBHDmp4FNlb59a5Vxf/czXVZ3IQN0y61vHbopeTo2lRpanoE85QtaQSlrGzecPIiJ
L1r33hisb7bNn3UyVlpjUe4LBlqfElNoi3mqjgUcCGAGZmNptNMtFabfECbVvDQCJokRQYMtOMZs
KbVd38UD1lf8USuayITVEaamBqEvfBksdKomWtiaNs8vA83Nxo/bFHsHUJzGUwO8nXzPisKtg/ol
mDdkPyDDIj7VCOnT1pCJfqm0wZCE8xhHvNYER31Dc9Oegro/za4hW7phUyx6yur1D1vixlTIVaY5
3d2BI/It6K2EqKUpiu8QlJqCAlA70Q7NXK9ztkzW5Fhgt2gLpM6V88cBhGX814Hjpt49NaZrAK/i
4rCIlUWOXxxVULAQ1q+wwbEMOswZg/5hvwb2vz1iX2n2XCAMnPs6pFTFiXn2kwgz2jTKZoVCHhwN
CBfcDJAuCu9SBOX5iAtvkd8tW18KxOSgXV5/xzfBRTG6fnXfuG5yPZPTdGTQWjT7wb/v2kI7cLH7
N78eO2CIx/Ti0qBo48Df2goZOXz9k64mPC9W1KIHQS10jz7MorQJGu7NAUS2VJKyM532i81ZJwoH
9B9fbW7fIVcCVpE1ZpdUEuF7lUxsq0UEbOsP7sJwuIdP45SWwVQ1HcWIFN2sETq4cAZqz+dd2NRB
hIO/bd5MEvc2gti7P9/k4jK0ynH4+lTA6M65AtO89ICCsI/Vmxv0zY/LoQkZYz3pjMEwqZUdGXww
B8y+Va7ZOtZe5GkaU/A/yBn6QGVzvDPFWl4zxthHcyrB8W2AQGLtpOmoPsK5McdbywwaUS6tpdEq
fzz/ereQB+xN2fjHICbFbK0jg+B1Pdl2qdt1dY3wEuaETMAqoxo15CjjNug/zLK1aWz5kAZwwRKJ
3eOEC81aywrFEXzU47m91G8Ts2Pcaj2mQHZHqvtzcM0hyOD2QfCawnhyh7ZI66PF6j0yAqJ0FP9z
tSpY+0wEFBGmltVeaGyqJV4FqPn6iVg929ZGusn8HDAkQtAqq+aBLNuRMe9tbGc5+1gm+4JDVnkU
YYtaw25Oa0FfINgD6KRZFYpquSdHZrfSFykNNZ8UVoIU0KYyK4inbxndQJ/ekpVz2DZ8WEbTX8By
Kp5btnZA+TGlFVQNISWPMxdq/oSmsADQRYLDz9Xg2LZtOVIB8dYmCCbHWZ7CR94D43mnNyAzb//f
rZPnvWiBfEL2iCXgbKd1PsuDz5Zxt1kA8xTqOmOn6EGQvCFrhQylA9pxEWpQb95Z0yFokHEXb0ds
/i+/6DtVcCs9zmFvrP++/7uBfmOy2PnPbM7kPdZu8ZSsjxxw+TY+eftPqNIxs6uDpW8YlwFj2ezv
v4qW0zQgBaz56bdwXdEpOkldA6pIPjo1dlEIOOdu4XvPSgHyS0Xz8AJlyTpWyH3THEDTNjkoVkGj
fn2nNcu8mQhXeySMDvjY1pc/UUUlFw42BwaUoKjA3JsG3VK5hcNamzGilqaeYv1CIXcHUsHWHllf
hX89Lwz5em4kdKYsAP9Zq0Pm3Z2rVcbc3FMNWMQZVf022M3RpvP3rNbwxMS8MBsydZrGF9afTZ7S
Mq2YBREMpi6b3GPPL0rjZjx3PFq5ExnV6/IE0Tor3wdHmFI598H8Ow3ahJpR0EnlbF2rGBypJpAp
oRtz0aJoiFYnmsIfZNCbmcLNRyENawOVbNgGi+AXC4EIxcQPVyLEGhyr548veLSksVrp495N3ynF
ynETdJdQ265Fx2fUXly1yTbxBUHnR2yFXBIOsIBts/X3tuVl3qVS44F/YX5dmDOH7f1ITEMRcRsN
rcGfjSnx2jp1/8JKmyYS4zjmvwNNHu43dbW6llyGYi4q1xRqp+iyLF+VMw9Pxie0YQv4/0xYmChm
PDODHT+PoaItT4fH0UmVEFjpTIDxf3Ysg/CFDQWaOu2os/dpz9QSN97c4B+CkEnUFwai9lbnb2s6
bq1kXvOhV/xq+8G21tyFg4FK6xxs5z/KXSxtwfcGsfXDC9JJThN4WyVWpHmnLC4HS35OBf4JQibZ
LZtoD6J4o3VeqgTLzK41yl7IzUMHcZuTDdRyrdJ0zxX3EbkgeTmo1bp6r8LQzv0q613m3svhGRYD
uqHQTLWwuT9stC5SVZyGLtT2JCiNCWg9miNaQQR0GKl7GFMCT7bhXoAVktLa5bu1GExAac2VNTKv
7eAaQBDH3zAjHqDT4KbSW193Kf2mAR43kTmiP5sfiWTV4+BCb8qFzmoDkveas0V+mi8Gm4vqG5D/
QIWyIJMvtG8G2gIKdQzi+Ig6boNIxWGOMX7IRgweivOvn65cbxonx4yZYtpAXm543V0KpsaPrCsw
OrMsfeJ1jg1otFSW/YKxg19WCq430eiaxv+/Vxs8j3YPri1fD833XfFiO8iOxjgDwwgPw50DKXQv
/JVNwEyn22WbtoieiGhd1mIrr030ctno0x3WnXKTpVsNZ3QEuDD6Ee018sWv5boYg1xoI1X+hPtX
jD7L6/esmtJtgpheunJgic6ZXFaRIISD63rEqhYH6sNjf/3L23NpqQRUh/oXuQfqhzy0PHob/Dx6
zUNfthOuq1Nv3hQSmQEfVLLeKI3lu3TPMWJqI2m3abtMbPEz4VSHlQLq9KTCItAchuVz64B8plRy
RbAKooL8h7YDK0Cgp9jt64HADuy+B6Ov9iV2FjTMQ2OCpGqh/5l2NhMW4Q5u8z+6QaOTWSWkIMC+
mjJeKmUlIyCSjrOGWG9GD7O55DQdx3hFSqjGSldG7VLWAGNvi7FocfqViYsGTdBCyLIEWjdK8Bc0
Lq9IxBKyhzRiMlFr0WJhaCebWoru2X31ayP0fGbAEDjxZnUtSz/FbBweKiSzl83FeqFpneaTi+78
CqITuKmPk7HWhWIlN6FwAshL6DWlwNog99VB/Y1EaPxCRf30QNaJN8qjzvqjQsLRS4+ntml/sLNl
wqnas3SXNc38LNOkjpcOVMuG3chgsjMYwaTOwGfILE55yu7oalPUc+k72pPOtk6ETN/qpmtz3xat
L6877XarELxsurKX19bg8TMIxZmEuoO/lu6JgK3Hw9MwFKyszto8a/KGmoUou6m2U8cI0TCMpMJC
PdHxuy60y9aG50MFwpOlCmJNgNh5y58wWBQwAHtVShD55oK6fI5hMb4Fts8YKO5B4mnV8SzLbd37
XrfulLTUCkfwV5cM0Il5W+Nv+JbPxkJhy+fcXoZ9xLkqHlH7XLPdtsb1rDA7xAhMGY8W15ViQzuE
CUfYpiEvNiQ9eAvgma2iAt2WbAhgJFoxi/iiYc7bOZ8KPRe3TQ+ZFRWc3l0TaRJwVmKQSe5InfDV
oKAebNMVDIw4LHemDYlWPXIjG3EZBtQ2im8U8orGixtL+361JgIfiiK2Z5Ged+XScZhXbGrAVRE3
5VlSeJJU5Mskyaju0ycC69THnXEInJLZuEwN0kXOwtMfQJVBnZkAz+8j5WUI8f12UHQdxPEfbafZ
9OQSdq1OuPi+P0emW+JUXoU5c1mhkU0nxmr/EtFGm0jfl1C0ZS6gYHzsoGEyFfObaMoCK4HCrrP8
LvJMgGNtPGmRpUOEKWy87Wwar6dBrQLj/ux7wa6Lflvtpd4JS9bZ2mqAy9/RSRd51s52Iga0cZD4
+4Rut81gSWg9YLB1h3UVIBVZw0zvgVCC9/Mxim8mm7+4kfcSsUXF/lPEQFCMF1LGMXcYSnduaSI9
eXe5SZvBrwd4/HVoHV4U+DqfTfj2yfqwYc6uqX8bm5htca/cmzHL8gJTPr4TlRLLcKM1Eb7tqevZ
R0wogO9IUouM+DPznaazkVSqMB557SVOfv6uj+rLI2OS04lS5AAQUWNzIpT0EtLJq2/az8je2qVO
SMzyhRLfmIXe6LqBiydi0nsUSt8JUpICwx/vpn2Q6aIWh+0h/UVIUs0psUamwwq2HTj/GTO59o+w
hR4+qKdOof3i/Kjl8K1OrRfiVSCMKDrHe2OKcYc5Dw5iTxmN+xqB+7i0P4u4I4Umxk2scnuxvBg+
d0ZJeONSxSDgD8KjizpXJsyeVkQjKlFOW9i05/KogbRHpaydVqYplGqlvSw+CZO6gwTDPE1gnuGI
EVequkWjXBkwN8/WnE1nBVyHHymJ4XQjKtnNOsK5XDM80HwA+7UmZRi7TYRucB+ZMOXttqiSYaBF
oH4KdvsLO3GVaXxWmjN1PNoQ0QgNKphTwK/3+zY8VTDvsaYycDfUlo2OAr6WDkNivKyOl/i1DIcy
SrfZK2D8Y2jVOL9EvqEuu8NIYE3QTGbb+gGEMtcMC+bELqMykJIdfwptWLWoBVoOK+DHyLCdiO/U
QLDnKDgyrokXDqCAPzs3+TBYEdVf1w3UF+D94yenUa2uHY88vytaWqC5JV9t/Ty47ok0aYyEvKzc
HaQ9mXHOPBjx6MDjtXB/Zd7A6DPy40XNUK6FJAPfYcVgRNBSGzQR36q/LSyKX8dUuwlbhWKmn3Px
PD16XINTrDS4c6yQRROnCTwEVb9eFE4cO/88zuUcMpvQSZjKdGB3RH0C5eQlBRCuLicACWidGDhs
SRmjvd/gJ6tNdRdOhNNcufe0Zu6RBJ295q5t5GmH1QnV6uavvW+fVGpgEWggYcwhRDY+V2jUEwSI
mvanvtm5lsKBhUAkIpxsrksI8PaZgxf7iRmVN9WVoAlDs9bjtwn5KtLp1tWFeSiP0N2P8VFwo5mX
JNRg8Hbuez4IJelKpSFW9UldN08PuhXS7ZsUMgke60vfiXXCGoIlAMsXRum36OqQwT+vmApn4MeO
0vXeeQjEn+jP/LpeckK5ttPb+IsYAtbHQIwThIdH0xn+ENncS+Mk1X9ZnSo59n14W7tt9/gUvEYt
s18weAKwBIQBAqYc/zcAq1EAfhDPLEA0SGtDTqx8SeMfNmYuZ/q4TWjQCCalDGE34aNREag+V7cU
IJ3Bb2Xd6Qd2qAyry+rb3Yz2KAWezm8Vp2zKLOlxAps7EnFsObNze2MqXAdRbknIsOaFUpk7Q5O+
Nzk7E2fzS6puB53XvpDQ4xrvbMnmfaoijrLq5obmbePFZjrYQs0fjZ/47STNgcxRcABK8Opevvrg
lS6oRN4+hXFZWgjRcSMDMULmGMvoZadwa2/35eCAg9X06yI45IjRzem6mgnCzQsL8sNJ2cLsu9jP
87kljhZND0iAUiqJMPk/edO5op5LanDQ6WAYvK+2dpHMBtcP+oDBV52wy3bNEm5k6ELGFLrzeRvS
O0HO1RPwsl/v2lNvXUO9ekLbrQCSCq/ZexkwYRZpcNN1Qc80NsrzcHyvHm1LoGVUI34NQbgT7Ip5
lw+bzczjWTTouLUHZmFWWpTXO0MoEBhkC6zUvVxyFASlC891l07q+Y4P+zSd3lLmg6tUFjR0y7kb
5thLCgK51msNQfLt06eXkTk+mB2rX4A7rAucqiyNem2g4FbrtG/3/X7n3MqJXBoqd/ACtEi1fY/B
90U8q3wkC/o3xrSsBydQPxJC3NPy9gtujvu6OEsXEC09Z0qCtF715BLk5Uldi593FfvC8yLMWSwR
37tbJUD1vb/qBAroEYofjayMdv3v+SgAgoeCu4Nkvtl2jlodFgaeXKFXcQCp5DlYiOLqZ7sY6WF9
HxKHUBzruCVepqdC7L8i6xElc/bFoGavqLJFolhTkLirud6yZVIVT7t1Y43SQTMfbElPTU5zfoCZ
HSxa4jW/BtgU+bjEzSw+nQm9NH8d6gTHbmAVNdRk7k4znqwW3BAEY2yoJySYpebmzqzRGT6VxtVr
LMZZSsa2aNVwWAfT2a2yiMRMZH70fExZ22vcDAS252MkbSmJXeKaj4Xg+IvygoHfB9jp3asvNvgL
gNuP6K8CQl5PxBzXNTpQ9OrBQPerSXe8AcXyvrfeWVgR5e8ftRQ9N4iPruMuM7oKKgOtkpvBaWAG
GE+F+CjJ2vL//KXnIUzHyCF1o5ZZD/3TEGN5BGij+gLlt7424aCPz2s6hKmflBWIZnN92pWO3r3y
LCu1qT9iCiLaFiEzNPatZJxZiLZltBy2JxPblZ0QM20Eh0ZStGk0d/+lLQduvR1Gyd+aF6uDUpEv
xaJY6xarT3/Ucb8Zehubyq7/WZ7izKFNUYHfJmND+ya4uPjVVRJrUquPADZIflX4q3hwZQSDVQtZ
gU9T9kkiRNMKVhRYcq9Ui+JmxUPK/6Og1/ndJSVbENWfFmKPyrxh6x/K1REOQ9GlIhInl3fR0bJq
IwADvwM6qjIrLayvvTNGiN8bTcTN1vY/xCJkaqGaVvL6h1BmBdFEsm43JgiODz0JnmjO04dLEXmB
8w1LdiUJTKUjvt+lYMdNvYs+jKC4+1tCGvtNYOjHzVfvn0Qjh5zaA4p5tn1eioD4qdwtefttMyjd
xnuJIN8MPGBqxSpkZpIeaPXn5okBG0LQELq5ZY78XhSyT87kAbET1vGGkpO4XbhXPSuyAqBxIvz4
wumvvUiVBUOji5AgHnmieXh9ddAnX98YhqRlXlr8l58/ZS1u/m0qwryXQX0YuWxtHc76mbN8a4ST
SZmp83b41UpZfrhSP+YGlJb2xGXGC4gRFEU43WwFSlcPIrcW2MpC0437dd/nBMED5qoCy2McgpCC
zRuajA3NC3ZLkrvvZSANF5Bp9sJOhG8pO1RVl3gHMxEoOVn5rv4XCnmofrNDMdtrFh46Q21KJbFg
7K6yFihTP2x8g/shx8Aki8aM/6Q3yu/rebnFedbLaz3/y78vDCqE3wrFFfPq8d1JJpgp93IK4Iqf
dHDtRNzVYzbhVTki4LCcgVXaVtMFeKXIt5AW40gvxn6IHBd6KwUCWsy73EQssnDNdnf4tA9zpAEL
9CDMPhijOOhFQts8gejMn3wHQ4XItvqSEAH7sfjbKo9OJio5TvsMskHcWQYF5fBFETUD3cO9OO6B
CdHdBdSCtnxS3nHx2HzsdxgpN/PLh8+3ldaAQqA9hTeFmxzaNdRLKPbJbH+35a2jeYf4NUNezsgz
XaE4KU4dsNM6i3OgVipPzVWS5ErgW5mu6v+p4POq50M5jlIGAcQqPD8wrTgbU4XaMfNQIQ3gOThr
HYuhc7FN36OKW1nuuWQlHnLUj5nC424gBni2A+jsoJevu2DaO+auRfxuOY4NV9IOsnpqQrHZg7d2
GrSUz+oKHS6lvPqhRWnlhUCOEt6AeYnsEiSAWfT2CuasMrgvcSwuGvXLxCHuyNE8VnkK8/j2bmDj
6+qFBiOPBesIDFHjbSPApioYHcT6PwxOpiOCXYqpv+PYwYjhJ8XpUHtw4TTA3ZeG67qhd8HW4neC
RXUa1tTpn1t0s6Nbh6AcC2JPg6mVys5aYAfLLAprNalhygwQzEbbfWW+kYfF2/tHXYEhULQm+STd
70US0q/O9STgGYmdi94wjR4dj809qTR0e5g+acKXNE1ATAAfQkAyB6kWqC075vbubr/021XRY6n2
V/2V7FN8SGGkiSoMwCOg4dfLkre+SLPa5GQcWdilvwXsTxpDhjZU9k7XKax6kpgVhBw+SvaLJ88b
48Ihcgc8HnkHMN5zuYQ29aVYzoTUUMmYKT98FVxQOW5a4J4rj09vxwOuqu4kUo7rEFq5RbOzoQ6e
70Z1yNA9NuPEPEH6+Wd4anMYMo8gtsgELH71AZB2uSmbRin+E3ysxm+xX/OO6Q9Ejz+o6WyBDti6
ip7jxIm5HsDZ2VFb/+k34l1KSwNm/OAhzgzYXPwQs6qViGTM9GhOf7ryI1QqbQPJIANFVVkM/IV4
uUFWq/Wj2PyHDSSSeMim4NYdtqE1k1O/0sXoODQW2kuIWsEeR5PVAFpbRERFsHi15/x/a+G0bpZ2
z41Ynr684jhAjx7L3aTlqMEZdZ9/HPRAS7x1tTWADdesamA+qUkwkVK9RuR2WsIC8UWg5mvFViDG
Ejo05KkLoGhFC/RR6OZZC2WY8xxL5aXio7KjwemxhfT32w3qGJN8fC9IZeUBJXd1ci/J32DlXcKr
RUqY8czLiz9BHg61iyrNkixIvm1quD/wazWXblB/L6tLtWCPctbw5Rxi4q71RTAcJK6GL0WOjRHa
U4Q4OgwlSqBzDxd+u2Tpk5ILdSy3LCcNToLJTAEk0U2AE9L2soN/Grig0dPYICZvyc+J9CBBG1Zg
x5/wwfQE04wfs4IgGfZWlUXWwI6FHgtftwOrnRQmwM6EDgFFVHcCxlkIN2TRiPT1d4eA4F18bqkw
nkx9zD5KjBZQyjNn8+fSbbg+BOapDl/f9KyN/5cq9b5e7DtobHyDShiuqL3ta4V93UXIy+srs4Hz
t6jObD2wKJ2KZs+Kq7Ukv4ZLWhcpvGJmeANvEPcpY1QqoNPMnn0U506IFts0wMIqCg6kLZz9EH+S
nCvIFIBbwj0nZgzdoSrdH6LksNXSSvEBppQrkR1qNfXFGCRkvCXrfASWny6wSwUCUnYFsj5/Df6X
V6zzMBdWL3PTzpb1XUpUy8O6maFNC9dRGo5PsV0eSnEDGHj6miAYRxKojSJ5mbhYKTXPhEbnpIKd
scb1Sg8pfJTlkbZUzC8digwSTGTGtrtJ+MTCFzhEHkoS1ZC2+FIOSdMU/3t0HUuPDBl+CQe3b2K1
LEzUHCk1gXl8r7J9366V2y1iB1yjLomxxRAFpmIYi1I2O14aXwoLZN31kBFpAf6VIslzsvTLWA46
H9HLREmBLTxuYLT3VNyVLzwzvsLOyxKrwzwdiAQc0vzTsGmFHwim78FgQlH7NBaOx7XLQPOd96qk
LwvsRcBa4STLBK5UqEv+Y9UZ/9e8eMvByL6BWHYhgGS40awGg2HrG8ZdPK0wG5lZ4lBT01GUXfNH
N0tejVuiOH4MCL8ZxRD4WcVbC6m1uIktDFfXmoGdagR5E+jZWEb1RmiWq73MrH46QSOLPbgy8XPM
pKDpjz6sAUtKfn0xMF8l8VTxuF9GIKUd1k8HbqyHJp+Uw1sYQDS2wtIi7manyiN6FIWgARl9D87z
DD1RB6qWEOQZwh6MjfloeYZ76C414Mzrhxjqjhe3gmTWJ+TM4lnZ8qqmVXzVRf6vL/rh3zYdrxDz
4DWOlf6ThxsY1ij898yuQZTLcaMgVkjC9CK9h4ztiTqf5uqo53oRVGWd6EYn3M3yQ0/BXMqInn2A
P9Nf86WqeIxQQLOdb5+rUNW6KhvKCQC7qzx02guBg0oHUJ5/JogHRdF8zv0HAVHTGE4kI0r8ylaT
umRy2cGpxylOmT+LVwS1odFW4wyZqukAjEF6UiOlh1jAtB337vdqtTRTl5xJT1BNIjnt2JmmRnMf
z6MQqR3f1fKUVnE0w+Kcf6Ya+JQIPAFC1/PoZBKPWISjD1aEh/LiKqVNA+pvfP/IyxSGwFRRSlT3
WKuSDaY877MdFNOVdqvkV0EDp5A593IuDLYXm8iRKgLwIm3tHrfg4rr4gR3uXmF4xJnOKr/weuSg
DwHvCvEXCQykIpVzRZRMzJzabPSYgTwn7uzbzLsMTsyMwUtT00qJ1NmAccvw25ldoTZOv2onYBCX
EzZvFtxY1jrRrmlu8Xp6miSaHmZ4lbKv8KEgkR0q7jjD2Hb1hzMBjcUaBIXtAj0iVM7iAAnlocgl
ziPABkrlPFix5Ti2xBJdNACY3DkmBG95PaAHgw4JPhfT2bbfIxpPx7UCMd6pEnO6SMLYJc4CI+Lg
1VFDa3KE52gTIPIpmqFhYqlccXCTQy50Q1qOSCS4kAU+CXDQDvOQKbYxd9Uo2CL98OXj1lXKwsr5
vO7zeg5F4qFHa7zdFDoeSSO4irOY0ig2xmVdT4ZW5u/2d/Lq7BwM2NWFOsbfLC3HsxOQaSTjaPMe
JbHgDN4vYSBld3wbRqGSYNlUXXyli6Z/pXY0DyKBH6bP7Bu6G9ZC0QXary9JYNfkxIXTL1xRknXc
Q0sWTOWoEOJNKO8qVNwXbvZDHLrYt172pYGbZxqCx/RM0W/M7VUkmeMXqeR/YkLRV5Q9d7kEnEai
BLoBshCHJcrDg5w8eWxEpgCgZw7eNeVadHZNJiOW4q/Mk1WR928k/GxsN5mmypaTc6Het/lRMXxj
OqHVB9hCqj/KXj2Hwn0ysp2KTLDKcaVrjbzvtQVng/xN1FOMUhGZJPas2E+F9s6XeTag1/xGXkRo
VhtwTSs4ZYq7VGOpjH04zbUeVe7thspteRgf0TSwKmgXn+73Qe0cAoy87d5BPVh6KXs7DPPB4lU7
mxyxr6yFfYkY2OkYk8yvdlaP0+Co4Jmi1WlHjd+7wkT06gKGQz84oCM4bwKxZSUN9voqkeWQ5OX9
mH6+N+W6YH2cR6seF4a4NcI+t54zogUvyP1bOoR0w0viiODCB12jhgOSYi/HCbwNSuxkDYQw6atM
nq0qTvWMtnpj/AHeuyrJL5TED/qmIJpEArB5U7o5xfNNl7C5hhABwR1JTmHz2xIB8n4uaOab/lBP
DmkhLIw3DV9i99c8wjNZNY5AWNaas8BwQtyOh3ysIkXAXjPiqUgfqtg7UCwU051XuNIVFMe5v9AZ
a7tgAGgdaXC6g3PJf5knjlDVVYbRmG9213rrnKihLb6cuHT00kdXfoCaYKvoQwwoLOhusY7pIjzc
h4cOC2oNTuIMMiyC7bj28a3CAHcSj2APkSNaGHk1xlPBICFCep4gc0wLeyOmiUTi43Mx1AB242zc
JTQxm/RrfZzO0Bpq4zRxKi1ggTCJ7XRisboJhQ1Gny7W9zvl9UBS49Y3xKM5wNYbF5XQdhwfOjH/
v0s0S7O6pq8XhqO3+jRAHxI70qHJj1/OgxQ9ngbcxUH+kvo7kldHfT7KfwiM+f6UOGFs+ci4XMEl
PxkqkoGna4T3xYzpokjbjyRop3r6hZ+4LqBSjhXNPv296y3kAKIPvA5ubTKlXbQBVUZDLvxYFwgi
n2QtxxjfQCjfEf/zXJAlehfORwVCVTMsZEmId6CeoIdMoDyrZRYvQdJnynf3OcT7M6zoVYhPERbI
m5EHSe4Li99WM+EIKSbIl/wRCTwmt/p8hE4rBXEuq6Mw0exXuoeLUeKxwjn7AZHnzNjshHrp2Q4o
hoW89sxtpKQs5M3D9I44fOfA58T16n+iWC0si91MgXk/SLADfygBjALrpbix4p0ux/fbHb3ApiPv
lvyx3DpTsvHJWHX0z0SQk5szcZvzE4KmrDiihkwopWdQ0AJ4WC/f+NPguOoKsCLs/cf1XMpuSJtX
Q1H8gznDHCPsq8NCZN0RkQ8aV2auTUzPDG6NFcq0wc8GrsMbCTLQ+4w4/4DlG9EVr8EGpd/dDCoJ
vzfcxEyl6xPL5SBeDFk4jQiER54kEfTBuKSyscdTBh18KMffgbg6RORGDjeCKATuRUjgbaYUiWjC
WwrV5N/UrqMcPgvwv5vdznNUsM5b08QN0CADUW2LVw+xKn2ZeC8d6vx3rtjkL3rOvSTdbZbgl3/Z
8+9aq+4VCWvGPVVPwDCietXsFzCmCDJHhd++So6ct4LjMW9l6DECJtJV2CQG5h2Y+LJfeP3ACoyc
j2EtR3asQcefEDuYm4E6W/KIqjBKQfcDKfWFuQNaOa1w5+07cH30UIdUPcFZpEB1qfaZ3vNUoJX+
UqMkTS92Y3LjYiXGROQEEs0L0GPof5QUiZEIYRfU2yEs4xsZIRhlo11jfAD39wZfIvbkOQbYPH/u
yKvE7m/YOQzyyxpwUNaUUoFMF8QMmDtG0vrkd4aXLmPB6LXKl/OSMXT9yvITx3sodBoS8xR2rals
WjeNYVF2VDjZZWUaK2fwFxBbqWbd7A4xhZ2SpC0FCIeyp0dXy45TE3B4aVUnaHxZOBC5GsuR5ot9
3cyc6jZVA0jZYnX+3v7s86y6MbcaV14OsQEKUbUCDAKNHSLvKreq3ONnjZe3qO212fe91aJ2rFE0
U+O4kkc8Dbm9Ltfewrje6UB9Ko0ggzEJLA16Fbk5xMryzevcMTKmfbLOXTkfGFstW2fTAFNdmu/C
c7FmTrATLDsIRE+p5B2yYEWWubyIi+E5o8d7YGvFpGqPjRHPmTQqhCBxyoI5hburzRUhtd3Kj/f8
CNm5EjTNrRvfnX9NeLJB96T1AOMqzW0CQA9C4TBZI+kM33d7gkt7NfNXLh09m4wQTzSK8Ek31ZdX
X4jCwY8y3bXJ5EIBVHEhbAaWLYVo9Ms+UNAkmuhwTOWI7cYhikdzE79A/Xg/ODvxvewjtbsZRen/
WaTfuJTCs4UZ16S6X3viOFxapnqtgh967fiNhcPpy3j6HeDy5PKzumvcHISXl3K7MRSj61zDwv4b
SjlO1AYGSHhsQHrPh25YVbUiAgeoISpzLGRFDSRWahplw9J8dJ8gtMMIax6P83s9oSn+Cx866Mdq
OjC3k5ntVOrmWRS+9lUOqtVjd9R5D/1TBonYCVDvDBycusL/VrGDJ1Cmj/LZhLuwsYrKuj4+zn6i
fjjCxjDqe0npJhfI7kMUEbbVbTBUJLMwzhVyhadGzLKGpsy+kkmrTnNRuXla65H0nruRYaklnUzl
7+rwB+U1PI2R9ptRvxd3lSzuyeekQiHUjGCgL3igRGxzBeityiYCXbRox0zhk4nnCvcgQNDYfT4r
HiKjl1WXo+V3WoTi0ycuRKMqvoAdkYGbLL1coE3r1tL26dutuj9B+U/9hdFMUXsB3EZ5j8AUpGVi
SWtjX5LFmmjeex3dds3jL03sE4uwz6CqdUPgmGP62Z5xUUVHWhIIjCe9PPWSitcvuJ3p1vbhXCCH
uuF0AvIXgiRxiTBZJa1hUH17n7h5NFbxYhi5TJTY2gSCmg7jHC0UADA3c6FqainH3w/CsSekbN9B
vod/xLHHjt62dzYGBwdHjllf73hj1RaqbYkt+wufVSIWlu7q5KD0t/rRdafJDCxLrhCi28L/2QO8
93h5ziLsRHo6Vex7w7eFOLf+swyVEIST8ktgzf9a0dWW+mZ0mKK3Cbijd+ZftgHUOZDpof4/tg6L
zVOBGOK/fTyNDs5KTgOQy0wm2Wd9jgHGVwToVr/mGPqf7wPLDNjAzKett/KzB18enWl0WpYiQGw1
mbBZTji6NZkbm5cE9+HNWpXPIT5nmP8esyPrXC5/zgaZCwkRfpq3maQvtA3iPXT/6CdSbCFEXkW0
jgZUHhkkoY46mugHLwzMzvcPmvVE6y48pzQ7WQrxXamtkrL7DjR8u2SKKT1n4iLQB5PWu19eaCA+
Xpoa3/4ZYtzjtvn+V/jXBnu2G4Ch9Wua71OV68NBZ90BlM8yEaVoJtZuZxLr4f0Tn1G85nhNqyJe
N6DYy+IRPg6xM2LiQ0kdk6Vi7nij5S6rn8ot0hXs2PgWiVYK9fn+IOwBy+lpl79r/rnfmmbOWd3A
ZpO71GS+bssoBx09zW9QNeSBADhLuUfm0GfHJpuo/p0jzwBS5+0KcMuk7ayVjSQwshr97tTfHgi3
Bw0Ah/ZKjTy+gqxOFouHsnk/bPvJI18IpcpSJtR0jBdfl59Cz708LicqsU11KLXlYfIR/1m09hdl
kJgZ9rXn7lEF+P6oGMftnIflNbfJD1INW7PMBXo1lqSwl72VpqklHqMQbV3CsZPSDX8/5viOC7he
15SF2zT8UmmXxBzYYCTlBQOQ9pSYUtCMtuVL5qCRfo47zabeGQqKA/A7YrgI4tBWMDS4OR5KXa9l
rUbCFhSNW/twvRHKkD0URQRvEt3bBTr+brREL0n5s5Z0hvD6q4AV3jUV048NMWSzxxhuDn1V3Jty
treIjSFmBsRPkuGwVipYR9kx4eMzRPQ75kSLEv4HpVhKp44Xo4kM19nnZO/vQm36dGlRbtfExq9r
e3b9qXqUCjjmcfYGGgY0eyVFRbMyjIODjCJXtv5UBd+ANZt3fUKZkG1W7Mgvti7kWrr86ueUTCoo
TDmdAnkFU1DCqsxghs9k1aNdb/jqxdnkYReZW9FsB3grDvk3yzzWLLuXNiPfKntfx6CcNSClkIKC
qImYFIDHVocb8Ab7wqTS35s9CJPhcvS4vpST5iriSDJc+/LlHzUwZ0t6x3xoXctzNx1gbzcnttQz
LIAefzhU4Z+79JchEUgN66DeUJ9oujsdjOwKwIMyZEtTzkcxvktZWNXKllkmKI3HLfquOdvgHtM3
6wBx+SAM8sOfFpkcGEPXjX9VhgEH6EchLGpSpg9JoEWTF9OOSOED+ZWoMBbPZRrDA6v2T89ZOObK
VkrIZrx061aV/ZXe2GteRk8AUs3ShF/ee4oZWk1oqzCvIG7ZoYlXAWVSBufiIp6OGn+8obzv0FcX
0KSbwQsOcWdwmjMD/CWROaZX7k9Q70Q6FfsQx7EWbPLVv6fkATRDgr/pkPPsoVGGZID7ylPyIW4s
bkf99vnK4viBmGIdQ4/6MDaRhgbrgmX3eIMMyctgyoPICqA6mSbgC4JCzTZIUUad+iAqIIxy7aRS
LLZUdz9kzxWhXM6uDqQGJo9vccrENrg9aaIIjMxbrgLbh9fX5/NtKuF0tuaDhKnKw/46Bv04iWn/
cL7MirrUZKJ75erGANk+QMmqMphVuYhzk7PnW98OELQXNnyLn/YtAvl7lvB9iM10+au6SS1fMDNi
U5W2e3dVLdWwrVbAMyECCdwRI7mrWvfyL4aVLA+UW7sLhdsLp3c8p+nWhO5TOeyyDdvp0nNS3stj
EOFbT4rtTPqXUrpugZJTyZNTdd/rX8shW6vwa1z0iBOeOWY2nSHkxovi/xcLgZgm+JFO4X3XoCof
QR8U8ujhRGTB1i8JTBaT3Rz7hrgpFUjgvLFjuwUe2LyIv+Ywv2Xqo+cgD9qNxCGzw9u7colYAeW9
k184BpKWYnqbHSXyoQghLr0EXuB+95/i07ulc46ac7o2FJQL9nN8XF0n37R/mqPwYeAXfnKjcP75
YU7Q69iszusMDYWShf56VvlgwiX7M0gYRFlnp/Q7zBD/wXVb7uFPVLNDLZu31CUpOC+GUMuaf4s7
6vTzKif371voJkFHr8Bz24+3B9dl80tvfrBan78QX1s3l++h6aYfRcEj2EKtcRkpWgrFa+o4F1V7
HHqgXV7XzyHahAMoaNGpRbsRbQnE47pkQZXhF1VSZZEjAQGKX5hq9AwFrX/jqv3fhQuOn+5Zhmql
ZZYViZmrcFmhnskTxSqORW5Q9+HpLbR4Odw55t1VpZRb2CIAISU6A8ewTq8MO3vTDHxqpkn4ks0w
SEevp4ZUbr0IrZ14M2Dj0A/fz4JLtycH4AZPAyqdDPdVV5GEEnNkZhtdWRXvLkZIo4frjwPajPs4
gjNbBqqhIiY651ttQ1WSNOz1izD+ZULWy717da3Ae5cHBaM3sXO46csaNwUn5rQgVK9yMyw08D+J
MdK1VBJPDCWK6mks6MB+DB5yC6RTxVKdP6gODlklX35GPq6lZe4gxFqOlUIaGH9sdWUUx1oveuli
3G0RLU9fQ/Ch0oLU/axLfkzf1O7xF4SXRo5LxvSJRk1BDJVRO8R/x5pXo4Aq1ImkaXDZEn+aEomp
eXook+Yp1iuTXv6NTBrMcm71rpfdt5w/GX4f4n4YeNP6q4XWLGcer7jf3ZLKR2Ddx7RAWAvY4znQ
tQ7uGxjBneL1H2fYPYGOpgxWp1AQrNuwLVC8xKggN6WxdhX1JrxUZvD5c3Yvumb1be2j6kP4A9MP
D8FBX+l1G7l7KFRo/pCEBge/KV616+N4mQypZnvzyTcmijs0TdxuskMBqFUjP/7JUxT/rO7MkDwj
K2UqQmz7GBskr94fRwIAmwvT/N952w6UjuW2+QF3xEO3OmF2wPAc8uTX+BXke6yj/8MzuwR6TXm4
Ob3He9+HruCEnuTTCJTqGuESmm70EkkBDJNW0LGYThn1pojA+QC2QNx41BOnjmHsUGh0EQAL1nHJ
b/8b6IuEmAOiH5iOHKyLu3VO7sIvHz9xG0vlWooINVgKzAmt8/+Og1UEBrjQxsO7yn6yuvFJhUwA
3ObynNd5kMz2eevljYvCi5xYXV143QmfLgF+AEcOTcgbJ/BFRY028dX98QyIpbBKgjX5wNFF0rL0
ixB9k3nj87hesR5Tdqexlb94PVxC0NPRna4jreMj9hW57NZSJUbQBPCCN33ad0zlP+LB3/3YdfVg
LONl49Gds9+gT47ezt26jVxOIQfRt4IIIq0V6by1APIPFaLo4cHkpy7qkPoPMcdY4dXoxD0vsJsK
+aBDEzp+DK+ba2Z4OhcZaGDl3OL88Ts23redX1cTmybgYcwEhtc2vFGKhJnyPxE+qXEELLq8/CWI
2C+ozWgSGlmhlhLGExZKGGntTQUtAH5+5VEnH/SeDeZ4ij59sxV34V0nTAoYNmxyJ7N2vbIijchN
or144U4mH+18PLwJc/r1GPTVyIvZqeSJUIdgoQunSpb+bftttpoZsurL4yj7/Hv665NjSwv/tVuu
zdTEEUdaYRCRSLn+1zmClZJ6Pjf7U18ZysG1GT4Kv/MOBerI0VBrm6/rSRJyJGx4j6ujPo9BZdE9
jOHA/7S/P7Qr9498No3tLNbSBqCqOLGObjJNpOuQDYhaYBY8onulH7pPB3wG/LTJrLXxRbTSYn0Q
wwF98nGviWohgPoVO8N3nzeRcVWWO1vuSYBRfLmwwZVxiJQ+GYFPlCN3R016FjXTB3rIFnLv03RA
crWaTWIwvFqAAVJunw1Vnwpyak0uDr6YxZFiFpxtKVOU0WBImInRBW8Abm8eyfwsdabXOjFI2yco
iEmKy2oTGjuEroRhnvTYhCDzVUnupJe+q/qldsKnz0foys+ea4tiHjcoxpKYajmDTCya7Q6NNeXd
SSSowdJwiqybLT8EE6PlbsM8gHjQ9ZIotenhzQTjuldM+uIDjcvY2/Z0TMedjxvCWzE+opYkgQtt
ENTgQVDYtFbYCIWfWCKqqat4YNtQ6JAOcMcZs5225RqA25hr4oQ0tdYsVPcAvhdDYqSFPWmUlBfi
5dwugHfrsPjI50wiL53vkaKA9wqaZVI35UPMRIbIR9ieoAVtp3WYhKdsZxrgb3M1rcr3nAAMmpRs
+H+hJiUI/5nS0T+gaMHQzV0M9pJjJ8vRzz0uDlXGqL9iko5BCK3WmHLoyVV+14p4PSn0sqk/bkIe
f2s/3ukKL4E/FlzsJTJHys3IwalWecdAcJU7393uOOtICbHZ+u6OxJMMeuNUXV6hfZSZO/jSumDE
ogtS8fVbj8FeAjyGWO+gbPkyp7fSzmrKa97gCXE7ZyiU4ZjJBSRBIegu7hT6OWMoN3C+WcHWsNM/
D1OHd+/g51F0Z8/DEA7KKWop2sHxPNPpkjqzV3WQzrWhdwnYDKP5oqxhgvd8aZOXnfYVUG9UbjhD
QTEkA3u4+5BnRZ62BNC+YaafUBg5unjTmvTJcx7JC5kHgRIMTnbB64W4tAgeox9nM33Uagr1xhcC
nwLjtjFW3CkkqXuoF14RNAnqp0YmD4Ge+JkTlP8jTTow1jsWT38clXHCEyS1DHhuHmuODG3N0LV7
jLNoc16hSZ8EIpc0b2TjFOz3lex1TOKFxDeE1vyPk1oVcrkcH41EFLdYcfS/7Gd1AgAzXFR5GQrJ
yBJOSkiEindLb5gBy5+ccAxi86u5eVwEwfB0apEXySrvsbiwH6qEhMWd9dsF2xRny5bFSVpoC5VU
pEBL/2wZ13VxCpDpDCGFPmKPk83bX5OpHA4j7XSZR++Evq0eCVq9KzOXYhSk4ARPYZ5400svz1i6
ytyUtjES2JLBoLl/q/8W1/N3zuMGg6Mnw6YoT25R53IhjK3KmgAMd9Tq8ZCBimolComuomIewFCh
2jdbALb8AdwaAAa1Zw5pF2wb0FPddQHT6gYg+ATB8m3a4y0q3c6v/qo4IyHwWmS7Dmua42yEmYld
jcPhHK790jnuhNxn6i1Kbr/2MaPBqnaw/+PIg3Ro821l81SQd/Q8eKJpy2aICgXfxqQyySt6hKRk
h/daZj5z06ZZrDqN2xwLnWMxIQBy32JEix6wOCPlQa1UEHPYdQkcGeheYPcJLrTyGrmfftFW+ZJk
qg+0HWcIiXeMvokObE1Xs8h3ZreYVDAE3fZ2oDs9u7tEwD8kiyygNZU9GjqKWCBEs4w3tGR9oAcr
NqecndveAVC36ggOVDrtk1tbZGB9UrO2t5m17TKv3FEBfmav/Hq6NJVJnQXhZBROStbh2EMWtf5H
+9xKQieck5gDmbW5JC37/VmcKumhlGuOPF2aqxCWXwXhvTMabWpWGtONBXJDNGNS0nI+lJz35n9Y
JBkVXyl/J2584lFtln7xC9X/A7cVV/h1PZA7SwXD+cH8Bp7uZVOg50LT58DQq0CLgoKFDd7HHnK+
P39CdNVZiG9YcLs4v21veIQgGELi0wy5pMmRyMLV5cOupNM57fuDr2cnIBW+dyISaRECpmgKFh7V
FrYvPmwtzu5zhfr6gUlJddffRquAWfG/omT4Ai6cAloMI8effPkXxpm3VQ7BLY/QFoT/RL/keC5V
EscNGe/14Qgqg+xntUN+MyA5yjQa6FqQvLRaDa+GabL25QRWc/Tpq+CCVA+BF0L8hqj0Vz5JRaJs
Mxm5wr3japnP0tZbbkFcvjXs3JoYSGvFKYS2usrSfVZ9hPfk18+gNCYKGtwVMdGNbrLFTJV4837o
FrC320YS6qHP5CjCaZJ/ykkhiUhU3xuWPoVEpHfkGvG62M1T8SiNW5GVGSNNSuSZaDPXrnv0peCg
WNM1g8h44b2RQFzqt6t2jVOoP+cvA2HKpgbhWmKlrpXGsJR7+80UVP5r+EzZ2AWZJTAEXcyYlhiR
J4YDxzy93utNrA1DrwR5FnVpdvuKm64y15zG2pvt5Ep4XNVt7I6l+ir9BWTYgU86DvwYioLvrqbL
2Av7UStYSFUWRNIm5A+OTOQ1Ntgv7fI33MsBskic/SVa+XgWw0vtt7vStuQdTBglXyDhyuhE1F3e
JBoG99W81vXJNFV08PWWiGihJiz6h3oYNc5ery7nQGsCtfYWc0xOS2A/I76W7UUKawKVJoPyHzO/
BWMmWBp5RxTz4czge6cWrrkJf55xxNhw7BHH4Dz4H+0v85jgKg84AGSTh/Op2t9XFp+2ykKDsZgq
2iVCWFlPkYloU5Wb99EWSaX2KZLM1PsmRDMFVooupAUnBevKNM2QqkVRDZJFboiHYYZjX4ejTDwS
a4WaRl3BwlsS07w295uu0saI0pgKyPN6vO1MIEz1P2Lj4CyKr+EK80jVL2mKcind2YLGQIuscbIX
n/V7B3xMR97J0kgWJObA7LKW1NJvxIlDzvU2rUZkVfmWCl4ejzCzuw6OOX1/BZ5Xgc72P+WHwbTa
YgYDnmqMZU+el2JL1GOonOvoSls1IjqoX3CwZ3IzaQmGrHdHQtWtXNH9m2nOy+gbV979wxIUyK3t
qOmFZ3B94Wq7OYgr7IsYBTTIuHcIGb7H/993/qFOE3gnEm05xZ47hFT8YXPsnBydadaW1u2mJt0S
/PodWp6HC7lopB3hDr4AENlIXg/QPshV3ihKjFg0a13kyemixoE6WEIgL64dWcDgvcDf2kwzJVBj
BQymQCnfE02rpUrLoZaEwKKWSxqCbv3YAcK6yMYW9rNvnAVgr/l5q32wjFp/HHQ0YkJrAkt1ZS74
DYzB0WDDoxJ5JHZkRqld39HUlVRgPuB/yeoHTtlrKyv62SxnFI31ja8BgBXSOj7EZ/vmvb1h2JMN
o4F4PRBGDC1T6RHnNmfSGYT/KQ5mzBxqv0ilZsqMBY3sZZAzhHqgtVC7DtX/9VLm98nQhTYpshWP
rFdbmhnC1kzhjiHokdGONh6Mn05M64CenNLKMnDsdQGA6cnnWLNic+/eQ0tk2Z1dpHxhRdWMp6us
p2mKyYnev+Of8chxlk5M3beh3utZTjCPuIoUO5V19L5vPsdgsiDfEBIuCPALtmfOHuVLmptiHZH9
wP0MuFFFUAOPAPGQbPlNM8ET+OCCU1ezcjQgshFHP38Dnbfnd1VaqKNYolxZWArXv9KNsFRHg3mG
8pIJXo5DcpM5ptph6eK/wkVO4BIdShadnKsRRYy9F5lh0/0Ic5UOwPgmaoBn4BSEh9ULV77IblIB
PX0p9QGXi/Vaswe+ArRT9dSIuYpKBJCOjj5HzEdgoDDxe0JUFFU/c0KCuvD3LVD5GohDmkfhfuAK
mdUjqvPHsCH9DkiRdr+6xJN++M9kSeopuujA4ty1yERm5wWLW5ygSTBc+gsvYN9rOjkZysABEeAV
2rWAnH4S60XQYVekKWP7cKUaiI+UV41UitlBi3ciWUC6taeMRsJCyONRtnlro4+izllX0sGC2iHa
HbMECQHdYIHwhRUOKob212XfJiYbHPPmuA8L/UIR8uPp4xZeT8CJUmEzul6WfOBUU/SbVrVMRkyB
ewotEmV/h0BUWppDqGd5wYIaIVfrFl17uBH7vh3zedRS2Z3AK/90YJvw0LVS686zS/iNfYpq97Lo
BQvavSglZp9/LHkIXBmAQ6Ac1Mq/H30RU6S10DEVz9D9KfJkXlyWQ/AHnuVSaWopia0QvT98XW6f
HicLebomLB9fRO6xsKO0sGbiVOS6O91x4RWqoJ3kFOe3bVVsS4RI+PLlNLKUanvG69W1VOWyWTw6
4io2+QwtQ9FOnmx1nQtiLa4QEB3Sbq7amD6Oq2aQvq05DiKKUhXzyKRLSAauGycvrnBdb3wC1PVb
NvQ/ehYPCm2ucjvr0BDIHqk7AGf5H1A5xTnnvPSM3N0NctYLV6XtzvWcZhjGSH67FhCZ1fgl8uPm
S8nfw7P75TUx7/DphfhmFFltLxkLvj3liCf3I0VlBCapb/qlxOvm7GxiLZpp2Ukl1dPSadVBHSXJ
tVHMK0b9hiTQ7oGO9sexAPm5GWIe7EWFLty4ItgLUGjZppBuJpZgOkU+MXnQFQ7PTTQ99getbzjo
NoKocp/NqbUxDPsmqKqlAlYUeG05GEEvjTzZi0pl/wJxuyvHX4lbB2z/64KkJvqZVFVjhds/j0l1
i1yLpxW0+GGhDDipyh5AGggwjrM+GSp6hohmIU2zNDwb39QEQ5UPIrwSvoucRmLcJjKrfoPplObx
ej1AeSkY8Bsd371vz12SFECYQVw8TeNzN3qhLVBF+nibSoXu6CMWppti8aD1i1Q2G5bhJQa+DfJ3
2o7Ruo1cng8n7EW6LfBl8RrHb/zfUTiUdWMlzBfdmBqPfBQICaw0KFkNkM+fqNoE7Lk6Wpb3dVFA
2JX8RE81pmslCFodjdHEB2nJxiLYjNDmV46DRzG1HXDDCl3FoRR+Pa0bHr3gUdcsdzfycz/C15Ot
DbCe7WkvuNT/uCgCSXDXWHnf26wvsfqv097+IgkahCHhW/KiALmlfZGGSbReaR2n7Y2TTO+bea/k
e0aMSEoZY9zXYG8PPAUhuUU/TSPJHp41xHU5MWMXIiXG8aVe4+ZntsGveFA27qaD6J4V/rGI3atx
rE0HO//0iuW99jNwA8dWyzOo6nIuB//eV5W3hevX+sN3xGJXvPttgLsf2LON6ZqEBPC42sahIe3k
ekdxap0hRNm0AUEVUjpR4BOIRYOzTmmNND8aLZ3V132e9cLrn0Lwi7kFPy3FtFULbV5pjBWQZxUx
DsZqv2EXtaB/8J/6nsw6b3ArfYrHUagGX5G0khtwMBiehPeF/tDSjKiREnvrKVIahG728euEdQoo
9NKhgrm9znMk4q5mTaQaNh7hQ8TZjM/f4ETY5yNcbwv2w4fLnI/UdObS4QLj3pTzWt3o+6ZdzXLz
kpnkg8TNtrcktMp+t7aWksrI/ofW4TsVTl74Jx+Wb8RL7U2w0LlM3NGhmrZYjhtO3vnU/IMnUgVK
YCcIqNw/nQijx/4poELvghFGYCmG3Uqspr6OFqfoUQqXldrhorKRsABOwrpuLdmlavbvyw42FpDb
tXq1uV1JvnCeFJC9qAnVvkbFCGVDNm0LQGD972czETNkgodSrMAUKs/X+GWh7WkG7wUvceGU8itq
2tOgzaAm4Hv8wBvpr9zCyUYOBkkPoEpkQCADw7eBb3BWEaMgLMPPebXrzdR+RIRJNz3NSGnwFXZ1
K/5xcIb1LImg6fAwUwWqe+JJa2LxWawzr7EKUPVIXmWw+hapk0ciwt/7eSaVK/zIgcDDB1nCqMYo
P/kXuLdyRdRDnazJ17jBI0gw2T/ogto/db0x0mHvUzu9C5Qm47Zxj+KY+N016wVAdO7J+ni8MJtD
0GB7XIKvc9qoE9un4UEAd7mFWIWst+gu/o43o4lI/0x9i3nua/EamheywljsADFU1F4jGQTNIFH4
Bxcdcsv81CmxfxLLKeQiEHNFAT8ULuskWvkceh6UdpeDA9Edhvti7Z9/g7fdjfabP8A/sy/EoqW4
77a1Dh1M16Q6S3Yrk7sA7gJ6nTiNxBVujYblhQHHR+ax/X90ws9cRkkixtSktF3LW+KETt7fT7h1
O0vX3104/Ajr2nrdlrVUgFASw31g9YKbcm0QxmChJXMCoapH40CKxYokYgRRSX1eQYum3jG4+ckg
pCjs5VUH87awDleuywdzURbSA1OPO4QLyW4gHH9kXsbcOHzKBknHZnWJBP6J0wARp+N/eS2Ch1xg
G8PZxUH0iQ0IAKPji4QGKLtRETu0Ub3YeXVH23S+GM/Etxkw++5TSi8ETeSvqFHiYRAUiV4m0Bm5
Ij6h43m8cXRhMgBKc5xLvUhYtINHHSFfs5ipU5f2EeyqQlkvX7tKpE7IxW3Rsq1odbVdme9P36N8
wyfyfcxO6etVVbqfm+wzz570GwQeUVLvh7mktxXcKXd0cDApFD5rzn8qwdwNLYQHwPgtZMPndvqa
kFhECER3bJFCFLbkv+EKFgfvRmkqpfo7R6WYA9+YsVOF75fTghbmacCx79+PdlqKe/gR3uvmo7i5
Izk0YddwoDvgIx3P0c2Ov4E9H3f3cyV7y6h3jOeMbj50SpAp7YbYstB/kigrDvR2GeAw991MlaJf
T3vXpKaC4PMvaPiD2xchWPkWznSQ0hrH/rigyfl6imxb4DRUW09uWQDIdyZ6n0ykso45ZKXI9oxQ
Q4iwgMANjc43nkG8/wji9GoYql8y/HDS/p7jftTNBXYhtCR5TzEesI/eZkjBIuv2XJ6TEu2hkKX8
kYIa4YUNnwRwI5nxlLqZag6rTst4g3rQ76+rB41QhA5Mq/Wnf18s8D+3wnkz+HkVhzyYgLivXHrr
cplTmH8ZQEfRs+BDP6liW/3uoY8mbJ9R5kwxirA5CYjH8n6hiS+KLMmeQfc9U1vErwy8ca4hSKjJ
Jz22+OX9Ileh3+lLt3RFofmlGSiZu2+xA+7Vycb6e4bdY+EpoZyaZTlamC7YSFROug3rjAVSsFkD
o5zDufEsMNKLbqx+2WXe27u9dNPku0zJ0wpou3AQS+L3564HBzKF/TxvABslEjw18+JHiES5Jez8
PaiTuuRAg65kwAdeJ8wX8r16fgYJhMcjRa1pGdaLHtzR3pK9Uf26YhDEfudfRKXI9DNlJmipf7oH
mkHYICB5bbE0ohhWjMi7dGZxhtgOG4igjvq/VMf4pYKc+2u9TdlXzYYN83qNyZh+dyYfm8Dy69sO
eveEp6QICp6Gw0YqQQyM0NeckWvoJS7Vu51/w75CEDv7NgkwxkgisHr3gqJ5z9fGtVGurtUmX78E
mh/wlkWdy+WSDqON02kWlFRY6FnCw/2VkX7/bnUuiza9GsuhYlDMnGa+m2qbUoqmAYjuifT6+LHo
bEQJb6kH1MgN3etbay31xQvpHlcCxPAGUzV8ZK5qCYsLHmYBVARE3Q4B4MndBGGCXARf3pdNlknH
liDF5EnEvzCuNQU83QsC99zqbPERK4J54KtAANpK51ZZyh1ea4TwamSY9z0SZnPgfpDfY3t1PKbM
Unm0S7FO6iG2BH647hCDMeqsRhsdNV6zqXNnt+e4iAMvPr5P1sInma3ahuvLUQBEH1ePYWDDfsyX
v0ubGyH4MMjGtSMDAXpgtVp//eVD1h4RuV5x0FAXgtnVxtsy6Ei5jVv/OzfhDidfbspy6nqaLk4O
3GIC9w1k8cXTG8C8rjRluHqNxyzsJxFyGtj60Hc/gefzun1+WWqgnNpKlwxwfQXJZ0oNnC09xW5D
XDPy+d9gskly7mTAygkcHzgQEashQ3pSfex8ForpNOG1QBWFay3akm2EVS9NVPQTsQiN1UpmyoS0
ml0DCqWWTuNHOybi5zswDYNLJEJXI1Fejoy9VtDq2AMLZ7R3eSYGoVehKnBFzZLSSHhVgY70FkJ+
UNPaBJvTkuNDwYcYOIapS1LgEEdDPx61QZwiIsW4kgZq0zcWiKJjmZ++xb+b27s1auvT7+wNI0mm
NGJbGfLJylDvjQa/wz4xvDGiAXg65EuD+v3YpklJJOL463z6WdsWfG7Gk4t3m5kRESi6VeSeTwuq
KQgXtGVmS/S4m0kYV75OJ1sUS8ZmjCpt7HferVQgEsCoKYIB+3EVm5rj/N6kC7B19MTut5M0zZ/t
Hk/XOgm4mXpFNjt/isZR65vaNo92i/NZjGSzeMDXW7pJlpdMSEmlmVJZlu52Ty8tpFOc7HbCQMqo
PM0ch/SMiM5HT1MY3nML8WUydbkt5UYq898SPg8EJR1FJ3qB6L8IMZj3IVJv7RGxlCHehmnU18KM
Z1MaaeK9JFM0xiq+c/h3lv9V1h5CmWQ277jYDIJLbWv4PguKqEhi0GP/s7+YcKVdr0W8iZc96hJj
BDzaRZL+IWZU0yAwifzjoWKrGpOIo4eGlEdE7VnQb//ujDdkNo5lkm6lDPfx8jDzoT5YZdcmllra
OEtMLXkRTNfQyvp6driuhs8z75w4DJGlGrEFoZk6R/V6dvpdYBOTK6ftn4eX89nOsWdp+vnWxfze
o35L9Yx1rVSLZ/plLAHyL5fn/y1e/pfxfm7PtmTFW+dZcCZbk+wPa7IJJ6Tc6NmzjGlSM4XuV8Vt
ZwDhvRSYo/ok8idgb6JZ1yQHmNQXeLPddHpycVHOoKyIuH0OseBmWWFRnZRS+n/i5QvhYhX1jFLq
H8QL4oOOpWBKKv60adunFTfdSxLFS1izDCyg83Xlmu+m6dnGmeQjOFQN5SbQBeFe37ggWr94wl+y
GhIAO6kMY9qu0pcUPPNupmSqOHNOO+RhTF7UwHbb3v66tke6NOCxRTuPWgdXU4GcWooxgluhZ/eW
dbaQdPjs2Bs73qyq/uVuFfIYRwjrSxKBnvIdYp5+ZPAsM6XgN6cR34+xLOngjCYwZ5Yik/j5KmrA
G4CfLqASgxGAhtBh2jKX6VAa/xoWYERds99yzdF9IjaOf/T4i0ESycsJGjOpYVfps67c45RBqLsu
vnz4f+std/Jgcpk9njyH8G5sj8DGS0VU9ZEfsfeKczgFRMruA0gw/mp+uWjjMUo7T56CC8C0q71h
RQoVmRkshM4CImX14VmoSxqyAAR8fkKFOiKqWizUw0XXf7js4iRV6r9JCRsGxgNhHHsUFzi1EuK1
CH0jLQu9bedZE2JswV0aOfxRHwKOIdKaH6S3/ZqOEhn1Llkg3UqfEpSyrJvhgcVR/oayrv0CUMzS
DCZgYXSL/TR/RLwE4kCwCdZYLVgYiXzD+GIkQMZgtJJaeY+H7JWT2gzqUZh+dtNYyV/P3ih4Etpj
eB8FC8v9Uu1lJbqbMfE6lY/ZnGClFdl22AZfakEUUfZ1xjhd3sz2/edwiJCzlPZGWDzRl82/s08m
pX59Lb2Dtd7hAfya1RLaEvVsVxRE0QzxqW9W6WswhS8KO654hoaX4jFE+v6ITkgDdKSN1ZoOrpjp
owox26bt+cdGSJ1nFCgMguSwSdR6Ve6XyzaKVRX//5+hkUVYGYzgN0XDhBz4pGU4DC+yYrCYnw7x
56sy+xQ8nAeWG1vh+g1Ul00TT599desJ0YyIrVOIq3RPt0cq5U20jL29Xs2lkrp6FDdoG2Ka/fH0
ekamWN46xNlEV0KSNRBm6xZFk7wVgnmdkaYAYKO00HYUPjIJ3Ak4HonPeCSHBYGPCgJ+NpGv3CXv
wGs9bKa96ivXjM62huKKVGz+0mHrI45ziRk4KIYcPsB/KzKTFnfxS8ckEksGNM+FHvTdeZYFpYX5
fNAq1NxFvBVRw4sMdHpe/E5n1CvYNU/y4Ryn3I5ps35jtBmK5rudu4vhbTl6AMU/NbrNVvs4ypTk
uSuIKFFdEap6o5IYEQyGloHAV7qDhBsGxbC9H6+/tAs8m/MOpV+OqPTs9DNfwcgEExdVlc4T/KbF
B8Lv5bx8hSVZQRVzjpeR4ZrVo7WjGRmOdblZNq2xIqKnr68xldg7GCdMgrmMHuVq5VgajAcerN+l
4XY7pfY+j58mWTCZjB2g2PPS+Icq/H5TkRAxVEVPcR6i+MLmlXvP1jmcQCYdi2XRM4a+J1MSgWEM
CUcJKQHMSFYrGfaWph/QXHFj7R8qKGCHToYewTlh9p3RQHbj+NqCHQo65RJhvGSjoEqL1HB7t17r
BsmjmqGRjSspioYW7pRzkatfVy2Vt+O94rzNCt7IyQ2Tjqa+oMHac2iFa1Kmwig5/dHE4+i0UdTN
I9r78PXdlic0ozfAobSwX0v+rCx5EbxPLZ3JLT50RNGozdVxuGq928nFTJVnr5EfrGkR9Xg3G3RQ
/tUWLfCeBU2XMC0KflHnxDrdeTBCscZ59VUPK7DbMAitE7sb1c1bL5UMu5wXDKo6/7NkBjxPL3MP
caw8No7hrMlVHT05Ho5E3JL09yafPLiFr5XVhOg5ViJiLYBEsVfBqCr7by3OyqJrprwtQy3N5YRj
4rQvMpvBi99m0KLqf80N4v2o+EgY8CKvzReltNH/FBBvqzEJDXNDg58nZIOFa71OKaA3pL+kb/D2
SkxPQcWk9LWEQyXV8irxJRO9187b8gCoN3LLKq1bssV4mP7xzWo7a84iKFHCv7t/EmvZf+sHel+9
WkAhn9utSIXpoXDhJFLcprb/ub2G212kGM93/cbM9FfFXojQ8JJxipwVIcnjU0OtNy1AwgLxr5hu
sIsN0cvtaH++wWBumHoPV0EVOL5OKLB+A+ukmi4WbDz74xi5m6Au/YevG/SGysX4ZvMsl1VT1/5c
AW39eE6zHntfKYAoIhPhvdCFWR3mZIc4Dwo4YMLiWevqQfO4kAfipEaZkHH/PGHZ48EEj2MjN3e/
RQRqzwQUle9RIMOqtoUF1yBNYyxCdPwNViuKGrC9Kv/JZ36BQYqknaMLIvT5KdklTaZVoUjyT9GC
Jr7rDWjzeuGKLb7mFQjPjFjRNwa3aByJhAeP3JhdWPVusjA8g1t0e29fkszoEtxjfjxEgbxRi3Fx
xgXSWzJGa7txqCHCFFtVc7eu30g40S6cil8yS4a40vmX/3BPxUtO0uEIBrd/GpU+BRxEZMjx4fr9
GcJnJoN4YhoHLVMEbNXF1hRw9zqm+AgkeerwH2Cp/KoT6C5ad18U6nmNZbHD7rXg1roL2U7MHmjx
TwKbfhZOturyPuMoHIm57smmRaMx7jVoK8OCDDImFVCWP0k5AdIShWT/zJi7RYBB2SvCJyUCzkl8
xxXqgTsZla0b9/Q1PRdqul6l6PyOsr8AVsTG3QyG+9UKlARs+fyS158rZ0DJpfAGnUukX06SAo6y
o1jqR2GVQujC8M9Vul4d/f9hMO62SMvjVVKM1sddmL7qpdzsJGO7EX/xg9jLTGJFKs8SlJiUFW5k
pbBIpiNcwy/IjZYoTvSI0BbnzyC87Jxyh96+gBUCUJqJbFqr5Xna0IvFXfdhDkgZQL4qYzd6HCC2
4jK7Sc0GO+47UQam3jpJCqhycC957lY/yc/HO8w8xqcFlIrQ5L0Rk8wvsOMtg2deIFAKS6wD632P
U2odihaMLny6l/p8RLul/+QevPXkE/KI9Yq5YSztYMGej6qgvcR6L68FodGcQQ+xd1lT7Tw6ME1S
XqCwS1FWg1Po8kKajzojztutdeyFTi8zqKJe0oE697xGlb40OHNEK0Ez1s4+shtDvxwRVeTmwX0u
G1IPA2Mx9d2vZHmuTbnsc0hN6h5RHqLhzxQfmAisFLDUn228iR67tCo4yJjWP6MsuGWEDKdzE+WA
WzVYcEM+NUMdqZN77fLZaBcAHU76+9yIGk8icp6xzAePTg2Dyi9U+MMl3GASNdSjZ/7hzk+wvWGw
5WVlth/1uoaNolIhpz2C9XFMUyOeTAdA05qLincRcej+DFW/+J2kdGcZeV1RzHJ3Tcv3yMgpalBH
FMFP+yk7BtJI34XPl82PzPFuS5fbwO6GN/6XfEC4SVbUXAxA4HhbHWtrFWR86Nah4cs2P1W9vCOV
rVhtZpBJnhwHBXezES2qgJcYukC3JnczAYxZj5t9hj3vqNi5OCze67gDegJPd+rPJb+y0H2nNPFO
BNg59JwH4HNi1F1kH0PSAyvQx2kVwl48YGFNsvmF+qGPyjt6/5oWRWDJZ5OKB6rxfob51qmYsbqR
V0icrgzyk/2g7xMJAFoQT038lttHu+05fWaOjHezG7H2iNpbxNe+SpRkfXc9e7748T5aLpcN7kMv
hA5HqkueDhpM36esRFOrNoWMIwM9hUg/EtWWhVSDo6VAON24Kx6b7Q6qGU+jqPacuR+QzODabZaF
sKuEEg7ZJ9LJrkW8hqKwZKccq4i7+xI/QVHwA297BjUUYvkbPXuCtOqhJsvwo7oIUfoPMbE9qTrU
JqAkOFCy2sjywMzkpMrQs+TosLn0lo/W4E4LqAyEZCvbuOrR1y5suMHIEIxvxAZ6Uu4XYJbBHCgC
YVQfXrPg5e/y9awADfFrOgDbuDmzSDCW0T42o3vhbAZsmuJi7fLDbMPAQnGTECTeGCLbQVM/iSbu
OvryfwTTzl/PlkC0Fv1GErCL5P2hVU5c56bkxOPvWZhPtMGP8KHsfCbSjGSjB4CkFZWpqsw2szUe
9C6Mduk8grXpbtm0xq09v7sNOyCdoNwY7idLrtL77Z+aesOEeqSzVOGKGLxjV/aXXSadUxe4aJYW
YO7/o4RgvgK2zQRxkQeS5y1dFytoVRU9zoovlezXyLpucSklWY+U6nuC3mIdk+x8Mg0iIWTw6HPp
WLG19nG94yZijnVf1NsVTS9srfihbTepZX5MEsehEddnwjk7U9V5BxWmL+1CvuV7bOp/iP02BPdo
LEXeYOtnxTw7UlUn3GMtZsdem15K9Z8rSaxbOHT29rp2hTxs4HFeoaoGo/qwD5R6qNVsWW07JUGJ
Q3yUWxGJ4Vv6Njb38sxNs+rFsIeKZx6cl2CYZNOyx7FC7LQomr19uE0h1fiu6j+cO2v5ycTpUOgL
3oQd+ps7sVYf32ez1Wja2R872SarTx9NpaO63QKslRZSOXwZMVkvzMTGNoGtg+axjHjuN7vm9kC6
hlSf7Y489Ayb8WqRMMrMfZHLJBFFfooKoKVj4RUQpaGtwOcQ45cM67ij86TYkOFbkpgiqPIdUxKP
OA5/3asdGvMhwBINLbaMV/RdiAH5yjZmCrLIY4DsnoYG9yrE715zY8kZ4+8QQvz6cUG1kC8lgTW2
Xj6PMCvXJ49wRDxNd902a5L6BdvsRuNmVOL+yDZe/ipdmKongRK1V8AF5WC22M4hXc4W5/GApRqh
2TFBVQsUIgPA6wabSVknYOrzpp9GSxUPMX2mW0c+CZUSF8yHeGUYUEfBw6hrJZYJWvTTC7JHT5L+
ODNlWVfehrPJjTp17Yeu8t9E1+ZDkFtB0/VDGYbg1ZuFpAG3V/Cpwpe54rJxkkbrXxc7K7C8v/ji
Pahx67VoV6VUtIhsFlTV26Axt8gTnAdepfJCQsltR/BzXyT4xXO9Lg/uy5eB6k7NkcbVsNGOvSdY
2/fPYzB7C31XUlzb+aMecOrqBsvO4ATJxbkSHrmhsWgFQTOCIJeS5+Z2++lybBhXWvvsu+DDk+Ds
kCeQ119KLcXiqOoHE9RF6bqbTDNdyj1GailikiaLHJ9HI6C8ynT2xXE0Shk3bcr/0waHISfKGOgr
ApCn+HnDCBead7KSm1bXFwVwcZ9RDU89qAToiBhqFK04d/kd/xY6lHuW42sXn5/xgERsTGjAtoIK
+gm3Xw3uiYpbQHIZaLPAi5tNlt4eg0wTBUtq2nP5v4/9Xp8rvW4CP48uVlgvu9G5ignYcRat0HMu
DdSffGgZfiYPTTeA2jLQ25eua9zz9j6cnpHsf6xKiRAPWWxXgcd4AVAq3tH6FcDDCIpyyLA14fMJ
6qdbFQ349cNvNzqYC207M/zWBRRlAo2MXtkhdYVyJ0viS9xWf8nJSqmnnD0tuPzimoUtHkDZ5RW5
uA+pPDYYvZuB6aXhlXbxuI1qMKxXmdAHCFYLqcpK3RIA2ExbqjEBDQQENkvRIvcPRaOKTw1GXKUt
onWgYOryjX4HZ0URxtbKkaZpBsV5rqUCTBpC+dlYG2aHx9DlkY8UdWA4s5DrDIhxDwXRG1umCapk
TDbmuNW4JUpGOF9IoyO+iSkdXpzH/7F/VSaMiL640t2QgHUZjTo3H1TlY8J7jxYbvCJyXVmYklbG
8DcCos+Y4UZW4qc7NOYWF8lT/N6uYpG6arPMlUdP3ta+RI6OJBQ9bEyJQrrA0wNeDOyul2j0aCPa
2KEZ3lEe3IjIsahmrIGn4LmbpZPwblATpshIJ+fOAEESCVzWuhWARvu2ZKPPVHDQpF3ahK1AyE8v
k2d5iljhUM0PQLK6CD9cRPnhVdU0up8OSSUwI5HMGtX1Iyvy8XDl1o1D8EhQO70RjojgNbq7gYXe
/xVa3f8o3fgKjZpDe6NbVttw3z0R9OI3Av9Nvm7mb/pHKfMSUQt8Vlnke3LlECtgaty+0HFQ9/TM
TBrZdbv7t37u2htNbuiiAGNZ+DjkaUxoz9mplZjuCdA9sl7HZHf646L2gPix2Bbnn4fBqi3YRDI+
yohGWafnygLud971sCD9Aq1RBwX192FUq/T6DZ6rRFS5RIXz8fAUa2Gch+mHSluxRoiOm5MHbY7S
nJRYGiCQZfgZMmCzQas0vLCXfz+u2oK3HYfndOKwniYFI5yf8/BV1m5HeLENsjYgMGv2fr9kLZWJ
yRGXBWzPNJIiBv/6nWwKDj+b9Pmqo/C49SY25Zeg7KtoIlqgtj2ArxUX4DLRJ9XbGoALQN/SQwuO
VXR/ksXJk/L9XDjSJCyG4AAoyUCYxO6ISyZE2MyhsRc3rl7jzzx9oOr/8yPw3yLjlmjfeDSjUGLj
uc/DtNBrYtShBqiAfWm3u2Mwru+4hjZ1swZ5POfBWB3p9La8V8XSQeoCnLIbO6HUcLohqFMvLQsl
4UGCeBxQyrJP3K6YNISHWOsLmZdYNaWzI1JJopAeG9BGOJhwJUWPpcN/dKM+y3On1r1B5S49MNhN
rGE8OAsZjWxIMqP/qTszbU5ufS8cE1dyPIPlY/dk5/ZT3y8bROvVVfE0GHM3VfevI6bFkXuOGZvX
enWPcwnBsulg2MaHl87QgHuJMHuYU1kKNjMjnpp3AC1K4DyErSQgAG2+X9k1a5qIY6K9C8RuEaC+
Uy+tp4p9kHLF5ir2Ij0x1q+N+LUl4i5N3xPKz4A8INGsk7oZGPJYPMdqhVGlidF3zsVKVYyY6PUR
Ptf1ulyQhFYPR5NEk0Bjkkg9COyU+lxAB9ajz321gKeSrV8PQS3GBbZ2/4+EbjaAUkZ3lDpC+9mw
aZVR0fs3Nam1chtNMGUM/bOkNnnf6yFXgZkX7oimfW/oSBc6c7ypiFDOH5EvcdDz71XusMTkPu0m
RwyVluHYDmTmwfbuidMwY7OfJ9f3vOTJYIR4+dMKWFGSmM3kDgWD4+GKaMoJE0pzPJPB+n52X2yw
NgYWr75Anme6pjAY/CeEH5fV8CSuKMJcLRo6O0J+ePSSPvANoKARnd69RenYT8FCJ9LEzjb1WM28
M02N1ahSwbIbk+vVG3ZEAHce7hOb/FiJFqe9ah4+/JzlPvkfSElzL5dAFJOjoQ5oqNI9Cup7lmDB
Yt4ujjohJO2mBymhhcbhd8IDMqAPy0ZEmuvD55621Kiep5NOZHkdsUq3kwjRn5lVoBKLVoHWGoDc
3nzvsOUD3HqMHtAgvU66+oRHFeCUyLGfI9PyY7hrj0kgRaqeuA8Rdyn8eijcOXMekfq8dD0KL8g8
fF/vdoW8WoPUdzKtoTuAfTPTwHozBzoKNJXfgt+3eSDyD0pL44t8k+9xTYqbk5KNxxS8y5zkN6Wg
l4lesLsygocKJNMYG3Q0UA3EThAt5rBLACnwm8caExJYXorNsRx5KbspIYKbG4p7ShS6MmNy3LB6
v6QkZDU33SJODwKyRabpFKDOCQ5m7lHc1HPQBkUHFDvNjDextE8AJiGn8gzncdziiSQp7jDKUJu+
RImdMSzGGw3JKbuTtqpy8OJYTwHuwKtSVRPiz2wpi3dKHiaY/X/H24M+8D6Ip9SNvqeP+LQstlJq
4KJLynLlH31Jr2AnfXK1FC0AtYjd1LpzOOQ1fVYyXv7bh5y5zNBjxVay7W4t+nwMXe4J5/ZYN59x
IdSNfN+FQZjNVWxxktrcXr5Jdn5v+CXzWazwk3ICMz5EWhgn4EDtNOKoUQ1qoPLjkaoEguDnOQ9y
B+QLU1f1XBpMgbNLb+7QixfOrrN+/XZetfEY7B3jI1Zui016vpR0SUh4PGV4dZJ7/z2I2xNS8ANo
hVffR4atZGpd6GT/vT6w7r1iX7nO9fYAeRhpMGb9U0h/cWLO52dP/Nd32eg9cnPdydMrresV7O0r
to6FLu8mJ+xGHRI3FONsjVb6e4RWUyFccB/0Z1byG4h4JCcRvYJ8QNUzIWkW+ip8Nl35CXfyuhDH
5R467j2CEqo+NjcCU3VYF7+7SVM0YBE0qcoeRH9uYcj5ejiJtmObnPtQsMRy5nQ61MVOx3lrxssu
IIKcLGnfJA95c34EG2pLA1vQsSWLbWDaV8M6kfiCAk0+TPbzwgqrCqadPgdw7vzPtF5Hso3h/VXG
U7PGRnduYFO6JYtRGFo+vM82iZ77LWwmvzl6IPfNaxH6XK4t/gxCeWhogDNj4elDeZ0Y5IXN50Rf
a/MBspsn+HpP4T8U2BQP8xbzTJSafVQkXtBn00QGd3QkGxg5igy5OyRHB138jQinoHuu8g4FKawB
ivqmNp5tS5XQ22E09E8fX9qqwNb4qjZzHQnZWq3fk4IYtNfsoyWTyw/+8q+DSr1y8XUb46tsa+R9
rm4ti3K2icKsc8IylY2tR168Bvrtk1Da+Zo4NPp8WFibT7A7+az1ca8884w0WlfNC1zd/JaMz1AM
PvVe2p1YLoKSY8ahynS8xrJRNFDiSMlScZ5MkHts8CHwkLFpJjNeU5P/bRFhVzG9aV3CNvU5J3y7
u5ej7l1iX07i2CIi5/KXx2iFEuCl5LAeiCTWxuCwkNOT0u5ZgGykcCpJWlthZYU0SBk+ML0pMXvm
9e6Uq+Sytlanyvd5IJ2wzCPCV+G+HGx+Jm852ISqjs8zL4sWa+weTASP3Pg92n9OTyQwtAj9BIaP
IzYvfOR0Fy6fe6xuWSH2HUnNQ4DfYB6YKVPFE1fDXdRUZ59LyAyb0bSKA/oylnGIsvMm8vhGksfy
K4A/26MwxXPyQ061ZjRQhb12I8YnhBmbsaq3g1R3hTKJsDzbPOh9KqessZxXqN3iRn1y1u0+LppJ
PLFl4zbw0xQX3YXpV51u8vvqcYCXEJ8YiRizUlVKEkRSjanV3FPBXRmIJ+weNEsBU7BzlSEHXhO1
x+hbvyhWnkfCocfsdAFhMG6c6OCyy9WpapJATpagsE4sjd9TtE1vLDCcDtcpS4+qxg1wdQpkYj/d
XF4zQazq8S1RXpCr64UYnNayTYodfTvYWhIiSkq81Y3Cm02z8hL+3GCHv8dcAiXDQ+7aJyx0PJlo
B8Ji8EpAUO7zMuWN/zXzThLIZAMhmCgFAneNV2K5BUfe9GyEFb4WY8VXS1q+NpEWfLF93sacZIb0
dWRZgZq8y30L+JVcclE3qt9TOgxtWVUyzF0LrerCBsIwary1+/Eu3rTJGKugpEc/Hd50NdoKgHPV
czjzrcqfR3RswUe9yaqMaFsc0D+9YQ07k9+4aVcXbYS6ZeOLLiWUZ3LXRVh1WhBgXw4uRrzQd/UF
JHRCCUy5fe22rei6K60fXHQBpg3JuwEitpeVnvShtg7M9OX890XPXa2XlDrO3tZw15iEDxgvGcNi
DicwT1rjM9RLf50U6GJTzpDnAea8J0T8JM8pzVt7bSFndBdI1kY7ASmnSjG3zTfm2aLjdMJoXNQC
F7wfYq5W3GNW4N0pH8y73I7GBx9v91ZckQc/pv4STcc0XdV7KjUdaYlq8yz38erxfxwh4YTptH/d
pKwXX2b2mYdvcvD7J5Bx23W57EW/GPoEYtT0cnG8lds2bDw1SMBPCXCsF/slfRmgHwJCubkqR/x2
BDZRSY324zxTjf+IFhPiKjJu5NdFpN2QNI+kYjkdEXa1HMdUDsrV1xOj9RuKTchgvRZc08WU81PG
edwFTdPd41dSka0CTsylfAhPZNn5iP5q4Z/MQ2TLcF2wa6oPdACQarkySdda0nIi+tJ8c+FoazOG
RhoGkduKClR44TZITQnIhZsOeDja/vxxAnMsw9gmj6BnzWH8mWiMfcLuX1h0cH4ATytuLk+SCy9d
i4rfMJcn0IcHE+Em10U8+6FpwXVWR8VFW6i7TOQpcqBhbYN4qeHamAIzcxrubwji0yl4my2N+Skw
A5+Iix3GcfbqfIzT7wtKzs7tc3TR3zC4uIEj7nOBty+rfcBa/pKRER9JitkU6RDc7bh04h0VXy3x
L9+LG3N7SHJczuXcr0ol2VC233nZI8BaDQfV+XiWhTF5NQDpjS21iecGC60/m8h8q3us6QRUd0A5
A8FdMm9bIUJVL9wFYioxUWQ4rtawJpbeaCOqMzvoVSQGY2ncHHjGBnCqHVp6/TE/MWE+jcXHKO6q
aX2ZSUhdtLB7m1vvfFwUC/mmIjNw12MY3ThJmZlLnC4m8B85MaI8l2cX1pD0DCQY3kWpPsV5BhEi
Zq0tVV3dXAmTfV2ewUVf4ItIVz3cnPn6R7rD7T5NYHEie8M5WcV+gi/esOjPnhl5I67KaG5t0VKZ
23b2r+8h+auDcsIecofiwRtPX+kpbr7l0qj/hTv04bcvGulcNRcfClhOfRQrR1tnK+DfsaMNOxD/
VFuRIs4IVzjg0jODqpabtg1MbYLYQn0WxMQLbv0SuNUS7vncy7Q1FYSIeAv1Vbc3V8EzWWesXlXI
SPlMlduf8qNvWgYq8DcRcf7k8/C4Q4SbdGPkqeI/gAk1n0yDXLgcct81q3/zUh76Orr3Q8XbKbLG
/nLaj/UJ/ijB6CTDEQLVsLAbSybMAlJvPysRuYX6bRy1VgHmrOJsBVrzabKAYAn02l2vYsYIIM+2
qLG6/VszPxww4NWBt3gJZxiQ4gWRc3rimqfhMRmHtwiEYBrYHYG0g6sgPhEUlJsI/JBBocyHO24S
/FZt1EuLS+4/rAMHYPisimeqzJxDnQQyY6clLynpLRnkwrDFrGlaKoOsq4FI9C9mNg70rNq0AMjM
1HQ70MbUCgA2+8S24Iy07By1i7JLtTEpez2kgNSHsaKagcpSfV/KEXH2q3xbweUHOfnyVcVV8fiu
SBYh+jsHJFo9DK3E9cTxjgCADreZRT+r6DRE7T7UoM+RhMQQCfedECV4bOmDQ7VS/y3i73Tp7MLW
GJSP6gQ3xL+KqUr5CIW3+Wti20qGL17EhZefZ4gsCuGC3o7NF6MXiXEjWsyUL3Srn9QJFwKxmFE2
AmT23PvhQg8+7es7JpNA+sE686TcqjFKD5hBUqtQEG8Fyje8MG576GEgxGnc/yrqNhpje8nzNC7G
IQERUmAEej/NcrpfVxbPU+bP9zepi+Cmdg8BMmvYrb1cKeUvYGZ9T40IyZUkV5c51aRJqgiBCI7T
KC2sGz8s28YSb8mShn0Ia8rWm9xODNiuIaMjIaizBBhN4XAlrCr8VYHPVzZ0r7HTWJAr7pWd86QI
UmJQ1Zxi8ATRqPxcEqvx8u2WxXYz76xsuYUu4pbHrdrUqdztNYc/EL31TlzjmBqqq9i590q65Xv8
X6Ro84HaLizN2Hfj5JN4c84nQXICYWMtatWwpe40IrXgl/SiUqWlJFJ6iMk6uMP+Vss5MBDHyHOt
dJPtya05AAYJI/peqHbYV/lNff37Gwg7AMsdQp/6/DiQa12dV5ENqMSzOx8232SErLaprA/cZurq
oyP13Uy9RdPNxr3ZIFmcSLcPzcYcA6w3s/4SFA96/EVnPii0onb0m2OvOcQS17rYMuZgZahbCEJE
FZ1XQitJgeYGzpRsGsUobFUgY5HEySAC4Ik7cyspW6fjzHEvlXdGFPm/WKxG6b2EXVIfja95FNpU
n+brp61BZPWA+m8+aky+Hkrymj28NCdSOPLZ90ZqNwm/SahXZuW/6IuhRYcUjzihUs3q4RWz6wny
kMa+D8YUWBHvVlO70l2aGzDEzNppWasaC7UAIEH6I0wb7aYQl5QGKsLrEBUzdp6n87UxRJUC6TKK
GTSjRu86pHYpFbd4mE8xKx+Pm/uhoVPg4q8rmwPSb4yJWAu+C6GVUIn6KytTCkFkici4SJTREafe
Vz6cViVWjG0pgmwW5XjbtD079f2+d8IWK8rtdyaEvghE/E+CM9EmLvXGoLcsUShgTodirm7ZTCak
BakweAUVtOa4a9dX5C0rGxvEHuhkLH8+QUE0A5dJV300ZEeIXJ38C6r+9/xQp4FJbtwy1pLZpIRb
W20hL2yDm+TRmjSJFmn1ZUxQTttFK1A3v/ppFh5bTJUDRyuZXnVSC1mkRdoK8iRCuERU0SDGpXYC
bA9gXIm5nOCOZNnNATu3D4MMBgAGeZyayEayP+p0qzq6MoCRrpZ+eX/VKF5ZDbeHD8ZZZ47UR1XO
I+emozNnEDJd3y6SghYh+h/YFHnwML7+OTrU/KS4MknKlphfyPMRxd5mvQ2pRj5O80RRXW1XbtcZ
pCzUrx4zit6K+xcMzTV2hJTvDW1gB4g8AvNxJZYNOh043voYb+BL5fLLKXJbv1ysPIDcHQt/3FLb
ydD8iOzNgLD+hIAIPhpZoJNc+im7eKLoQaMc960wbXjyzL+o1aQIJlQBlVwv4nCaFtk/QHp8k+we
1BHCUN7SfGo1AqLMEe5ThYA7rpiZ9+l79p+SJF6pSteXKO66yclHz3++9SRqfNjcRBv56NwzMT2E
bn5l2amZ97aLIW7QzYZ/C8Cr5UfaGdzMIJxCA3894KFC+HLJtBSY6keeu08/LCT49abztlVxZ50A
sCUzlSYyqPCq/68mo9gCwsLcfs3dGoKqhBa9DIEZf5yM1eWjXeksyENUgGHc7WGKFyyKyL5wmE98
dw44iHcaBJeQoQAOag45yTdT+jxcyp3FZ0jTOplmwUU21xW2GpIKkXMZFCX2KqBsCMh9NEgk4HHp
mcFAk/UkJ3debBtCF9AlUAbbxxpdiwLolWGkt0IGoENghr4tVbrACwICJ2y83trcVMC7rMxy48y1
BV53V+0EM83oKh7XoQiWdt+LuzDl0E6/0yEjzsOaA+Z6jJ5XXUADwz1uwZD/XKmBznZG7vv3q20u
xJePGGLYOvE4+qlYZZpR7/AdtsFmsL69KRGp/EDIUoWWOk3HrKtKLkpg6W4B13CCySC5H0+HIoNN
FV3qmOQFRWxURmYpHEZwA74u8t/zAxv6StA4nUY/OayJY0gC/ZNGbq5q7wUUmGBdnp1EOp2U2Rdk
CPVnRz6xB+KY3Pmqphv835uHk6qMnNJo8fKTSSOMg/xeTHVY9lK2y/rHRlCcWozJGNnS8hj3yW3c
H2eQczo36zaroa5owMI/7+aPhfeC2rBP9leG7VncaFWFglWPgrZ7ynySjwhHz2jDgRpVx4Jw4dvS
uRZxaPiet1dvkdYAiLnPxBgXvi9l1JQYR0z9uK8IZ7h4FriK9OclAhhD4nCWK4T844A7wY4jE2J+
By5tC3UJrXw02Yk+HiFSnyIc88Xz3ty/gSYS55NAYSVAgmk65D8EHsZqPaRJLPgrVjUuASW84ytA
3g/k2cQiqsDU/BBbG5ghwIna+0yjtT6Oh989GO+3A8Ak+IKJaTkCYpmJnm8Z7DeSkxhuMf+owdM8
5th/1utASxaE2zOfnDlCmo5ZuTM7f15qyRQ0MJ0rfOcLyOXXpgqXwhr2QsbyIzbL/3N6dWrwk3cc
PEQwOfRr/NhqWhhuXq7EOK6gdvDzFL/o3dY2LiZdQK3uZprrLZZ98MwaJBYytjzWwJUpL8dsPYf6
tR+xb/H97d4ZQUs4kCxNJceY71MS0tbmNxoYmEkO5jqwAEtPvNpZs8jEndFYz9k2+Ol/bMSzQ6lO
eW2uIWexpD4zQzNqNFVtND8eBQk1cqAxUn20v+6IVSDIDU0myie1YS1zwkDUvFlwgANDLF1cXH/W
o2WcdBkuURuLBZfOU8TrHx9hgc86/cOEfuGEV0uR41g8gzc3BkDPLnvHJRUP20lJPqiCxZ9ixkNq
3FHKIbo4vsyUJqBwLZ0RxKlAOxBQXztfEH5GjoOt1F6THSokIZXheYQreztN10sL67rNYKAKJnIu
NqS0tpP1hQB9UnlMlSNH1xW05rON506D8zU/JkAxq6X5BRaCDxxkNt83wE1YpnQRBXkCpf8gFnN9
aNS5cl+Hgjelsu4p4BjDQBg8XgW862Iw7A3I8pf96BklR1adUW81ZgwnDZ4+E32rbjQGCj1HmLPn
LBMuN/PjUnHrLnmL8yVlJVQlshMAWx6DyGrDxr4IKHRyRwOXKqIHQfLzudgVXDeqdgmCHVU8MbBb
onTPdW1f35LRQ65lVBxDLCHYaOeMQq+MX7U8thu8tDpLEljerIiOoin2sFvSIWXnVMeuPfgude6P
4jUW/WZFJAZWYLZb5n6TMMU/LXwywHbXT84BAr+5J75xd7Gcd27E3hRCTHXo73ic0a7X6DzKuP63
OJNhEcJvsDxeRHaJoKCyaCuCFwB7xWWmr1k0mmz1Mghs4lJ4gafi+aENNZQ0sItVedE2oSvPiT/A
0iGL3CLiVavmV7m4NmRr3QWKc4ReyLAc0t6wZRDIVeTG5NqbYk9wSi20aeuRnnvSTKzuzlqYKijq
4yDgvzhP31zpHczIFDn2nQTskZbMcmpOqY8JhdJgK7ivsqT2tEvmQ7mAcdYS0l+TYpaIIEm6OuNS
2Ij7/ymZSMghuLGHaReJ1j6ddRaFQlVwhf7Hou4RjiAKskHwJirBWPeDZ5TtYfOEc8WTVfkX2zao
dGw3aOdwzwLQ4yXUGCqNV7+gICLhB6AMhuE8fy+4ldCYr/BR1N9NDexJJJ70iml2Wus9WTXc3cqy
ZjZ7MZOZYflyzfqmeIAu7/dntHCzVhYAAfQIe5nGwACf8EL+XG3HFvaZdz7H9l4Rv/z4wBPiEeZk
xHOSIVI2y2QEyUANqtVATZOGgpbcpnkbzsfnVdEw94X7vK0G7hG0xJG3gmckHsR9Lg9RtQuGA+i4
kz5oX0ruiN2M2fEyHHRqFOFWVa3tjfV/HXunHt2JNbVPVsTj4k7kEmXUaAGU2qe1/9IyNCg1wKnZ
uP0KGLYvE7Fnk2oIyqoOxyiQjLJC4uxtctVykdgfpncuCeJvEEiZG+BGxTMiuiY1AnQXT0QIL/Il
P+HTcub1gxk7x2jLAlno77alP9zRc6825OLePN8cn3qCoctQ6AEJ4Pm3oGVbNdxIAJ3zI9GfXJmR
amN3Ij3Pe4NbiIVw+8FGsuNlFGzt4IGUIwIZFTmGnxGVAUwnvQrUI1NEh6R4vnmTyMQqSa2fgkYF
VeNVYoTIfm9MWtA9eWJTy+nVREC7iOGmFVKeKWHJL1Aob1sh0wR2tmEJ0anWf9OAtGuZ9C16FsOr
hzCkcKzWG/G++rF7h94vg/4xr47DGi7L/pMonqOYFnKaNZJ04+kJKNoR6kwNWQZWddacblq+9Y+Q
eGfkbJg0RSHV9u9CB82mGmUU77hxyTLf0dLBIWy1eMWn08QwkeHkUBW1E6/DPhL3v/S8H+FTlH1K
WUHw8IswV79smGIKJZY+AGUMDKNa+t9XIKlI1ApmXWB+S3iocRQywMcK+pkZeLoe54MetC1nPRup
5qdsAsLDPU1gyWPUluOR82ROHslt2iiuMKXEcK2JShnW1V6+XYqRJMLPgQO0AawTgLFtDpgcHro/
6OWL45kKsTugbp7v+35Gg/O4gdh1Kc6YW8foguBEGXdLwjlJlPV38YWN35t8+wtIxGW+DyKH/vXL
hDKdq7hhsSwTNjOu48rxddRCqUmbWdwdJujHui1O8rgWywrHzPoSfMUy8oTwiEGInuPNK3occIji
VJLfTH6xZaB+mOGdraet11YNa44SsZPO+6C3xiWZzQKKKtY4lHjlvtCsO5DOP/cU83IUqpalcEIN
V91bQRL9xRS+7tuUVwmYrTjcBisbqT83ezq5NdUYDm5nUoNnLjvdkX52xAdC91eA9aOvHV6esb3Y
qFrKtbHtlBliCL6nfGUY/aNur8cP7Nr+Lr4WVB9w6byjXNEM4sfo2KdMqmhhCujaTozv1BPraX3V
8u2mIXC9tn7RC9o5JObfmoMCeah0gGgfbkBub5ptFoOoQ9mld8h/rq6BvzroI/MVrlDZSu20REsf
p7g+blkAi12RlGNlt94R68ud9BarU7Vih0hN7NnZGsGqfjs7UfQ3LZ7Lci+rOVJM4iPUSdw6ghNQ
2PnQGWKT4PSJa961E2qlt7w7lOtOk9zXEveZLdjl54N/+q12A5jwKfzStR/o5XPmRt06gGeilR3E
OLyWvqkRu+FOmjof/VfuqIM/e/E/TcZJ6G+cakrxhnR0e92WQen1sEpxiUaxQDD3Y++A0U2yVgxt
GnkmiMWnh/OpqwxTyvbgvu3v/kHNQiW0efgjQ/8h6oV9magKBPfPTw1RQOzCmpn3neuQMNJv7G0M
kx3kIFvucaPq3+bsMZbmLmb3zeTrCymuKOEDPAjH4idL4N80t+8xNfYWBJ/xgH3Dg+ES4ZUPUGYG
GIzBaF25HZtNRr3hHTYLQ4mNx63i0Dcjhnl+pttEhx4Fz1TUoLxvqUpbwPx2xKp/Vxf9inHxwZ3n
crPkKs+s1pl2spoJR/O/lIvbtKKep4Nx7t0pW7jDPTDl/VRSSQezmex/V4x2EJfbxx1nFXfKUmor
4WAAF4vzow5S0mHLuF9cavEvz6OECQDj95ZpUC1GNmPulVNxj7KcvRovgo7T4cDS8+Xym0CYMbH8
tCoZlRTWP97Yu/7jUApLy9IziFityITfnHATY+PmWzG7PqUZaIduwkbwTzODeNQfgKRP7XR1dpT8
p/uIYbJDCLLMw1YNp7WJfbuYpEzhrQDkHlMWPleNrKnLpU2JHJ74suF2JjW8DrNcXlX8E2eR2IT8
yKJnOSdDIyB2UbaQQdz4dJz/6Pb/dcsZSg4bSXYQ3Cr5XFXbG2pFHtY+9TB8RfgZ/r3gRkgZiDOZ
1BD9g7BjHArDbpPRBjSkOVx3vkLge1bmEu5aq46b4CKLyPCytfWXhbpk+HFUEsDfBXABT3ASraAr
GHcD5sJE+1jFd3j1lYbzFaq4XUTCe1ihBwJOe4Sz3fgd+Sav/o9IK3B4HDJ9gFD/UTfnCViz4F6/
3WnhorYPFotg3wq5Z5ddrhA5oz4tGFK18QymT+/V74ovRNubeN9UcQPwJ/0ld36Mbb2zTr+S0MSY
o55HmF6V2lyRLbFT5tfQEr10EQX12y7WqajuGX+TCTj0V9pjVdFpQcx2Y+wW7ULrw5kJIgmRCL2P
PTlkGga4U6yN0W/mlE2mpU+7DSWjf2HjiCU8p+x7eSQp3DOzdSD+IkuHGKJmQx9z6k37NYEVT680
BMDYlFJftnG1/cOoWRbfAnZ+fsYMAQ7sSrtg9QpW2OJ/BEBrGbw8X8BLFYRrxnX29hqbOu7RmhOx
jQjB4LmlVSjYtWgQcujeqheLc4VMaC0OxwlXcSk3jM/lP7CMEL/PkGCQ0wPU7uTUACOnhsNd02Y8
e2TSoCkQkfcvjjXPZlfoVoMAmtKttHskdwWaBqiqU63JwZkM4KInUPXx/Vli7aMAvEqrLTp2kSXV
1L5HeqJk9T6uHlmgq6FWQYyLWX0n6vfa8+XpkwxYqwW+oW3szg5wc+cMr/d3WqkKCtQBKrg83CIF
GhsmSPZ1ObHbbo95RvKuqAMt03GBBiCA4mkJee5HWSZPfzF9YneO1iFTmqPL3AEvOJwlE1eBa5I+
WAQ/RYvZE4ov9tgubpjjBx8L1fSUD3JxEcgRinmVdblEGJtFuD2/BLIcrKxFbwlSgKgiSTUI/5/P
IfXY+cuP41JsNmkIj/Xl9XpNTFkhAJW9RPkWxzSfB+UnWh6R3pgyma8ivHwQJVf4tQDVToNr+8f1
zltsMs0rAfRb/oabpv2b3Fknxyv6V2rrzj//+pmUuadVz48JHaChXGIagZAW0kuvBQWB8apCvhwr
TgLjflEk9bXxE/Uuaq39Ie9jqm3zJpzaHDcM0t0kkooBzf6P74UusZkMpGw5oP8E/Q8rt+OPDDWu
z+y/x94tqZlOdueHMfNm5VXRjp8DpBlhbYPds+/Ox8u8pVyLw/AnK7b27pecyBTjqadD5in0Q+gu
F+jaK0p3OMYH8oIXyZdoSqB8lFFZ+NDHSHL+CgzBlRFcFhZFc3kpFe6j/sPQ8DAUDA11/HVGilp+
5UzmOkim/Oh57Z48guclqqLdfMppNC39X/JcUIXiyupxhF2qNJ7RlAzfFjx9nvKpQmdmu5tMDqy3
tHCFtqlNFC1gyoY9krLdtb7q9AjhJqinUjMFnEKW4Gx/c9tGG/umXt0Ue40H2ErUhGosXWH0qCVs
9RZupRXR6GblXnGYmE1n1ml2zV5x+f2TVE27vcDMb/wwgE0VBlUiOnL5mKohHVdIzxwE/8tTV5m2
l0jdTSOtCWOSGje6zUbk+BvRFy48wfx6dCp/4A+caB+itXLdaPWpv8sEsPBGb6GFH3ncnNjWguOf
jrb0OQT5Ll/vTlYoJRbeQ3wHrYnbXgU8nohuzGaX+pBVBKgY5tnUlvzp/M9yn65UD+2zNm0NrO6j
wv6w4vRCyo9G0bjTrKWC199mXUWqxKw0WYrJAf0fgYv9OYajkav9f833wJFN7BIvPI5u72+JqVbo
Lp04DwkxSulhYC8XoHpOlXM5puIFyOr38vPiBtbp+EtOXgT5iOTLOz3gEGeKW+J4i9b2N8IUx/hh
3aod9AQ5M4s4xSBo2pEKzrRZgu2N+hsKEy63OZFxBo1MS+9jIzQFKXVl1YpBofh19NUEGcD+Tcgo
cB3qA1pLQTshndPHH2FwuCC02iHXiFyYtdL7rOys+MtrkWvTIMzJbFAaNP6hUlSNg2G9/H7cjt0h
oI/zEt8IeE8/M5eyUUIMgvQWNe2douneH5hHWdUjZqZglpuhBjQcV8bDgjSbI+hE1ywNuJtszMoN
X44QxR+tyr+FRAm081OLjSv2qgjtxKgg6aAjHLCXpFz4AsMIqr+rJsSCk6dEtjdcSLykmdnHkFy5
SyjUcmBZRl9mH25QfQGFZas09veesIWNuYoTKuuXzWvNsE/7/q/7k+k5lgefQxyA3GaEcCXS5A8i
56X8gdxB2vCS930Zw2e3dUJFHLJqo3RvmxdvKOJqwVvANUEkFLd4LFtjZltyF6Dla9CSPOkG3FuC
zWxCYs/ljMNv7lCEKWD7/5fDVTPIH9Z0/xPhqy4vO/voSOphxBjP2YiURItJX7sjhjlyIuN+pZIY
E2xvS8k3zfmCJt2y/BWprTA7zmfKGY0aaOmpGuhAuIoPEx/t9Unc6iaGMjBltpkns4SruVJhc+8S
DuhhhaAl7JY5DQw8BTD2bHnBF7s4VxuJ4JzMVwh+Ddhomrpwo01QIdFp5HzKgESN2YcJEY86abkx
WpYYP2uzZmimDKkfpS50qAkW7FI+rGj+Kwz+mS/TkG5gO2le5+jsk829zEr3OxbtiHcODsdzzyf3
DCGKirb6zmjLkZgIqndS8NatHFC4PthjNlhnD67PWdI70CHyj1CK12LijoqqwEEEjkoq/8CaMqDJ
cbrLdFZji43GIjWJWvd1Mzn9sdXgpajZkpRPzvWSGTSzy6+PU6/e+w8SAjYDcZ9QDOF10+g88AxA
wNeQw5W9eE7HHiQQzicGJE7FBWzmggAn/ceiVxOL5LBjLMyBdqmkSnbKgnyEPVe5K9fd8KzpuTQD
WkESXeqHIDYmwaGBSxamk/ItbEXhMLZwIrNWLxvg9X48hKuZgrmjBYF8a6IZTO69sH4PQN/H44Tz
mFxhqZftQGKttPGM6X2pKN6YTPmTX1jmgNK+3y9gX0abtSOJtVi+Ks7vrRmFRsqTweAqfTBbCiS2
Rplbz0umSqlEtAl78en9Fv31vJvxXLPCKt6J+4u+k9y+8uBSt+sxVHzuIIn2iZwTL539C2n/BEjr
lEpLQL2yWtmvpc67XAjop8i52jiznBnWoTzg2Gv3eMuO+zZj5F7elgnrDQWXJQASMffRQRwzel54
4ljA/xzjaNu2ewfmqD13N/YdkAeMxUQOXOuGXlEAliId6b51UFg9kI2KuGAWcbcRvPcUkg+bQxYw
ZXa+FyJey+5TuWbHF//InP+/qDdw1aO0FuDo/wzktPaDXZhx3V4xe7TIiyq/rZz+s7VycwQ5S4Rt
NQyWfd7sPW8CgZvQfQb/pTr5fhNGL4yZh0GI0+P9+RoqeBLeKI4roWxruMSReIjJ3JSiQnncffYe
2CQ8EFNdq7yHrlU3OyqaLEK65m1zJYIe6xCRb4YoTxE16EbPUV4QzNuWgnzIyHd2raHeNlzjYZAP
8yOH1Mwg1fBx5MZkfaqrcflN5Hn72Kiov4CxkCV3DqGXiTY/p45YVwfBpRtoYeWokIb0seWNl0tt
rL65YCmj5hOdfv2n5wnp8yNUt5ZSqmNMoEt6U0VenWIBKBVCEOFKfDqTexpi/o8d69uUQIa4NyeR
5fdAABgs0yjXFu6rUfH0Eo1LZZopRWOOP1DYjig3kVQJOlrjzJKOL7sWWChOOeCGJ4ao4VsIeal6
wBBxQrIHMwOaLjUPMYTbP/TWlq+QVrBhsq32n6sp7kpZxbfSWGnSkZbKq9AOi2LOTMyVn73NXGbJ
3mW1vMOs5pjFSZEXeuCmHyPW6fuceH/uLIx0L4htPNQjt3Ee9j+laiy+jMl4Tgr5x1CogecBkUFM
TpCJfMxDJvtZTZiUu8prOMU6xZl5twlaeKm//jK5nV/YN7jS3ll3dkAQyLRMpxFbF9VcnRVGQWL5
oqihZwJvUIGaPgatHd4E2kJHRxcnKqp4xAF+hxp4UX7qgsd2/Yt/gyjzEuFNHVNwIfX0E/vmgOtp
3AJZAUNVHKkRNhujXup3qEL6RlhIoc8bJT+5qeHK9gAcmT9WEXEoiNKbefn11h6FG0qIJbZXuhtd
UENRJl3ZX/hkFp2iSSrf5pO9A7SxB77daZJyc+R9J8GOUnifITI5UstUNu5UcozKWTaz28B1JRqM
WQDBmGx/U5rmU1xqStEd1rd5CgQ4HH3WrGCG35ulD1zjaz8ykgm1xoIDpfV+KTfewBZppYJIDbNO
ijXFw6edV/WCKummgtJccYey9BHZX9mg7cgn/ZM8Iwgo1vWz6iwgpt3U/8QO9zruLsrdw66Nyv4t
5bekR9P005yX1Miyw4KkvIVCLh45FBphL3pX3xzcx6IzNGJIjtJQTkGaxyCRH719SWxEaBqNo/w5
gTxEATy5tmtORjYv3Ig1T08RCMSgD46w9Yr3F7vk05520ONW1Ybw/jkvfH8gCUFw5Hkvc54XwKlV
83j8Mk68a3TkSF8mZKIOh9xNwsH7sruDeHYav9H2GMQSo7aWX7q4BrwBY1XGZq/A22S4suWrJ8/a
bgXl+DBloTpSF1K/RhyKbmGWWkGsL5QMm5XO6ef2bHmpt82FhOngLow9Mii4rSwiJOuBPde7zaCe
OaOFr/niEd/ETn1xxQcq8J9tqhNTWuEEOnAU9tsEDoxaNPyplcBv3xV+g6qqQwsYPAHflWhkafSg
bJIg1OiYWqZPW4kSNb1xz2lfkncoVQoYapZWfIVMxpAw89jh7j+HN4DUVSoGRnf2pVpXhFdug0aR
+KAXHhKQapueb3K/TYsgPJYvUm7DUlgDg+adRBIHDrHj21tmuEEdzLhNSeosIC0NqTyq5T7RiOKT
s4d9XmFM027yHFWd8IBRzbOP/IksfdjlPLyMIC5Uve2e10VZwLzN2PTpxH6KwV5yFI46LfEgKPU1
eSCRg+37cdTKox73OCfsSUsR0hqhoqUQ1gldLZYGgewbtOI0heCiaufTUgS2ydSA3CPWniS+Gps5
tKtnI2fQx/frLUlzHcSF+pun+kh242WrAXStIRy5lzZWH0ofAMvjMxkT6am5NX/3jLC8ik+x9ziP
LJUGRbvkY1lSUqxi4E6D+ntBqsM35pq/VavsP15PBDqYZUJ3aJP/+jxhHWAV54gly5MkJdCAYAKD
ymcCQNbPXJvmSqYzLqKlmB+uVrdrRMWSLH8OlXoBTXu8LEsdZ4C6WhAtHi2MBoXASl2iViPwPejP
FADfb+qF6DluRoBTiyatpiw6ewcJYlZvC3pqbuqsg06zI71mFRCriS/chDhPUTGzp+ATWrk9Co4n
F77uLDB+7V2+A1z7yQV0rvKt3niH9OjPY6+bWbk3PPUAHVSeaKwpcz39PoLWvIIS2MFYM+zITfhE
BM/55nlxN83hEmgjJh7HdkZC7mANjCgbfrZjSxUnQOZXwJOEff5ZrX5S0LBiFCTqFNG/zQDlrnsU
sQwwp9R1Z8lHZp2Ts4NYqE/edq9KCKuU0qAH3U+R2H/W1odNZh9/Q3CXu5V/u4ViGaY+Yv7Fih3V
WaGWVSmAKjUHsH/jrJuA++m+tQH2coXgybyNxBvUHqsmRG5gXBSg0h+D27WWO1KTd4wte7BX59Hs
K/yU68C5+CBJiyva34+R3nsCrbf4M+RX83TWmGjrKl1efOwMLFEI6LzFKc8Kyu5R8tq04ZL/zG2E
xbmB0wahqKQvMES7d241qS+KwuKAg2DQ/No509FZoh/n5H2A1i/u1LNtwt5pegcJc1/X5NMdotr9
A/i0T1lri+B/oVXCR0+kj8JL5SZup3npEpOqCi8LzGOgjez3Ho9ze9l+kkkIopx49H1+Gywc237h
+nYZyEvrcfRg3jcuc/hI95uFjPt1rvm4C362sydJXeylF/TqQmO2giXx8VMSFr45HCgz9O4M5lrY
frqN6NpDkzsQfKvJ046Re7m1AP01JWsYbKciCEmelZ+Etg12OvjpAco+Eaoa6G7c7y0BFbNLWGOp
1kx/jsKTZlPajTyTLuGLGc6dRKZzUe01V6DV9IlqFcOGGPrB9n/yFP4sFG41YhyVAZGfFLY1oLub
BOOwxuXQJHhztU8Sc9sAEdfdIoTzxd0Oe8n+6wmrdB9+jN18dPPknfiWcgKLK4SBlw5S+1YniVyG
McVMhhWhgDrl32w9bxOmD5cwAx6WXrCV0T4GEy7RRthDDDVGXGgF2QTFfQxkp/9ZQHNm6OkAVa0t
0iYV2epGKjJavvRYzz4Yx29Shfwz9diOs8nlVNK+yb8n/vScwiGTZGBfnFIhix3rfO2XoM5WmHuC
d+rNxX6w1tXeJfgk0YEiCAzJ5hgOcY49+KPtf5F0alRV3iVC2gwhtKguQ5YQSG0R+oapbIhR5geK
JSlA2bwIEM4O1GU/JR0V4pJJJ0QFE1m0Ci3fUBzPSloWP364ZehbnBIgx+ohSZ3Csn4tw+vFwEVb
GmXe96lS5/05VL1OwXyj3gloDickBa4D41mEOGM9vvbBHQ2NqSoeuXhS5KoiK93GSIBxvj++m1bl
y4rEK2yV/C2nYeHmxKnB5/PCVXsu9chDb1H5nzPt6mr7rhtvFHGez21DkDPyBPAwEwFgay/hueL0
iG2d8C5aYmCh10RMGm0fuOYHE2X8dAoXe1WWn5E/GntYDJiOZLRAYl/gYRRHCcbYezZJ2sxkGrt9
cR/pk+xBMq2Ja18WolXGRjWEeyhLWgkG1UUUgCmob9R+UPWE6hn/GqpaTGMf+NI0D+VLLZe7KYlc
wb3pBfglmfy72+ERIXQ7vdvMfru1Ixqw70cYCgc32ALAQNixlEI7xQslxbTjhCWlA5FjIEGMWoIm
HJUNPQYGbkVynGzLK+rIp9z9W/8+tE0qWTh29bV4TeTfkSRpGTXsU+mW+SdmPSUduqZ13uElMP/I
T3eXZj+03XEjax6VxP0C2HLeuLdqq9RcMhcSu2Ca36iTrB+tFaa+xoOXtBg+MXaQPVCzB8k0PEpD
he+aVPIBagZaU8yoY3HDdJbB4jbU53V4q5Km9AVVkdLkCxRzABXg4xSwO+68DdQ99ZdiqFrnxiAA
XibI07SF0Rzj7wibzqKB8Ne0AUVeYZrUQNovjPJHjyPBOTgfpCNAtSlMUwWVip/Fowk9RjUbDqhI
KnK3lV/gnYH+Fu2026uH6OxRTqC3cJ0eCyJtbFdjSkd3kWZJBZ2mOED8RlFJdze509tT4E10tKNe
4jolxdtmGmAN3nACpDhVb96y4jPk/+MEGCyR6CXB0IlIgE6R2Qp5hGMqHlCO1mIrvNmKCp2UyAjA
0RH14Fj9B57fTmiyedyu1QVjkJOC7J5AIo4+cnl5f4cIWMmA+LKmwT9Q23PvQno+EFaP/gv8xFQJ
IKOPiinN6qIF+20OfEkCpkloa1UEZvTaRr82QJdBXJpGrfeZ4k1O6S6ZgQ6wzhfGu7AQ/hQapAnr
neBacgLORH/r59jWQR413pQAo5E/3kLNuheYhU2nsTvHZtyoP426ufMJ+lGvCNKOlMiHQrmA6Ikd
7Vy7L5oNxvla9xQVSnGP1Tuuyww/XaaKkBbNvlXUOsyqscVtXn9LX1M0/B9kEAQ4gAjwCbISJ5Tr
gmYk3fL2YY1+3+ffhuVubtRPbel1wvlEUS0z5ZFPegczdjxBrD7whZyIgfcxxdTp9+n+0hopTol+
RmC1Jqsq4D0cl9irnuwjJzC+uxlegfO5FTncncIHS+qmbMxyAFnYWSvawCsrJSdKjs3YHi9p3ymL
yuzTpwjHmbG7mWJNXDbnlaiorc/yXmb1rQDgnnlrBkYipBq+yuEj8pB9/b8Y7D2OkyqVnkphCFpZ
tNKS3Wz6v8UtrZerd7HqIgKWKAP0jOjGy+KwSfqSpJKUUKQUF9WVIO/3+saLCpiJtTSLNXrD6H5l
QjPvbmH70bP61zEft8P/jfTZAAa5VIyQo2KrcsPLdAjdvh2tdkSDviCjIRomKRlu+takj9M2r3e/
JQNEFd1o4QJ4kICEz5fzn1q5wMBteaUz0aZzvepZ22agksoOqWW1fdM2fvyA0o9gNgTS/p1ML4BR
tvLSWFDfI012HUxeuHyHn+RTt7lelJWfE/JeQSiXmGafDeCsNuvExju5WewuSDTSOQzB3jkdA7Ni
rzBr4F+EyfW5iUjto9swmLcFA7FBR+7ASUvYPPC1ZJquQIZ1P+sAIfpTG5BuRPXJ3a0kXQYyoleZ
PThVjDFg8TC2PeA+TAd2CFBPPthgjRHUnMGZ1bRFU9jAl9p8n2WFzZZKYlFml2uBtlp9hPcxk5Lg
rh/daP/N03Z6yUyFvDW34l1m+sPrNUSwDWvcAv2zQOKFAZPfSXgq6VS8dFhUGkuikCM4DV4p/oS2
ATzxIGct6IXIsukBz3srzOhl/3Rx1QDEWsARKVFe3GuXyQCil8NSDRrSDRDnqUhK0zpm5oTSnP49
4PgWPMiK+n1TQKoMtReDLwH/pyBlG3al9udT4Za4o4jNEvbG1C9ATgsy+HAUmZ1On9GMorMNk7IJ
i1XFHCaQ029hdQk0tAt4ERvXc2ZFPyD/6U57Pc4qI5CSO9E/TaUwccL2eitztkhsNIWH+Hrhv680
YGdiN7Yt6blC0BFJ8vBXYQD7lcR1JwmiqugQ/ql8gJfwnQPV04l13kpyHyxRXS0MKnzFMJjgy6qF
YVCf9dhcLoJViNdWXEseT1ED6m+UVYV5N5R7lloskiWfW2JW8d9ur/njnPrb5XSmWzzj8kcYg6g3
ozv+dIlgUIpCbW+TxIQRiCYnE8huLxinwWkrhENuZQnotoFihWJ/63VZDdNwvlOi44j6rombjTen
D8HNkLpeqhstAoe4Y6xHK2sBH+1YiCLmNSxyA5WOzYcziv1zXs8qV3u+9fRTfU55/vQrgPQoWFsT
5LZPRvF2mfb4WGmsRI5xzB+2p3SL4+1IfuhLzByW5nxmMZ+YZfDyLNtLUEiwJ+jTDj9PDURR3D7m
6nv6WxqTo2MaNagghg+lcmL65vCurDDlH5vIk+wZHH5aPTCs/Gm4Rix0p5vracytaBK1uFBu20ZB
k0+50/I4HMzqn5n7qVIGAk6v/LicZr0I2t9wbv4BIDO7XtLL80ZJyJkYBiPbqRjScBSCjdaIbnyr
C7ckzm73weOpQTnEkNekB3gWmGCA1+NDg3y6J4K5gxTRH5WDiv5N96CWKcwoEfeeExkVqaF9z1i5
p1+NqVLvv8mNGsEMw9VinaC6RInhpxvrG+qgT/wiDLCtrO+KevasNNRaulpmy+qm62+aMyRVtqMy
kZlAy4Q5BcNFH6rgJe55QTMrRgCaJ9lDUHPvAk9ZlbvkYVfvuAEwua+B5w6UXec64ba3aXcKBBGu
ltvNowFi/QOCxAc4qFq+bjOtV3VYZtNwVSIhK5lEJz76CC2pTREJPDdpmTx2xk8gZGaZ0EaVxm2r
s+XsABa6pAcLjL6tWu70/crpgbH86Tz5DiM8schs/pzMutGf0b/TPIxaE16FnI0l866J7FwGAZRB
zvkD42KQn6r9uqzkUX7lUzmWzsIpW5dVk4tuqoyPm7Kh1sgN0Hd60MAoKIyyyykyvh1ZcyU6MYuR
JlXZ6ccfP+jeIUuJkjrJVn7M/IL1w4/8ltVjZmT7ECgX5VezBtSTULx89Q1Bsxw3hZhjbSHmpBHt
AcAVg/q2slYW1sp3d+H/a/gRNCTEykoJiDQCd7NTeTAyDyuHqzmZd2mIpq8ZdtAk/XfotdW9IFmj
9Ey3AutWdngQbahsdbNZSk1j3VsZ2XxAze7v4vp/hiXUaoqQP6ic9mENw8nt+01Csk4P/C9qidHr
fFXFS6ioN4I86ycFEh3K7XZYs7f1KiOVhUcObzuh8T8acGXfB98BQ3Fh376tf7Y4R+gg5W4mqPTF
JdwZvfVbI393RJgZSUY/eLIr8SFOpUJotzdAyjQxXL1t0apWLn4xgn8ISOJqXmle1hZQg9W/spf2
WRvnGtHlUi1CwM95+5+0C1n/V3Y/YaD6P9N3N3/s7xwvmzJZO1fikZTZh59jbh0nTPkOh5gqb9Ir
4J04BoVfvsl6c1iTJQxsOSuY0pypL1e7bsjKoeRf/sropnvea+vpIvU9ifPI84cPhb499MB7srvt
5hQ9UCiBoJj1aoG0mt9+x0EMggvZQayUagMPb6ER9ng6Wc7o1oL7i2L1JL38yiobfc2slounSddC
csdinChoZrKvmnIQ3stgiUsqpS6aYR+j32t6y0AXZoIk5yExReOzu28vq3tLOPEctDNpyhuHSrWr
E+7U1H2NXp5F5IrUP4RshWJiizviDMhaqLJwU5n7zpHqG6Y+hxLIvhMEL95z5h2xHvZWjDYZ1f9j
HInigPtx/FqLtxm4TL/M9PVLezVYlgn0ka+PCPx/0a5HVPZvfrz3PrOCR7f3Aydcxr1bAS/uUMXC
FZbTuYUxjLEtHN0e3mi/iGGAhTLGYPJo3aYyecBKaAW0twwzISte+Q2IIZz2CeKsFkuWa66T0wdC
wsw5gbLLfQSxYSpGd1DbzVNfQx9SQHLeWEZSWkOExWdW62iSCO7DDF7NlKEqGdzhzM048uYXNTJL
R96gs0LOcf5ojedF4/SLrhrmi2BHR6nH5YZL6JPi/kH+W57hejQemqC8H66e70ypIkz7b25gdnoI
T/+Ku7mdq5ylMLugbGqHSGYyzIg9/4+SVtJnlZReHn9QZNE36x3NZaGrgoXhAEBflpRLyHa6QqzS
w32HiNaRAj6LcN3Ly+mbxtK0mrUErglNuI9bDRSfbIGZYDpTaNdB3Gi/aImnfSHrOhd48JEftLEy
AJIhT6NI3HRvxpVuJbV5iWe96bMLYiLeSK8mvPhxaBaMjn/IXZH0SJDwbohq+miQtrydvVz4K6Q5
HufF73ZoK+T7Eq+UC/qd1mfz+IlLFEgcY8xVPq1NvUGAT3hVK+q6AQD45NHAlrR6QEhHx8do9sEc
1JzxlYL77bUY1pwwQqqJ5aULtBrzsp85Tj9y4KzopaAWWSTkTocbFIBwKhdtwrG6bnudQF5U/yuj
jO0Lnt3oOpekdgrHNMsFHpswmEORBjHIyiqUCUHr4vFXvs880JNgshZ8wyMpQJ2M907ZZiVRN5jz
83Q8lHk9J9QrbuX16WpF1t1h82IGL/tIulciwC76pUOvkTz8/bN02JZHFHyysU4jBQnXJCH8G3bI
sqSF12qc+oCWv6s47dOw5XToY+rGKb2zAmmfniVNURsR7qxfyluMQovQbmhPoP1JQCLM4d5B+3I5
513UPfU+BqPqBZOh/1I5fDfo5VkRs6/xEoHCkCA9rNzbbethXShRFhkLTOP9pZJAj0wj1yrKCfoW
C4h65DqbWdmag7Iaa9Onbgp/zOIuCPBTHd35iFtv7zHSQ62i6aw9fwpAPuHD7yJfeI/65GF2aiJN
EkxoZIbNq7muUddUSsAEdsbOvi+rTaSQBaaonjqiGMsY6JltLJZpCa0IQoLlOqjC5e2lK4nS5Lvs
s/Bi/EJyKJwp2VfHNl+Ox8sEDmbOX4m1apgDfI/Bqo/iRR5HZEC+stSysPRZnn12qFybBDtg/1v9
p4T/Z0AJNix+9Zc+gAvfmRQSwo5tTpSKRFmeTRKydMpJ1SM8KKRuZ/o+JzYkOkhA0RSRQ2gQ9jhg
4G1+ZRxSbEMJcZLgJedDQDSfpLlfuqkgzsN1h3csG8X+q9us8lmDkVS08TVKjDIt1Su5Kli4UWdl
EZqNW5UO0RjfjTMI4Emdftqp1ATpVj/gqLcWRHtvfnIwFSp2GGXtsYKYbxaZCiGvkTr+2ZRBNsmj
FIZwAyDXzq0nYWC8fCFc3EEiGy2HcVqg9r2HQDQMjKyKcrIl0c6ghWnTEfDAsa9fIdQecpk1dbH1
GEz5cVqTUV/8c0ThwPxMLwfSpShEtGB8m9ZIqs+/dequ+L8yQ95HGIR9cJpM694gbOqfbCGHTX7J
kQsCOHOyW03AtHaJnK4l/jDl0kHasY/+uh/uxwIy+pINr26ZeUSB+9y8I74QNhp4XAwMUbj0+Oay
1qboqM2KG79SHD8YyN5JR2erVntDxjyh41f3YX1vZJDzz4/tEObVqIjzUIHk4wNXvqqdiQoDsJOU
bOxIhOxn2Zvx0Zg23qI0GqM5Z3YA7jNko8H4NKCAbe9LtU47AJp8nT3t2umRCeRtV94i6Qvzg8ln
XDHVXOxXn2xVJItT+f2vdX0ROJzxMQTvwYvkGhkQO+fl9ePysxij3Pt554fQ4X0osk/q32pUR0NK
lQhI2oyGn2HexoFAAh5oR51+ayASF/GOpVbdJT0C4x6wE7B+88CbzuRiFCaUoz0pkDQSa46M4pgW
cppGJc1OyNhMvkZtK22M0I4qXnMjigypbluU4ZqsV9zjah8BffYwtklTS5AMkbf/4nrd1UA7l02Z
U9xS/LElvXab8kUJE4G9x6140mrtYTSOI/4yk5jNalb7pztzGikyfQTWEqq61fmpTc5neyhf29tF
Q4y6C027IYzke2K0t1oy7q8cA3kxjS0hWh3xx0TovfH2HoZPpRvM99VXPTNFxiYwLHhlTY+IUwH7
eW0zNXnf9H39uQH8RNNphicbSb0dWt/EI1dqv7cQhrDBqchv9qvX4SfptIADDHpYrMaFWTX+/WkR
MMafIbnHbVLFZzvbKRK1gje77wmgj4Gt6VKs/w2Re+5kALjBxI1qaBHDjP1K3qswW2DS2JtYN6rA
gt2Atwc98t3+ytVRgB3zm8NKi6ZH5FF4f6J5dQRl/ycUiX9TbMkZ0xV2N0dk7SaDDlRHDg0wt3ts
Gi6pkEC6M0brqIHWaThcZGkQPhuPF792Uk/RcY3Egq410k9NcjA5AqGno5TX8IvOErRy6/uS3qHW
RTlGFal3iAaDp5x6DkyI7s73ToMP8RfnydiqmDcUY8bxOfglhp2rZBa23nwIrm4PhpwsCIdjbDIN
ZKPM47Xa3zxkCCJD0hd6QV1yoeuz62nM25n5S598wvvxxuXbVPjMJ/dJJlNAiQUGdd981gsOZmeF
Zf3ZaRkjs3YHwBAUBQjgXtCk8CaYefcFPeM/KUm8LfYTfbo3lHHCc8BJNnJFAOapl8h/1Y28Spvt
HC2DvFDZkvezVCG5uxin1BPCwWBOn/xtFjNblHv79sGQ7JXAUQDJdolCJJ5kppHlT0foSOzqMfQA
l9quaa5kdYNk0thIneqvS7A8RiIVEqep6agSBs2/MBvsOgRg0p0qOVKHLsAA1GlS7SsCQlzK3dfZ
A65eOLg9ybL6PM4PIOBRADtvcjoDhAjDOsn8prv7xy8wQNhjDyPbMu8OzqCAdPD96bu9fEc4dAGX
Nlp8JxSi+++nuw0L7U941OEdfuUswyiwcCHhSOeVFwwtu/UkuqHTUcSq2nMKA3Ado1aSVI0LipsO
HDa0RHfRr8YxkOxS2gKBjXWaoFIvwCgE64kZTMqIKcOaH+sjrPHFhweEGUTATzC1i37AsvXPAdq5
9kSpMUW0+XZwVU/pGHQb2myIJ0XfhPD4V9yBl7FJr5ObXm93SngTS4Jz5MFw0SqaQfRHxEgUYFHf
xpSpj0pH4sJC3I5zu3/V6MtjxyDqaaPxEQxR2qVi88jGRdPbuAOotmdhx9EtmnigCilWa2ZvY5BT
ogRpwq21RLeHygfKV5OZyZEpgGZbd67fvLb7KQrS+PqishIUyBd/OOUFa032cnUKbEsd2jNBSshe
A0j/n98gxL8nHZv5kRs6WvXL7RaS0XZSl0K7GYDmbVHMXrYOLZzwmBMt/Z7guGGpu87ms+5h/yYO
DtfOg8oc3BLmsjG6FJ2bImxGTwSeGBGoyFKO8M7lczKFbeUtxERUPFSnaXYyQLGJ3Vee6GWFX7na
BCRwXoHfX2HeGhzOYWOmxthdJuj42WQSHjPfuerGM3Wd9MlmSgxiFj02HcoADRl20fFKxxW2bLyu
jUSX/aJjEOGAOUhwyr9tZtlSdqr4kiE7yVDFeuSb/uIaxOspwQ4HoyV8uvMV9lOVV3ce+UhmDg4H
TQ1u5uTCF4bcQQ+ZS71rkcRNEEPmOjmPcMWu4Vi5iW9X6rcJgBd0DKVVltxQ7k0uOLEJX6LYGckF
5pZd/bprfvcwbTFLbBhe/BKSNr/qfDtvknc5tZGDImuoQFdQTKdFCY8BHwUSkW0jqPBYskJsXmN/
OEQ2tURV4QpOh7k67QkrPbGaEpIpCaoFEzHAviBVQqCblFGI3uKuFiiGesNZyCrjvihseHS6j7tt
KI3Ks6b53NRW5u10m1j6U38BFMTGsM+F8dyo3JPFXzGq8+8wVM82i5a6FvebNcByv+pNb64VgVFo
eTc5ur6MpSPdqXvFM+MFUfUFmRUX/K955mU8b8wMwjNtBXFjbDJIEbn8t3d5gRiqpElMQwVTz0Jz
W+JWVhkbmeWJ2g5HglXBWVWrbVQNMhLdAAE8VVrC+IuUfANDZ5ActThaxuTLAjmFm1xvPEPiyxKN
gGK7rjUywUwXUphDtI0YB4tI8ZHpzbKHPaTTx9bE/5AWzOYoQ3u1KEw+scMk+QVOBYnaA5BqSmc2
m2UwCKsm5hSJTFRLFLS66voT4AGPzwW/Y6uPUU9K54lIKNfWIA8EZYc8brBAg4z0O3IqLF1zAhUB
y8l5ZXEF4KhHDA+onwLyuciaNZe+iBOskzVQB5IlKmKxs9Ps0u7oQ+q+6924r2tPR1cD/YKLhYZE
N3VAWrmUcTWKrLyuBeYN8N8oZlFQ2DXMVTJ/vre7fHzBO2w4Zj89L4KrMEq2mVRVo7W7YB9OM3VN
DGNEXGxbFBh5jjq/jhffc2VKUx28i4sT54Oh982wVHnt5zufz/1+E3yGRhSBBDzJShJIR4tVOUGF
XhNa1x8hwV5tzyd0ZPzLvg+ouNruHIegTyJ0xTAzSS4OGCdqHusX+aT58dzLeHTc/4mxbcB5mSDD
5lOE1dj8TeD71ZJ2bKRzrz8126IM1uHkwUKLYF9O+lnf9HOVqs5Mc7YjZVt+lfq6VIhEmvbGxOLC
QnvnhHf+ZepD2C65uQVH+vumj+ll5AMfkyHPo+IeDCA2zZU6z4kwXxI4SHSeWEYBrWMupmMtSaer
cDKqmJM1f61Oh9LjEfDSD3bXIolXnbKT46DL2LlnBTbjBOc28cw34G7mCx4YAKhTv5kynuaXw9Xg
vuq5yDzJiADecipqs8mjfB9pNDvpmhFiBMmeTuSJvLTI1kbCNVN2bHn/faoJj9wR6yXVxTf4lPYk
YMZCIYKz8qqEgTrl82RKQzJZPyN4+tqijneG1JfVIN0L7/DdXdhYINsXVvoYPQ1sNMpmbqaP4c7c
1Dz+4fK0zLHX/+cvQ9YQcyCgJ0eH4lx8nv1tZGx+na2NQr6H6GK67dQgaW/ceR9ofXNI8y2kqkBz
S9PonXLxa15NqbSQ9AUANIJQLQ5AZO8dkBdcyDmPYGOFryg6L161c8wSj1FOPHVz60vkKH7ASsDT
2hiQAunoZSRMiT0zo1XKNXz/k9M8BlG/ST/gndyKc/FWq+QxiTkdLQaDj5iKMjaxXxqfHzndh1Un
m/M3zAHGJQNoUoUbrYrZ4yYgixGLPOI8dUzVYYZxpktSFK/rsfl9LbLB9szZ3gIdZPGciSgKDKVH
pCYcJ7dMUKyyWAEgvmuFDpqybjJgISjchT3P4d5vKURh174eILvigKfIoTsMYWFdKcOENs7KGMso
rAzxoTs66UeUpZwEbbbat9eOOMEskXL4x2i+3CmIJiW2n+MQBJnHMqCacsaVGsgZLMxImOy4hzQi
rzBCEV96WM9f3Efe4dYQ4QMQfU5axK/Uc+qJl+hXyTmrEw6LiqZx0wWvIKIbgNskWzV2mxh1s4GX
uMpqJqgpwMoaKfLmljGXuWASFSZRFCzj2rohprir2zsO6nhWqXZRzW92w3pkSnercYeVBsKe9bw2
G8+IVAx4kTBxU8Kb4uzFCnDmIyvjRKjouRb8oMBfHggNss55QPHszArzWJnNs+2/aBdBBgGxn0Mq
GaYMoc6/QNndsmI1ls0MRaS5IRVVhE1PfdHToAwIufoM+DhRqrH7PMKkH++8xvupirqAf/6RCrLD
Nb2JlQ6sgzn/6B/74CisBV7qW7xbM/r8WZ8LpYN9nri2fA0IoiXLsblmF4RAFVlhOMkx/L78ekO5
k7yf1U4vYPz0jkE3CrPtaOIJXjxsM5ezvPFW4vaalflsU5Y54Z/7DSnjr4GYSQ+SBTmn+kem0QUX
RAXxSy82Tynuq87QQmY42AsiER++UlPTUxiIiJE8g3VVUottB1GbSyg8yEOp7QcbnMUI5GICft2d
0lMrDmGYm82pb8Zf4W3wi2bhIi35nqBjMra8JcY0jG0nPCyYJ+rHMEuRyTknRuNDRH4Ks357rtxi
SFBU6nG3xBYJNXrmd4HJEB0Dj4iQVts+PcfVshW23KThV2epGwdBm5eb/rKBkhY6lintp95H9lcS
/pQlFxxIUMLaxQ6BcXJe3bGn4wevo64HBNAz42cWLp5+JX+Wdnz4qgTKYxNA8O+HQA9s0xuOaHar
ki6d2c/bvGhCyg2QQI9yWg+PouEdD4PhNRTGnWZFZBgv4JgrbDTq2J71jdz5k9O/zIeyur/Rkoz2
SDzhqMPh+xU7Nyj2AeY/Iwv9xUqNmA0nxzirPVHB1+qbGmkJOAXdPUSRWxwQPghF8VIu3TAGJQTN
XyKaoiN3tv452P/8a4LzvAoqig5CNdTVZIMRdjP7iMG+YSEqKJICrVJaHRdk13ZDrkDsPWfGeB+U
PCUHbvL9u0u1/Pv8LqXxrs2W7Ivbg7U4uPb9OPx436s4jEJPIwkzJ0iOWCjAShtKfr2NApzRxIfd
uav1xFzeIvbRRq7x78kHI1Dqfa4B/qFPiuR+8NZdkwE39Qg6UBlL4TxuN4v9xSfOJ74PDxAUBobA
EsedFtWq5M3BnLyuE32P4+DTgKW7Tw72R2cJ8nOIfXjKHHQ9vXUh70klGJXjHeKk5XxDcw2Mun2Y
08uRNmWnhvocnW9tydTsyHxdNLtfdS/TUStKKVd3V6ZB+LO/v5CoPhX9QFaHY3IdKycsMgQJJrqd
L+LPSI83H1CgKEESBw6toUmuzEU4yhk/VreL9kdpanf554p9DulGR9GmKuzeyAl8VbWj/ZB643Ov
37e1TWd80fZOLykyewMM/uEYdRy2YMXFpF8hWIMwspDGcyo88lxnpv/UIytE/kI6TxNn5c2hyi1h
QTsvdoLx3hi+TmUP9NJBlRYHF6+KucIJ53JtFNj439zuOkxFx5c//nfBp6AH7+QONT3+EcnluLy4
7HYEr8j2KYp2DdoTniRRMW4qYHvCgubS4TC81RMq+KxywNzcR6RJGLcPv9eHTwU2zNyAl54aowIk
gEOTVls9GfXXIYbw4wc2Us+Y8IEX3KQvpVV7/PHEYM8MmjAXLDWHpD1r6nchVwgbVswUf3a3GXhD
Zm9bexdSlszEicFGbQYASMwc0CxLFPKghk+XS3lIow2E610kvmq0aTfcUdyd5gK72qfU+X/fT1GU
16G+5nVJ1KuygOT4LtWzgUrKdlWYIQHR/c063DEDP1V+KA3j/2C8px+Jn3xcJwWustplH/pJ7coo
fancbusSnDnvPqpgysOV/fHnyko/H/fyoQIwD8mxBhwwbDqbuRC3C8d7GDFB586sSJI3EgItvasQ
+Lu3Wr4ymsK0OBJTYXy2ElSYuenJT9mtlCUgcmH42hxu5/5pJKJwcomLBKRjb5Ejheccgw18Vg8j
aa1dEexsHmLzHPksNolCEKJ6eknvWv1HoXL/FhEFTrlsON5TPqd1MtZtjiaS0zqw8F8jGAUhf3DE
l/XQgCi65BNDPluQu60j7pQD83i9UoNefILlz3EmrTWmFlFeUCkzgOVDfM8phU5LsuzE2Otl4Lo9
7BlEAuEl2EtC34lV6628oLvc4q1zeV2OSni7jd6FyxsmKSfCC6egaUJ4r1c0GZwfqtyvfUbQmMww
NemAb37cZmUfW+gHvnU+jjX5rY8ALL19PB6k+iY+X0jQer0pf6v9usRy0kQqdBByLFy9aLGYQRVx
FE8BoQK4SlI61oTfgw7RJsNjdCtKbVRRy8xJg7fErgBhy9JK4hCor4IyDUC78OsZR+BcS94L5a30
8XKzXBS+V2EQL9zAH3O3ukz10yWbUFNoIN+pkO32Pq0KoTFr8wMpWojyYvZ7/fMCunI79CD/h/AR
eEJhtWgYnzgoYpjUuNbG2Eny/2nGa9zwUD5Xn9QQ5TjrYR9eEUlNvN833fmNE1b9w+sjbhsw8yAq
y/RkyzEYptmn/Y7dRhxmKGVEju4sqj9FXzPBtiDykv+YgR3mit86lzPStJGYQb9Ma8UIGeJ9csP5
law2UqmfVybDXeFeJCz4IFKHOVl0MMUKj8vje/z+LpbB8jsntBTb30AcikPMqc1bokrwYQTnMsI1
RkTB7amGwg9aN506+eg818c7vHVqbYO9xhVDaUO/yIURp7xkdrR4m1R0w/HYqtaDbebo5pocms1I
MXXqaZv2j221FR2k8GqlMd6b12qDzO0n6THtYTCwWeEVT2QzcheTYv7wF5+oWZeoKKQ+h6RB6Jb3
Ufn0h7I/vrCxcMdhib1Add6auMkOibAXm9RpdiIjkXuOKIjiWCju70B/JKKZ29Jjf1zZtyMj1oQl
8R+dTbvRxDLCdprmzNuSJvwzLeRXV7ZIH1gFQvzvz48uIE6VxWDHB0BtFRN08lVrf52iiL42ENEx
ibRV6QYX5GQmhIv6JTwNO/M0P/xjBWkl/gpNA2oGHvxb1JGV4HPQlkLwrgyDMwAAN5Bmge9synr2
88CWkErctxHBIZU5+EAKPlz4TNo0Ronejxxhm8ZZLNtj1cv3sRbnW4lvNYpk7NdrkoS547Uvi3k9
Cx1GIjhfDIcTfBeHSFhPOvnV9SoRgnrqXyYSCIRDhr2UxfmJSeLCUlpgWbjgzOikktquZlMKoBjn
9qtqURdPt7FDMtqE1Oyel367VWlZ+EiEgNfD4QcDkLeexxCOqO5JzSq5d4tRMLVPG3DfuwGvnxGc
Wn53pAOCuios1M/5BSwacnDpxEKPqUGYv7YBZEaCKZ3XwyTZvAx4YN/FDYPPrabzVsPoJUKeG9Xh
jNrpKE6vI364uuUuh0YQD5Uebky6289ST3rqBmnsPMp+s+TddpkjIvTdLtS235zaWeMARu8GzS0X
8fjXvzxm+NQodqmoE6KK/vIBVdR3GnKa1u9kAPAP+ET8024nvIILDICZnHxdBwQDlZztiCplT+hL
NTi4h4FMxt50Y21udKwtsXvUCHddEqzuibCh4AencBgGMSYpMABmti+l2fKJ+TFK8+acNQvbSZzk
pzdJeScMl0cHcHDXeLdX9OZyFVc+aN2KyJELtoZCDf8tzPcCEQiPtD+sEDTQYep2ssiPy3lcEiDp
MOKYmwupML5KCuis0r4u/FD7as83GkV20U2AdkhVEsafxMkAXGWHuOp7CBT0R1b1ere4GknvpqKR
DlCSNsh6/IGDkRHT3yQoYmIxS5z7RAqLIWHAe3Kky7lhwJi5dp7DTcRdZnUsfcvQ5XFdS7ukg4LL
AenUcV4D57rf/WKjhAlaXfYUYrpXYNwaaVFy30OnyBK5CZBMHEYtB4GbVBloZg6KP8ubxx5iqO6w
DGY3QFmKyQr++FYPgVbXyjQp3CbDVZbNSDqFxf8RN1emonp/PBhlCHnZmezPq9pew1RBkRjlfzz4
7FnJ7LJHM8GL03Ezz3tF7+/GM/zcuDghvrZV3Ix4VOlq/+4ZEeC4FPMMNSr5+DRr2IQLkspzH151
LOXK3LU3egIF1mBIewP18n9zinRkfxiey9jlYJYZDc6+YTUBH7+II3//451AbaYi+q3QJHknliwP
NsC40LZZKwsxOpVUv14DHtstXcNaOosefIhaKwHjrHbf2P/YSQP9eJJB0wW8Ez4esqCLK8jAgQ+e
MuwvjGYWwSR0Q04Ymivfk9WrDSk3+aFixtfGXQWFzlg+fmc2tH4FbAuDGuer2frG3B8Eohx9H5yS
HlUZtBeNX0n0fX0KDR+PANn7L40nN9phTuHaY3rh7GQ3v9LIw925GDsFk3YOnwU4vZOfHKOk6RQN
atRXrjlWkuStZU3nDVYVmvZBlVk/lLHG8/EXmYXGq/tUBqv5vnSJYg4rwjjOkbg4zceP3tEHSoT3
y3lZCmp5Ih5ju0N8xLKrJg/6I4V6PB7aTzUhl+obftymoLSFissBHXrYv4g5gyhAv4FUI0IxRC/C
NDZQt6tl8WqB3dSzp8iaxUKNf5q9HiCVfUPuMiypz6wWDwDbHmXP6iAyev6ngv8wx6KWaJLE9Ttq
2TExZXXccssiiGWRAdSQk+RWnGbm14mrBpBcOAv39A3sVLQzoEKS9dCtX3NEJKQK/NAH0lHs2yf5
v8Pw5jQ1I+PBivl8l8gsCjoCwIyWsGUzySU3buE4O6yHZimq69opJ7BmyXtoITjO30GzyVdReK09
raWecPk6KYxSQ9yK9EpxFi+3MJ/+wR9vsrCY1cB15tcg1TXc1qKlXudyPJkRXqxa9GieNVmahFOd
ox6TtxnW7l7MwJEisNjJSNB+vSM9FZ4a6EmCgSu2ix2FwkqNYORChPKBMJxlEg8lXx91ttm4mWx8
NtqyN4aX+Mge90cB+PuOyrrYZpmUhIHt+ve7qVUbTXpdIdZ2EQHLbkpbLOIz/Y5YmvSeKnIU0jhs
gIXhhba4tVvlz2+3cgiSsmc1pz6zUp921IZrBT6SvVly1X9JUTyI3JhlgrukiwX8hQUDn3jbcuvw
oSuVKi7zUajfNz5j/qHaW3UZDULzpv7wXfeg3zEqUCgdNCN9heGrWz5C8ooo4zc4znnQxatgV4MQ
TYzlFtb2NIHgk2X2wAzuoRb8CYzbOFB4KCXYIi+Yzyg4PYh9Lm/ShG4zABBKy3MndVw9NXneL0Sp
NY2Vprg5lDQnAXAuoaFXbKtp/VOes4oqphEY9RcsIScyo3mSyh2hQJggfFgqpPDIadTrc6MV8/ob
I8ahOepRfhtTfpLZvVcRqaJtm2jg25iTQgoB2mMWM6yx0BRvgdNtX6fS24F3k59MFzoCRNTWJK7S
nZ9bI3MCTKgHSWWCyKJy292UvU6vYOCa2LBxeXWqT1ietS4ZnCCZZWNTCslWEyxrP4ml4IK35wp2
HR56wAPWEMuS1Vcam7JHWEIuSCAtPd0c/OpDkH6jTR2DMmoazOgrgxmdl7R5hE/GP5X/ekd8Qa4H
m6tsvcWjMjmjV1naPrguauCoFvMEqP4MCqHXf0oDrIWSDR0VHE5oMqNBJyJePKFAY2lSE+Auj4fo
U8+KwdlRQ3fMPzUDsP7gpvBW42RroGJgg+mxpQpeXqRPPc5BexF5LrEaJS49KSL9m0CFeBUrH4DH
/iSGWG4cWygYu/flxVmU5wI8ua+wkTw2t/ELl3tmtxgcBPQBJtuNWDI1gEPP5iNV3KxTEbu7UnSO
n0ckkDjg/+ydlwtIhSFeEDfP40NRh9I1VcjDlZ8mzJQ/KlDAKmLZf5tVghiQLUY+CM7IQRYNdlwy
9vep0/jN/tV3/fb3W+WDnsrEuM2CaH0c3Q+UStMYAQXaOHiaFnEHZg/IbKZ5+xGEgmW6TpydALZK
NgOMWJpgqFrR2oeF921ZA6WOQewMD5kjEOg9mfqbBPbOMgiQgH4A6YLEa7ZLSDrCSzVCexrVLK3M
lSmxTCzd3MDtMxws8Tv0U/oqxQNxgiBZoWBN3iGXhyOEVZ1T4lB5VDwtRbsiKxCcI33z6xtm8wqE
F4iQ0CXRObfK22tZpGvHQMrSZS9/5IlHpRFhzmE82kKH4a4nW49N/YaJLmezQu0AEf0X/M2HVP7x
DGv6m4jYVoAZ6rfBQLTvjJisqh4jtcF+8+JLeNBuaBWgaReBYQBFjoYlLOeNPxV/QLG4Wo+ST9MB
pLm6XVFMQ8EfVpZ+FO9+73kD/QqdWwJAYHruWCLVRhAPCg0oIbdUqkJkyOMG8ws8uu3zfdchUQsD
RBFMc6eY9intbl/wmTWi/NLmnudWP+sXSMoI0Pcqwy/XUHvVKzU8WEgZ09AGR97ZeDPIMqzuBnB/
Dp1dwmIQdGdrTZn5Tcn3DqIS3lpz+Pl3IbAGYbdArU3d7/LWG7Za3YKYdlA6qM27v/xqsIvdSFxg
hqMUZ9oGWW9UysDQr89HPRgdL7YfNHnWNmHIoDUz4MCjP47u6dNeTb92LJGML0VFcQ/zHorBYi5r
swNhdx//yIIRBaeeMDrirywrYFhHXwfsj3wHyx9BBfCauiQhrz13VpA9M40s7ad8/z6QElEQdEhx
47dl1ZkU5f7g4yq0xzu2AEyFLp/CWH8O2ttv9eLev58EVdeByxk2tqpiQix/7g35y7u/nf7nvYT+
x6W82/kjvX5gTkczht4GUjx1CvVrAcaSxQquzwpgJj61eXoXxuXiwvr9F4OGZwTAGwWa8WhyVeNt
2yd8D5S2E6nW9eDx5VQag4aAJ5ncDQucr52v3SpoxC149UWh3W5ZDaLQMS3vMnhziAmQKDo3tvU/
nmMwG1LkB++LVYh/M2FknaCDJgpS0XEATga4f1SWNx2VH1mtwqXiaTRUGhqy1uPrD8R45iP19gsA
v6S3J18GsjUhiBt7JEoMuVLDlitZlXtGrCGrPUXU9pOeUnS60PyvAiJ8YhEfyh3uD0ryTuF9cko5
eZh0vm+La5eXosAm6IvdPJT4gfBbbs7jhcNqfkpAaaIzifZ78JY79C2aeIoQ31XcmHcHC7zSt9MJ
qKQ3UbTMCQhoomKUuasKZvqfSmrqVQe+TrEMBFWJ63icKOEs5GN3kL3/3YfZY36dzNGs2zAe+hmo
4xDoICFlU4vXVaLAxBU0SM0KE/ZnhvCFGwME6sx4V/KScInEAG3pvhI9VQIooVlawEKfDHZRHsFg
JK3kQ3jhKUpc6i9/Zjey0FzhSAT7hrpCbrTBk+MzR3chgvJT/MHRUDDOqBdP1y/CoLqbJsdxcGt9
MHwj2I/Gulw9azedJTNg6HhuRGKbEmM47/BSi7Z0xK8DFHNzGe4EYp6XzaPmYWLp1D6ZRXu8DmSR
Y3EksCJRaqj/Dcnd/cs9UFEjYn9PAZQNZ7RFIO+5YGniU8jkxKbm8NYzzEb5uea1AXzULpIklKHk
Iu8vSzZtaiWHrKveJM67ensaHu4pOXR5EZWP0/e5enww9KYb0jLNBFgXn0Dt3EY0sUianAmnJwmV
GEk49bDcC7pJHtBC4QyRz68I40kOYkSioCumNthV10g4yFECJwJOqcecQe4jVGGdqUEPRl0agyPW
Ock/wXZn+j2KJWm5wBN2JvG1E0QewDcrxqTIk0x+YbqJPAUN90tsxr3G9M56zneq+A9/kWcPtkjP
6j93m7JyoSkvvzqI9FyHcWw2tX8UghbVKi/pE5F21XkGJeZb6NttOjIw5MA1Ra04olfpqVtea6Ww
fnbWfsgFOFJfkj59CuXyUq38/G/HEjB8mbMFHocxL0Tb4qJPBPlTUqfzZGevuke9hx96E1mOAeCM
ZouR9dqFHAMnTpGfqV39SEm0dq4feNRmSKhG/MMAwqSz4qA718u2JSMXe+9VUmCk4989GqGRpAtU
dgUYWDGLpWvKs8y3I/M29QTPkMrl/Fda1fjtPkbbkm4Wt/Ek0My6OksqepdRrtVd23XjRwZLz9ZJ
gL3J7+kLxD9zCAw1XrT4oaZi/vwA58heUNdvIqVDlpfFO62C2mDz7NH3+jcIF0Y8DAisgTMTj6Od
DP27kIAv431KGMPppFvRbZx5nX9G+KIrOF6bZhigLRtaIu0SuXHb4zvSTwmllb/6KepcHc3OpiAf
w3ahcbejwb3bYTfgEy/Fj6+s90xp+SfaLYk1q9DiXbF1A87WD03YeoG4fnI/D8gvSIewrLeCoV0p
WGKW3is/Y7izP015Fodi2CGkOGSpiRvi/YqS3gHBuH6scN2gLo97Ziysq8LvkNbGkjji58Y1wK/8
wzK7phdlDFAeYpScrMLoBN3OAD2oGzqyKx8bfRGrudJqP11PIypDct84v4f6jYKVKyocaBrekOuQ
t1klvUfT6NAiyaKOWiot6H/iPsDBgzI0yuc5GDHGjODvZBMzqbm3qhfpvACuzcrZ/Eu8Z9QFVmI0
INHjPWBatPOFF4BE3+4gx5cNEMNBjqxOFOJClT8JvYTfUlRfeL2/NIothAD3s121Wld4Q6Hbo2su
kgGripCk8U52XiZopyLERSwKAFa7aJrblvv+EGtW5jpbCrT5AXzpxOfK1Wx/Ndh045swqD9ox5pB
ZrQcODjlH8MlKWDX/bfdwT/M1qCbKi9UvRRA9Gv7LvrgBEtrCuXH61toDriaV6sFBXukRMN1QSZI
HX595Ks/8d7cwfraeqT3wxedBdMcc+MYuFvG42F2xbUKI3Yti7/sKbG4bBMBKDw7euTroZbLE/qo
Hr3WlLNNO6Olf6XJTq6i59IKe/Cl9hwxWzHPENdBC35nQQCZMcbSkzfLpyN1cP8QSrPkeGK39umv
/VYBN9y/VMB+5dRXDVGOlbpBFaeeWGnukv7zD+PU7oUsgXKy9uw/AY40zUh5PY0ghmDg8yMIE4/2
mIISolwsZjit8sSGXxVlacBQB80EXuoYSyuZzWnb1L8gY07fqXSxIUCZhpwwGY9btdbfCu5brFDg
gADpo30vuhXq5c4XMyVALsRAWMJKfEKDr/+ka7XxHaEW+HQ/+5OSAV9VQcdB1N0schKRoE6kkuoU
J080SxcKQcMWjH0+pKhp7QBxh+7qkKc7v5CYO7scEyBSvhjfr4rrybkfPWl+yEj/NBSqJatrF80S
WPjSIzwhJpxWwgNs/B5qbD2zhZYOAWCB7XNImMK3TcMQb4s7yjBfqZD0XS8zyMlKZaL+zOfHYHvo
DgIZ3EGbz6PldG5Fqavm/otuRINxINW3uH337FYoJAe9r801p+olCfn8oQ0/IGhMk6w4UCJH79x6
rJXJShPaDZJzrXLG4h9gdhuNjBEoR0gt+xNgG3DS2MzE0k4QMTz+GKYahbqK173n/vlr7dfhwe0H
VeABDf8oiSVZhIEdxibkQKPJ2ofStjTUAWsf8n/j69UbcLLyWMN8fEx+zmoQIQ3wx9fZftZSEjkB
LKRY9zrWfvaBfvUGQCVmgnUcpjcEJfkdDNJs7PyuybZo7ABtkqoeMhC+n4Zt90r4miRoyR5ulPBD
7NvgIEy+Q6mQFC9m05OIs1F/MlmvNB1+Pym/LqHpyQGMdz/wREtkrBh2M4xc8IuUIZWeceBXbtaH
u2WfOuVsa69Os9+VPXHw4KMmBelHPP6BN/UZzZw/OR1OBITWF1Tq5S4pg3QU40rfmVtxoNSzyPEI
sQSfdSiNHTe/22Im+GLQt3KCDN9s8nkYH4w+InjzIHI+CLbEqvOeVEfV01pX9mwbTFvGu48cfW6B
LiE/pzTMBj4s7MkOiMdGgfzufr6l5wdUZUVvJSmUwPd+ZMIT5U37irzmuAKXIe9viLWwqAegntPB
mY6+Kxh7DRsFY0XObkV7/SJIxstYIpnIupgj1xPg8XR+2iih60Ifvu5SQoWRL5bpvgx8/5r1s61x
Y/YgDXEore02b8DRHdxz5Olpg3o8qYZSsi5q+BZ5t1VWlRrY7tKuUa6Ofwz0XTAmUZjaIxsHwOFq
CwvsF1ieikxMv4mwVhW79aCcBLedV44DCq/7KH/M3EG3u9DCoiyOAMiBA5gWtJFM9O635tuhH4BE
J8C59PIklsxYM2slLZLmlA1O2FaSp0K/2Ibtf+eVeynFKVy9GN90N1YExifrSePiiB0GkA+H/AMq
b1CdS0f9y8O9V1FWG9pJ5vZk0o2gY7QGqDZMpZVZ8nYdTad013ziJ+Kxz2+bOpl172yvnag2pLf8
4daDYOkhy3amtOwWoksGdaLoosPVE0utNs4KuONENGhQTcjs5G2Tsf1xYg1B4NjOSznPahwYCrJQ
6kkonWtpdh6t8vWEzxbtzCnUHRgtdjP5k8pxUsUoDipO+cyBHtHhOddEpLcgc6LH6f/DF4I6Ad13
rJmDa3mEjf1+WxQ3T6mggPBiCrUM3+XBFBNJFmhscnOWg89F/C6PMa2vkv4CdaxVsW5SI9p2Cq6y
1NoG34AV0Bz+dFrkXyLeQ38L5qFDI+mYd5aAOFOsXXzKINfEv2uXfgnu3fwVMWoik1MUf60BSN2Q
PftzjCE4cqJb/dqs0winrn9ABIfDHVqdQkuYwncVl/mb/lgvQn0uWvmzMmGtyQ+LbD4r+1bpsfQI
cpM5nYg2hWBZQyXmsrxML2ncyDTg6tOQLhnnyYFrm18NakHoE30goh7TJY7xOShl+pW4ixavNBsv
wm3qN+xXa+SuIbclOphxwS34YClpEBULx9+cUSOCtO/kMrpv3HHga76uzJYZIXHu0WN2LN+RjWbz
e8MnB2UVvLzfOiL6fmps1aWQTdsBES+P9iLv4hTPLCBScO5eK8IGDh2Y9YM4S3dqIFbzS6+irK4K
kjQeqsgvpqBUBskMOEcHqTfsePaOMb1EvSXvm4cPsXMQRGiMpQV51Rvu/wS3L/lDNDOrfMaftTzL
bzsL1dBIL2TJ/2cGh03E6UoGEneRoCtJiYeCAZyTl5ByPlXfbPbwoB3pJqpYxCGBGWaEAuUvvfh4
XLocE83CsYy8LSv7iI5wRgJkESnViAE2AJBUmFtgYuaBZwUm84kOYy21QpSinjxkTyoEbS9rBiiC
Vmck/FVZuFD5J7LQZblUac2sPnRSi4hz67F7oLgZmFlOeP8PGjcyLZjPq9SlUnZTXnu0bzfaVk9x
jDPune+dEepP/vvKov3oHsWLI+BzQbQq0ekKzu13z4TbsnrVQOaaGJcK6akhV7+8kaagbjjKgQzT
qLKnZLKTf8+TQGijuIGMKFMLRSXUbVSyJb/bA9sfMAsVnX4A4ciWxF08MHcf37Fh/mzuI3RVdZiV
dkIIvV9M7Jj8stBa5idD7rskrU3UtYGgmfl9D3jyXJJOfQsZvESv72B3D7X61LB0TqParQXJfY9p
D1NTqe0wFchq7OMHuAyjsIOXeviB3p4Ipokfyy6b9b6Qpsd5Ejcfiynozg3Fw9C0vnKkPwAk+5pO
Cj/6si2fMP/9Ufn8fAbfkFZloWInz0YOtgCcLeZShTXBEmIew5yTmZ4ozSrxbNd7o5fZHN/xAzpi
y2pK/xpCUZmzlsmruF5W4JykrTeNSrdpOtRILsKu6UKYdhLCOkpJVFS8z54pawqdvZpjYU9pR8cY
4klSwy8QkyQv0IpAq7VY7wucRagPZvSE91+UZ9pTeI+knVFuvljgVkoPbMmbhFWcYUVEk4Th5/2e
CSF2Am8pGCyp0SJ7BsyVgDR1qMiAix/PdmXm5hKxiSSAV6o7B8fQlNa3xWHJBC84ZHJvquZAVH2s
xi6hQ0Ld6lfaC9uV8zeO80+IVwa/nZOCF4HlJ7ZdRd02S8CTYRgLTBBAHY/BgI3nbMwxT2jG2ZI0
NwHqQJniw96KJRGCy1i2x2IhJhkVMXue4y5vqiQqLH+IbNCSgewKCCo5ncfDz/lVy7KqKrVkbA1+
MX5eBIhlGzxBDaBWcTul+4bW+t4pejhxMcz+pYZzt6KE1f8jX72w1yG2qtxDtF61DCqizzokLzOF
9P385VMJfi/01e3DMYNRWt3QB9XegYhaUWdmsaCqXfm7y2HYe5Q0ay98VfY/jrz2OC4oPi7kh9us
xbuJviHyDl7VUf+M3n5wwsvlZ5/rwSZ5Hsux2i1weuTNa34lVcpVqnCS9fUoSUNv0ElCu60Ce1J+
QaHFmCbAXXT5jTJBAlu2gKE8+gTHKJT+SRac5ZQxWyWNrXAWXBfAqMyiM14rhPHZ3LXEH2F9Ftib
/jc4zJdPsKUzg0u4ETjqj0t15OEH93bYciw935ifYOv7XWGS0J6J1YDhOQrpIISew9/uf+fksQUP
1pcq97A41ZYUWmyMPdrGiEuXjv4NAVQ4KrGpVQXDigPsvCaL/UP7M6o7hijiD0N96L0crFfve7Cr
3kuMtUaxcPpQxA7IA6GD84u6AHLy4iDfitPrvDELm58MjEOW/yiXR4BNondnZf37T0yJ0716Ix8f
fD8FuvX+XIMYmh0L6oFn8L6sjw0KeUIRXg/grGfskhtd69tjTePcQm4YdoY9pSu6WGTIfQuJEW/T
8va8p9Pu2vAkLwI1w7Sue62qTXT+yGLVTMeE1sQWv5lcsTBSzQBzBas0HEMTFduen6ha9EhIjSmz
MJ/RiFzMURffm+0kV3+HFVYKQyR+g7CMiqJCLn5dtsNmuPWf/I19o5phIlc9+7X+yxEYmqBS2Ekf
Throg4FwhaETivtTVTEedQGDnAF2QasuN4mtNk20sC7vD1CwIO0I/bHRmLJFxNjXeh4XxiZTlMAB
SJRtnw7g2pR+vjh6DcI3B3ZsbA7auJJSRHsydKPIRnf51yH4k6JbPUdcv05rvS3H4qt16N1HUbv7
MaV6OLmXBZBzvwAzUR+VkhTqSEnpkqbR/kYQzL0XqEz3PwmqpTZ3giOHAVgMWhDRhm2bKghV7AJn
JV7bYK/0rSBWvAGdRDzkrzFWcMpT7cr4Rig4aUEmqb3HUc46QhKrHE6EjYSyTUuO6RL+uBnTP856
NA/XNY1zCPbUw08kQ7BsjBpGVa1miMRf3NS77X8/TmzAnl9+TYSHSP2m1wOZvjvUAhIn7jdV0hsV
l0I4YhbWpUG4i8uOmfT0Hh4a5XHgrLSXVZLnwLg7kvoVszD1nNNYMnPfBz/K0Xv9vdWZXvGY0NNY
Wqu3OvqnH+5l50HDDNTQ3l2D6DDj74tWFiLt/2TprWBS7y6gdYEOjdwF3B0zyTCiGnH+aISI+zHh
BFf3KKmipIALPI5U3ZB6vLZlf+K5cjZTNgqNgya/MEjezGU/DdQ/fVeSGDLgjm/G+3erSXTFlLxd
DsfbikSywBB7Q4r3yDGbS75AhS9utTwKEm3Qy/EVfefU62/piYX5WPCPavccDM54UA2Lf6Rj02A6
leA6aHzR1R42eEzTY/gnrSQ7kS7XjsGWH/Sg6SMhFHBoSs386G3aee4VlXrSfg9FwyOZB8Tvda+K
U2VefUkJQ2bOpFP4kGp7bWGRphlXAOV67eauhqLDrKcfBvB9ZeRl2uD9WJapUkCGAxk5GCuQ1eTX
TmrmqXEAwYi04wHHhg64zy/CRpZgUFstmS/SoGjVCzqzhyPInoMGz5w9XlJSgJFUO1VQO+nGmavm
m76j5Zj5HpoZSE6MIlzhlkn5NPLNMHdv4gXB/bSxaGK32JC6L0HWtVlFALlpYnXXg1GD5qpzyCNt
AZD3EQ/C8ytxtfqCiom0NmUa4M34o3IduDiYZqxLM+AxCWYk2DHMt59kFEQo2iz5/r8kc6SPDdpw
t6yB5I3YPM7VHbBzbLQqJcY99ZNd4jg6tc81ZtK0JPe+ixDxhTkm8w56kzPARwxj83ROGs5ZU50q
oAhfzbqeARPATBs7W/EVbYNBCeYou319maVVXqqLAMB9hsk7you9eA06j8xf4IcBhTJ7uL7oPHmb
m32rEtvB/ZAJ87L62PogV/9WAs8TD5l5mhGMHW8FqMCiGySM7CMQqcCXP8Xf5DBRpj9p9pNvYkU1
L6KewvUvysCfUETADU57ZuWRSKtb9Lmr3DDm6SBWb5MtUJrNODJIVkQUMagjKC0t3OuYR3/h4+tl
UTlfRmV2qn9SV1Eg0tSRdKWttBKPJoAULhF3lKCOXL8SiBAsQZLYh9fSWlGnyfeYgYHHcD3Emi1F
lVl8KWf801T0PjDiIUgIhzMKvtqD5wZcYNntNMQCFUDO64qZq1TyMSfreDt0PzQT5NQaKxrw9Lpq
3vvl0QG2Xb/eeh93m07BrckbDUCQNp994gmjFLmqSEjOt5s0s3QRR6iGSoVl+L/9UNTgqhBS6644
qkgOGjwLYZmTMkPoPlPs3BawNOeBQjx/8D76jbhwj52e51j8jlh/WjzjOf/4Oti9JX+rkmo0u9Jt
xr3H9OplNC1EZiImNPSAV8zqLMysOqmn27vilsUplWUWskwN7O3BaU+NZF6Z+4qn77SrMESfpk2Y
XEW48vVNKRC2oiSeNpjO95Yk7mqgx3HjqR+X+ZddHELN0RopKIocaH9GsriBEzFQtQp2w2PXVscs
f1BK9duWPl+21xyLqbwQEQoo3lrUYDaEQjgy2e8woCu2MBbWGtjm2hiKvqHzBIEBYW98UE9mpkzU
Aq7T4q71aQBVh0tPX173lBBVjBCRfps5C2iNe5hM9VypZkbeFJBIRno0BrrNss/dCA/9TioO3EPm
SjL2gxn8B74eq4rxftLmb2qQCzYX2ooAWl/iDEF2BD+S9yZuoMIcXojn/hLFTUsRJ5c1W/thEw2B
ruvap+C0n6cKU1mFfUc/ql5FcVM2oTWYcsBabUEDbm7apDpo0E97woBCVdQo6ISRNJB/r3XcPJp8
j24XDDzQtsXhLg+IUHegA1rnqKrqbA6n4iyCnkMcJDpmP6BhD75CX+PhMxxEXymhowM+JHSpol71
YXdu2DH4JK3e7h5lWg3oQr0bSsHtNFunTfZ4TNPYvONdDMQQBQ/RU2pdCcAf5ZDP/LGq9+iRW9He
H9ADTvCF2IQPbEcClXC9dpaO9Lv50oa/aEoLGiKp9SjoVjW+R0wL2XvG1MFJZ9zh3t60mWyDGzns
neeQQQwZCRR+atg0rYwGzSm3SndBYX4dwWUWP5dNLn7EfqrNqgy5U84KBaQVRuK/4a56VSX2YAx7
8AGlLCxoXsZXQlwPW4348a3Yj/D0Lf7ujHG448g3KCStUW98ynEqagzuVej8oxnCh2fJy0XPwG64
+lWpu9Jc3WV6HaofwfnFrGTUbsDYcSJOcJaA1DtYFM4p8tZZ7j+Vy2MDC4G6EIX6RnGgyTeT7SCG
dDTtE1aZaUHhzsIZXVuOZxZbhFX8lCTx4gOdmmdBQuOc+sHtDu0MMEJ2jK+M7mz/99D8azMWugXn
DhjtpJ01QS9/DgTWJfheJRw5amj29fbM6LYStH1C/Y3XqcLzNcRlxNYd0jBZ+idl8DxtWua1b/fX
8xKsMwljK0r6gYKVRdMFN8iASZONMU+n0FPlrPW6U6NVmENLnxC3l93T/8zD5jBoi44XQ7HGqlek
KIAQPgnT37dW0LoudcGxSC2MEWkDKXTQj4RDaCAurbsISaykqTWUB1EoJmpkRXtZ+NRUYyc0y7CZ
QsHLmtmtUARM3ini1W/EojdHoBaXda83lKRa6xTvs0M+X0o66Fb3+zpozOMCexK6Xj9YoyMhPnL0
CeoPW7FC7aHztcs7SKIhvKq0Sjnc1X+oOHVJMMKxSc4zoy8qJtj/8qOO00SoFeDRB5uRHWuUvaaI
2jpFXziNNbSRsrCAvrXNGSAkIK9+3cj9mxeUjo2eez5Yd4yzYBeZbh10GKyMlnxlhDvY266Nhjzf
LGPKEVPUjV+bF5DqW5chx/S/mVLmPR9LfChlF8ya8QWY9MsFkF0nzJyCdIlyn8xvyQYei3wgDobq
Fl5hZUmXMWt1G+CctAHOtB3aqkJl869jVGJodVogEY+XApWLuwUlxw26GX3jBY3JXIn6UXrfVSdn
xuHCjoskI+s2zmPRutG7RDAuswCygZ4Io6cc8MaR+uyeHr3iaH6UIhA75EJVRwF32/Me7bGsQECV
8oq7nccTL34nz9y/YPjQR3D5jP4YEsSoHXv9qvKKzgeWowey83eG6Nht1iFnbZp78Po6b8+3qcyW
cCvl2txzIBCG+cRlf6xU1wctWQkC6CT1PTMpW831qMxZiD6poyyRMS7Ilyd00kncbs+m0Tica+uI
/PPCY1bfA7Mt/KDo0/RvCl/gpe8vIoPUF842tN01FuT15uffUYLj5bLwNh3e549KYQfYjtRsxQuL
jj1Mxmk9H7pls95Kz91fbwVOGPWxU/l8Z2Ub51Ckd1oh2r7nMGui2FNOKdwPx5bdX3zfDBIOcqQP
F/7hqGX+MZns0Thn3mlMgFcSre+kqKfztD9Np5DpaUD20F1IkIRAsi08Fy+/MSzVM9ePqxuRdy5H
UKx48521zQcz4hHv99QbPpvALCYJiUORQ+vTwMj/uDg7U08gQ2nafQgFkjqkaXKZtsFqOXuuzPWI
P129SrLL2/cXsG8tRLLjmpd0zwiHSTK+B7QHSPv5XuNAxsVymvTqRs4MtHbkD5Rj7CZUIb4zKSIh
rOmYGG53kTQ4dIA3GFzhb5Y+eS66VaA6x/9jkQNzvHNhmQHCwH1QCf/c5/ckwUtwDg2KzsuJfHAP
AKMyfWS64mPerJRuZXU/2CiZ15asJvYIRJ0HOofrYsJU7H8vHxfKShpBMDd/LBZZsD2FDeNXVbfl
cbX6JX6GKi7Ce7MUJ1EcDMmfolgW3d7Cd90WXvvb9O1FJ26NWgZa2yD8R9c57zbiI/gw//q//LDi
QttPl0cMu01N5I8HdVyEQgBpHubVSb0VscwOMtu1aiwsWMoPBuDmYBZwbzc11X1tcN1SQ3M80d9N
kAFsclyDlEu/uEBA1voLcAdfnTlaWvDW6xBr1Ara1QTv/Soe8h4mowxDliucUq+vrxEc40dwTP0E
tezP4VUgH7+BT6kz7sDZUg+WpeAG7fYvoXhNbbPeNHmzHLIghblVVveLBXo5A0DD17EM+GriD/DW
urjmvweusNh91qIgkg8Z8tnji1kBb5J2DSUpZo4tO1/7XykzSUh4lcdRhwyb3j0kH/NQ9dKeHQfx
LOo+5ArAKwgwNF+mXxQwXzf7JM/wK2cUFKF+/l2mfF7l9TNdTSDrh2Dx1rrZRpDDlk8sitt+KPIF
IYQ2xMKXXnaCWjEeWw7aNHx5zuvM/gadq1EytcM4VUbRtMXyhGuCfvg5RSdngI5/N64KSzUB0mjp
4LFOFh2TGueePhlWsnMW+WqlxIep/L3lbQu+8EcD0xgsq1TKM7HtFC8i8k7ZikHiPAPFI99neDM6
vR9/cJWrkCqQkiyEH6AOcecgO6Uv6wiT8gvU9bE3MhGN2fS3rsJWrsPnX4uj3MeFF9iUMkBAV5p/
wFu0DCo3gXaNY6ltkrgEAy/BgZkDBKTmUKQnUYUH6TmViNAhWROu7lzqBi23dQmLuyBJmTjgJvK6
U38CDwIL7mXedM7d32vnnIbI8yYMp8XvfvCvfHVRgjO1a9/GrPiie2UXtEG5VJLjCzFRUQ5TbIc1
CJyKiSO6xo+1ouKA+Q6iet3P93FoChJMgVswwQliuMPi9IQ+8C+++ohnTe+zRhpVuDlepukhAvyA
l522iBjzcadU4tEPMdH7oAEdHXIjywjaNOcs+1n38AoHEeDUfYdsssp9X65EHm3eJ83vpWhWlCMs
KgAz3/bEQzoWHDz0anpQlhN03RHAHaUqnkhnQ0ZzpsQo9nvpuxBQDtISbR0qXD47OjiKjMoVd966
/gX/xv/E2n/NJtajOp9cOmu1gCVgqKJmnon3FzrGQ7H52B8rV4hhA8JiSKZnrHDJRUi08rVMDT3/
WGPJ7A1/rqRZ6WXglTkQRlPcApglxwaKeEx+nGv5I6TQ062v7IS2hi8yvWh4G+MhQ7qEiMhiABBj
Eowd+oS9WWzRkujQElWYuu356VkkBcxBwx0O05ffCHzrHoYEIO5HQh1VuJZtPoQFCdsRsQj8gPdh
U/hK2m4Htf+CNHGMozmqmwCpctU59kIIvlpCTCWxHr6+8QNwWkb4r7AFWu/VdmdtRnr3VdEVYuIB
OzILq7Kl1FWND61uH1Kp+RBFcNHOSy3om+XyJlNjxdbcLFnlGHIsUOPF2kML3cTtO7UNwYv7Uqrg
gYOritO2yt6U/lXoQThp1GX9FqbofV4NzZCSXYF4ovb0yiVG6TWFeipjpIClcl3cpzKOvIDkoiUQ
TJYwphDT9qje+L4bTP+Pxntg/bwR/5VSigvtHmFLGKxpFv2+GyG06cA5Dysqh0TAQPHocUw6rvwZ
0Cd7sDpqq5RbUejRFY690I2ctL3J/rtD9Wqi66YiFYUpy55f+dxnUGpt6rR99fPewIGh/JST8p/k
Om3YlCTpn78Z7bDzzVTp+dr4QpUHcxsW/vlaCSM7fVSZo8KKYely3hsQux9oMaN0YIVFdVvIdsxo
YseKoFWOejE31MvbBz+EwyJV6Rwmle1wUmSi7y8mbiUFmQ5bYyLdiYNZJa9bddtEnoX2pz3KW+Xm
4EqKkseD7fSCK9VdttKb2atSXNtYdigB+WKrYI2QVcg4DpR8VZzn3Wng5Efngpb03lJdTlUIwNiT
JXGAkaYfEUdQE3twn4FCN4ztgwpE9uPpaqse2my7YhXVv5/nfrz3Y+Pl0tlvBXvZHLj9iVwLqYQP
tLDyzRSpyaMaXd+9HqPLmCh2ySxD5u+vglCHvGv7AZwz7gXb1MY4e4dfSnrqJaGXHwmbonkiws0I
cDL7Z53flnXn2sK7sdZMYmRwDw76Sv3E3txPKhXSR61+requoiu0BeLwBwvzltqLbOD5TDnPPI3G
mwjKyVnj78L24gbMu3kpei0tEaUuZclm/yLfytAB3gmMfLkXWBH/RQu7JYbgiIqSkWM89vGhCf0G
SOGEIO57P58teYpW7K9akHeN8IK0SeL2Q1NrelgEI7H+ep0OVtENJs48OFQgRsxAFN2oVsgEDLGc
3j+wzess2s59DZANnXhR5EgxzreklhphU2hvnf9iifjH3IOKVyWda1WJR44gp9EmagdeGsrQY3VF
xjfinTbVENjS2u4mTf3x58gal0kCrGFecAlB+B1vez4MivwJLx1U5xxTM37qxlDgRDm3X8ZjICK0
TX43zuTG/oECThazpkvkkCQbMd6g+Vg8FqYAd1maFLVZgVXB/1aNaD7XSLbPHyS8wq9XRtz2pFkI
KFfmXpVr6yVZd2b8cTwIoVI5AtuC+vboFsvnTcfN3MLkA3Jp9UFNU3hF04O7Mw2mS/1hGwV5AQR6
r060RW6FJ0rwXB6TJKanGyPqul1N7AtRTMlaWKK2UaARscXcamm+Cg4O8DzAnjoEP+vBmFLaVmkh
r+Y9fSgLKi22ANDpRXU6roDTgOfPUsoxra6wsQRjtMYGkHObViNH5XBIa8zq0EhfOJAiZiazdkPv
SE36XbCqMncpARA38zQE2Lt6GmOm3ThFnWaIHe5c9f2GtYlMPBHuxUUHBdY0A+CbcnKaSzEL1H42
yYh+XBlntho6nC/ZDXk/DTbuycM/GN9zYCE8xXTlhfkFqsNFaP9jkjKn81Ks6bKm8U5nIoOEWUXG
fKsB5ItRIu5lV2ttatYeDe2BSuuM5nWkfi86OnvO7CiG40oJg06vNq4L/Eh3epRI/A3X/GNE6Z1h
At6T+p5rR09M5xHFEqISsW81ivr0i+Trw3oQ/tYnUiyMan2XzIo9Ka5JAQihWS/W5Quz41x8GYP9
aDOpbCLh5ONk5Ak0mW1YAOQo3Sjs/sW+8wXl+POPt0asXmzrO7ECaLwt62+ccjYNhGVSmxDgQ3rD
U6s3f94MJm//821r/TMGO++m1ijOmz5fsjO6fv9nXKmDLdrEyEHy2foSLgnSW3P0n5qLC4E3SEkq
El2UR84s87Ot7RC2MQfx+oSdhqiS5A2qD/yEMtAFkw8asrKVem6B7DG6SQ5S0Y8lGMJ/uDZwY63/
XUMI8pu9b94lNEFYGnOY8MJa0z+yWMrzWg2bIaVd8O2+UUhIsWrDQdfncDxjQb3vlGTQfPDUWQks
a5hTP0bMsr1umnLrIHiP/JEQcFkx+e8BXTFwahmaQ3dW6vq2516TicxFOEkb3UAsJswd8sOzx2MV
3g6CX+ns335+o8wvvYxp2Y/evAaGqNqJOw88EIQEtDFQUUPsvllAQu1mnfizy6q1dT05tTjUudr3
42k5XTNg+QAwtA4aUcq2APIRZ/hwucWft356bpzHbhtK6bJS4Lqxfio9vsLrKRfVyFuPIXzvaAAO
BVD9V9sdaTe3nPmBz8fvNuETy+QTMmdAEMMAP7OuRtuXimlZ6aS1Jtju7d3zlOWA7f7dtwyMxQag
gPWaGp9LPFuPWafkxYrQD7SVhQAjF25Iq0XN8XhBLJ4fmH94owZTlKNpdSLt5FKbQwPZ4wYTQ8TJ
4ev23Dmic7+wdn+Q6U40PMAgjTzynqMTow8zSK787vqN0nS9jE2j32gaWaCsjYZa+2gvwq5TZ6pF
uW6XPROIXQzwkJdZVsGYi1ZCyvgwY2nDqaQxTF3uQTDRy/6A9g6Iia8tPVie7QPhCflenW4QFkf2
eeAGHz5yW9oOSMYBQcazA23FRvCT3SkoYAe/skWiAYDCn3pH0vHo0LvZyNJKXMu8WoMDuvv32WNq
IF4dK4sc7jmR9iETUsm+8bJQYtVZh4cvHJFp2bStzqNnR0wRnN6LNlBOF6Rn6ew9eJ07BbY+ngSe
RX1T95KkKJ6wmVyqgukmfqWCdXcTlpYJ4LT9VYRl6xal4mYHu6fAU+gOBbg49iYMcomAqHvs2raI
COof/rSfXVmQfSXgeQSPWYlzW5l8x7gf55gtvO6W+cWoRAMlKUJCijHWgHofnwD2Ts0T/RihpZQF
HjeFcGBXhVaIYquYSH4HjRekilsmorTbPzjbyZiFTqrztw7G/QAS8+x56a8/SncRZCJWJCEKjpJ+
9RqsMrMuXm5jKeSVCrOuMWFS+zh+QK4DwT7YhJ77yHUXewF1l5B/Btw0WmJLkweWA/aihJAFGR56
/yiO107jnkqmVBO/HQzcM0sO70wqeq0JFBV70EOPnRoDy0FYhsGgLMHQmhY0nxsET5h1UEpuHeIQ
FRtheFeVhkHwvAmROz8GavjpIA5BnJWEQO7CEQAyzo/PPVOGhXuoa4AX6Z4db3UD6YSKJ/e3lgaI
alBxOmpnkAyXWzIdDDsU4WaN4UEvKV8djBR3iwYIO39d11ilsk+crLuoPjNBOTgk/+BcyeKfZZC3
TUoNEj8H5gUDgk2h7ZuOw5yxMGkIlfpsyTvhV2R3zL/srpUhrL3jATWZEMBw6+5p5QPmId0BizTn
WZ7DEB+YkZtgU/mW4jO31soE2cOyLqD+oX5C282IYqVi900o4XDb+GPVFr/3b6oFLkdKbeX32i9z
yKUrZfxOJk+JHJcf/dX/lCmYNdPrYH4FF5ns4jTzUpKMD6G43kTghrqaMEZyBHPMdJ7jFNwiJ6kC
uI4kbDP/TaPP1HI1Yo8Nl8AFzNYXZ3pueaZaVATm4bv/YWcVWLqsNuSEfiytz2v0kevZObw33GWp
u3QH1zYn2OTsh8a22abIL5sUyQuj3huq/PLSLoW2PiN4ZV89HOn3XfyJC9lMX2uBdj0Ksm2jSkmv
qSyYQJHoIEoyN4Z0BhcYI77eo9cytlq1jcDKYSDKHvlpXIU9ktINiEzCHLFlfRXgrjvvRekc23pj
+7K45z8ffr8gyihCgAQrrpnEmK36P+k7hvEiYs907b2HCXl1Fk7w9OoeTbn2BcdLnubxf2uEzbJI
jAuRl7PvaUTG6ptbX0t0kg5kIFaD/lopQcL4Nv1S+gmy/oIYx/7RjxDIWW1Ytl1uAl9EfB76Af18
KQ1IAzMxS13elXI6IELYMFb0SYpzbC3xNBFguuX/4QT6Lig9pVk4TQctPMERvzahuAwEC83wDCnj
wyCh4xbi0cbeRPFC0KH9TtYUAFjSwkoMc8UzbJk1LSeVPJ4utx7NfeU9IkPtIX+zwLk+PYsGAzs+
DffMEGU1d1fVoRlWaXtrOvVF7H0fIUTGPlSeempRRzFx52d3yHMjOgh/ZoTmVQPz0BXfQ6Gu+hqn
oJhmbOESDBoRFScwCpuXicL+YVeYFgUwxPEMgHEG+Obyfq2+C3XqwPoB3R+ZoDFMAZZra86BQnU3
o0Z2XDuxPkGXWyFNqoyX98onK1bPc150lKxb9NudpQ44g4ZtAuEDGUFr9zrXVJXJM1WYM3LEDDS0
XkAVInWqTbxSs27TiL418pBT4cgRR4tF6jxogGQeUkGvyoWfkw76FEl3MC0MCvS3/VsuQRa/oKIa
YkceNsxK6Fi9qWjFaMw7vu6tZQDM+6D60/GTICCUHl1OW0zcqNIcAkuN20h2GIimZ8PwnxGuXOIg
P63N9VVziEot4vlu1d5peJGwkWO2aHNd9o6ZhRS8QRF9lRnrPKIRr1sWps1PtXQaQN1k1B8F0isM
ds/nTrvqI9q0QWn6QcWhZdUU8YaeON1Y28tiFubChTR3SpxOWbSjdQ86Mk0RmYv5JExZP4JglWWT
fr5dzxH8vNeMzNW4xJzKiDpnRBNarXWFVHhpzzbFxCe5XkJyrOgYXISZ9bp34ggozLwr2v5AcThM
52hwINCw7b10SeVhIUJMTsf2MJNZLl1A5nOadQpV5vwGpl1hgOsgqwGvfit7Q4wwXmQvL6jeIxWh
uyNK27/3j/d/lETdEnW2hGzbmXOMXb1gZGLTOCB75H36MwbzjjjQx9ODVDBLLhgF8/jp608IJz64
mnkIJjD71OTQiWFGYuWHCEbu2SMJ/stbH9eG8LA1iEDgYM96TTdcJua7CxmlufgMfpzPXkIta566
sAVzp5fCUIwKAPs8WyFFI3dhWQASX8iMH03/uruOi/oOKPCY4hiJtFY1W6Vs77TmpX+DAPjyaW8I
9K/hCHzZZbsh0ThCEUKLljdg4N0bBsYZ6/jr26MbjH64ocFatm7kQtb4YMoTEwZ7q2m7rPbRNuuW
MfLTmgfPbusMwKIVZ5TduQ+yJiRN+wn/H0b+WUTICov16pxcuaq/yuJjuNdSmNxjRkdZJ6yKWfu/
Ro03ZX5mgSbbAmrUTXzd8RHS5FOILEaABZOoodHOTiGa747B5LPq6j59v3kBWMvl4V4Y1Eq6MNx9
WKXdUbynhJxDFfORSK13tP1zh8Os7eEMKFeScCuSoN4UJLS/nTr23hkG+8Y8XYoD+oEoo5vRlVpB
joHvlbvZ41MvGybwvPm1ZMIKUpSTAXYnoTlbq2PoC8lUq95HHZoZjuJUwOViC9TX9yZQcdar9mAV
WTBbnzPUgwX5KQ2E9MMcIzUnS9yMWHZiaki9Q31o3ugklF+vf/JKHWpipwl/FmOl0SYRL+NJBLgA
LE420KZuw3IKzWOGEjpeCx/nJuyJco5OHp+00ClJf3yPkLlrRkLzXrE2O6EZwGKihxPkcXzvFams
hPisHGV+RmXQDlIo57FAkFr9PeY4XPTUYkQvSZ4g0A7j3umcGPdRK46dTp6tTR18omJ1eBGWdriT
xHtXthEyJrJI4CYEVVoqqQaONReII2bqaa+rZmFUJDm+2Gjvfb8b4n3ZPlTV7V/02jvOPu8m9DOi
673602w/EXFLcUt1ggKv5U9D2YG9Zq50Iki0IHgWE5tuYV1Bs8vo1beEe0dwoknNR2+prbC17NlF
sI6Y53LIyLnOH/JiUPCtmcRYaKOmdY5fFDsSA5zGzDtr5tlULQYcyfbyg2c++hUr0YqQSzyyN1jS
GmfF4E5SqZvzIw0ccvB0zuTU8P1BqVPA3hz4mE1653hStTlcZuVp21U3cVYZBKlEwA1sFnerWliQ
DP3xvtGOa5qHmhOkTFlmlYWPfS837VroLL5Nh/Nrcb3ffTXSJi/mzh8h8VXJn6BY+VAdVmKU9S+I
+DedWtPu+X7bI6jvdcnIjRR+6dQh4EyZlynm5PGE4EhFDlPAcZ9g/WE6L2bvus1xnA3rk11MmqYm
JJYhj8lrapPHdxFfWk17E03xp7ptUGfjosEDT4U0BEj5jFVRhigovY946hy0VAvqy+24EsJYFf5q
3UlsXVTL1BQvI6HUaRxwJjDL0Y/NNE9lwgQmrapNoTgDnBQycMazEIzuPCB48M312f9HxkexvEGa
UsLQkrsI9/CvM9FEm+VlRasI3ARh2J4j/g+VNWf2Cv1/btZ6tcVQkivk/SXiKpYzUeFyAbUZC8Eg
emL0pNAepyT1L8Lfl/5gl4oSwLXZ/UxZvfazoptEwUsBuVnATLPYKfblkNRJlY1JDCAjzgEaKzHR
juZxWPWuljp30aur0rxjOzyxmdT3PsU/tMCqPW5hYmOpnCkvQDE/t5kXYEMXsJrscWSZu/1pdBhf
Hxoin797fbO9xb3kuSiMABoBbYRGv/RvJe/oBkJ2upw6hpWgrMIGPKecMFUFcjuno6Nmi6vamWFG
cjKNASFNByjCMdM2DzVicgxKuOOxiPtMD3+4lS3wcBy3z+P2ckmoYg6M4dEHLEi+m5MRJPjNwpDT
KCguaj3RhKTEAmYkxa+W484IcM6ZFk5cVMS7Uhs3YI0O7nnXl559prAqZjUSZjyLZvuxnGxpHY5d
4QBPHqdixnUPax3f+bksd63bnK0YNkclVxVcpraPumbgpR50QOJbayos/h/0JmRgXD2TZpYalBtH
5KDDleRZV6+T7HkXQ1ReCEmpeJQQdVKGWf3L6d6qDXC6mpTk47IX0WGC7VzOjwB0s9zpxgZ3sskV
5eUqYTndTG9+vDxZteQz3loa4ncN0tCnRAmVXKF5pZXIhSxBpQOPXf7xdALu02IjzaP8TCetb9Vm
Y1AnctdUce7abYBMqQua0Tye+UJgqSd7U9dVz54454Ru6GMgWjCv3I2VkMFSlOIErskuW5+XoJQp
7Rqe8OeNxGxcmBVjEEek3zdg5GKgX0QmQWcO/vrP2iVtQFgLsTjeLSy9lwQDSnE/SEX0PHU8q+MM
0hEpKaVuA/6ITULTZqLgsxzERuGF7PnR/sk9dVHyyK5jBQqlr1Y+wl/FwrTSouPFRE3ZhbqMpQmf
UkXkvWhj+IPMaa9E35/Fxx6TaB+KX4hgc5fxcspvLuAl7GJUv7AbrV2DQNHpKGQ90ubU0XZn1ygo
baOFpKcnl7JwtpEvsp0eNhuyKo2fmwSIbGRQfVkgw+EtPcpzl38GSa6zyiDxHkcyeHHoLshabLNx
w2pEK6NmaqgzHmXiOyFPauf1gcT2Z6Yp+vhmHBMOk6qY/4z3UjjtdkkHzmqc1uhk7wnAXFqnT6Z3
UnpWFvtsgJomXE8d7SckAT1HsQJw/JhUH6zujUr0wjlyK+1yx+GUHY8RVinUomVh0f9+GA6c8m67
6DYcBEpe39c2NZiHXMIaQ081MNJr9asEX8aKA+vXc52rAInGricsgQ+0D3j4hma+93MjA2DMSeWn
vUe58LEj0rLRx8/UxZ76k2y4C+LoW4/QzOGVtRdOyu9kxWo5G4bNuWvLeEcuCH8nxNdPmOT6/mxY
AwW8KgDukDdkCx2ZhFq4jaSUQLfCTVfDai0IFH64XkM5xIPw81i8EjLE+AZy2vxqVmrQEBUYabFJ
oPUpyihJGZTMML9ZhG0nkwBxwcYaMi302T8ssyC00DxWubr26dXtQG4CTMV3p3m94whtXQGHOlKD
9hvIaKyeeomtME/nIZWo9+7sfkelRP5vTFhXYS+F+SPVvjE8wpZiStPaBIB2jH6MSJffTV7toqQZ
Dup13dE+aOHOQ9Lw9AY/xDXFpas5GOCCNv5m0wO3W95G580gAen4ZDvZ+GjFlIvat2dwrR/JB3jb
usPdJQ4Q8HKYrnzJM5932PS0VBDE0ZIV5rV53v6dnb3ec+G4d2UWEY0eESQPVL+ciw+BaCi+HkGP
FTKIa3KK0QMx/LSIo/KtKLWFzMCTckWN67+NdM7hq/G2ykKxK7lPh6RpyqWLtYt8aLRN9rJIEUCQ
aYNq6W+K8T6spgk7KJL1pfJ3AHkQfkNtMBVzssgByPnxMJZta3Y4housU919pc2BXxJTcYcEInoV
9v4wu7qSXQMTcakWERAvWmt3eHWa3LNZSxWtwmxA2jxnsKi7VkyxsfzJny361q+omqOUsQf7vK3A
5NsoYTeGGbUgpphPy/fZ95QO6tCLVdnbsnuSWBQbhhF8AxB9ORtY7Ctx13LkdZl5iFnvk3o4hk4W
j8sRkr60PkqOX+IW+3DT4fiHj2SziCOFooNVa4qZnFRWyIJHiez19xLNSTnVqZPMvsBeuP2Ki9O4
xR2A9/7Ckjv4cDwRdDZB/o/6o7pjlaeVUhDVigoOewP7bbIoeu+bd+72USo8RsVCsxNn8HRorYEC
OMZ8iR+TdQ4NEYimyeYqqjeQLDOHBfhcSTV0AoGckB6ftqi5gKDTGSfqkM74ddhRc/Tdt2eCE4U6
hs7RwAae6RHgOzYk6Ymd5NKjrDx4Ui9qBEJbC3MCMBJrhAvEFEoS6Gpv6/+tReWMXwGd+w6uELFM
VsANUD9+fueKhpOLvEUyvB2beE/HKotIpQa1ouLrI6qMykUi3LOgssoBdRBCDJPKnmyasB+pnTLi
p2a/7QAX5qlgyt+MhyBNeqKeGxQXvVYgaJ+OSpzQMime/5znu1uVmSV//2sj0++tHpGgM8yctr6t
J/59HZ3nQuzafBuueCeIwhhc6HGMWzf5jb9iEb+KMzYLJ2Ur0PqLu7oS/vSlM+fq2sDtZeuTfTz+
kaU1DRIWY9djbmqUzrmeozj4ibjmkT2bgcjlodb1PySszb/jXYPun5BzPmTbw2EZY9jO5S+YSKlA
I3mLaCHz9E920+12dCBSeMaxX3RDbeynUEpRgdwp316Zpuos4i4SwAD267BBzY8ITmsZBcWZv0cd
uZeVeXCIdxXrdLjNMQ4qkSv0eiz60Tiz8NQdEm0/dW29Fg3Uuloenrx3mHRUQ+qV4sEAzqf9zq58
La9RT8SP5YIaDRweI6lxGiFn17zd63DBDXH6cznj1ewqZ1TXl515doTaSeCDl6JY3MRam6sycu8Q
juYyyncyqE2sT/jY/Le7GVe0sL+Jac+UE6Jg/72uMWcRg1oHovWPvwPMTDvCp0lBQY6pdNTKehty
+1fD1w4LFG96+MCsYUWym9y9OsqgmEZwKSuZQpMSXwYk6GFSPsJJPSFI/Clg5MiO7j9ogr4cYc/J
kWv8Zgtbyavj3igucNZxsbrUayjtdxa8YYlPSGVM1nyk4mSAM5JWy/3Fx+Dwgv/e1jJ63lS3eHbo
jQaleaAycyTRaWoFux/ecbQehDHZ9Od5B4gRdMnufS8kzq9YJ0lzdIuAC+SuRbNgIlJAaKOF1Du8
x7DzX8lczBQjpqPIgD0KZYSoz5c2PnNoHQFTnB0RL7vGsOmNodSJqk6MtxV4MI883o94CPHOTaQ3
XZWKPLDq91xdfW9JZvS6122x+VPaEI1FhAdlj95WV1DF0IHRKKRUctHGKqIN9k5FVme1JHdHv1Ic
wd3WPVbGvZ8Deg7bFRU8DhPRsFF5N6Ypw4QpePGbSkSBhiQg9h3O+DHI3qlvIDhULo59BrhfQbLt
KEWMqbTqY2PxPkvu65R/Nk6p9i3sVxza2blz6cGaabRwlT4GQRVEu7FBVRNsP0UcWTTZQiqv2gsY
fQZvqBqNFKB/mRHDz/HCRf1Z02tiOeAs+C5cXsr5aXrxKqwfEsPP2rh5w6bF0sKdn3+E5saiyeGD
QQRD2QmqRGdT67pBDegq8R9l5hauQBEk6pMxYIqvGS41qeybODSU1woj06PRjAIX3NGklCpoeycM
7dSDr9MUdnxB08hMErryugmvfo19lrRfd/YpXIEmco65rg820+mr1TPX2TmQQ6xMqVgP78g3X7lH
7f0n5e6zsu/zsmxAr8eps2NG6blnHEQ5CDpiTwMPCT4iqSdvMOAeDVNSWkEVn19UEEhGsIE1a0N4
iqqIagB6Zrro1IBtb4l0Jg3rE0bh0yvtJTF7JBG9Vq2dOpbElFUtevHYL/b3EJVSUWoO8W6rCM7t
+nujqhhuxt+OKb5CiN/A8g/lMhShXzIUF9jp+w2rw6XCZ4bhdzdjSW7GpdBU6AmVQN7AhIiVr0KV
AoUKyKUE1C+7EJDAKV8QNt8j0/bv+Va3HV1b0IwHYTYOyE0Y9X61T7S5QnZ7THj1yVo1jZK/yWKs
dacyT1kQ7AiiNaCuxRFLDH5K4TKlx4dcjC2VmLk3YYfGdBLv4/KYH61iBaNjaRCa94DVhltI1eGO
W72IO+zImxwuMEJEharEhStZ8fRydgdPW3BXSMr657ipPk88B/nooan3qABascGaKoJwID+9NOs/
dJOY+q7KT9RmZ8ziIrnSyRpSJYrUpuS9vwHrGze8HavtfJKhcQwoetv83XtPPCPx6h14ICHwk6Un
0wrvX2KwcVAZpD+n6WPPGmdeAoKAD86mXWszHQRgd+TxjcPyNgTUbVogQ6l6PBM9E4rpYEOJ5qap
nz4TGZnQa1ujqmChghHazZXqtrDd9W9sOSh78DxY1SZpOO0+YFVRNTgqxFuBV8J5GU6akkcjKBrJ
xnrmS6tHckOiRyE56AgSDT6VyBxd6bNgjC4DtC4wwcuIbIK0CWCOZBK00wgxWQ7k0HIh74S98yLc
zwUADy/38U3sWWwkCHdxwKCAl6i5tTWKa1HwYnyjXXWO6wQNRH8pXLtzeNGiyreyF+wQtHN4zDKj
QJdks5yuTVTMBPJVliIxZ70NvzceuAbi8n3dsQnU5Rbx2doRlxHsxVXSrFPVDRcCYs3Q8sNNUBj/
8hraNkCuTbHGMnu+KuZ1xah76D9Vu9JYoo7qo1zY+MbcnlwoA/3bGbCWDVvkQoD6Obu6SDhloTeh
j9T4hsoPd+ueWIZEvOEQ1h3akMzPmelETmEBDF+4mSbgQmXgO9mZCeSzZjUNtyr37MYthjB8kIsy
yuery43hHB7DByLljbKMa6mf3zzG9zNmqumXQrOq7v0JBojxCVHHfezmZ256/UsfQw5MNDBx/TC1
e4rzGGHwXwwQHHubYdQp2xuJ6oXDbfk0Ra6EMwc0bGiU19nTHzxwLhRL2aTR1Xk06j5Vm3uwZGuv
rm5dD/OAoI4vaQ0cbP2kxpiAvXW9rZt/3A4RNDkCz4kcqK9+hlnVviBOfA3mvwnQzhAlvk0hn6ku
eJz5B3QzfJ+hymG6tldJnj+DXWvXx5r9ok1HyOK8zoSSWU9ncVGiVifwXlbHdvYXHqrs3wSVkErH
GLu3phmNCl1q4qs4hDd6OEyb7BBsKgdeue/cqvzZFY6rWBVWdAMVz7immw3wdbStAZGM3wV2Cj/N
sePJ06yn3nd9V/FLddEDS2jo0byn5OhW2tzMZ+WAx+d7Mu9xOV0swEsMdE4nzkmDReFSGkGJFyZk
mmqZz4DDOtbfPHzIuTYv61CL00Bk1BPD0gqFptqLU90QRabzqJM8Yfgm239ft2yHmYekoBJPhXdF
aezF3BAios8f1fJhHqfI4EvEeiEWhjDJy/TqawJWmYeDuG9prZ+V+/6wvGjflrNRNrI83FEyjgmP
tbaay+l1rpXODIOz/gV4kyL00xJeLMBn1m1xNqkDIYGEScK0Ogm+XMlN0YR9uBJXXsWn7XlNkWRQ
yn3n77bxhm6g7XReKgSatRLrqlRFNDgvUDeUVUxLsoTA2t+ai0q1RWc4yByrGCWRzAYw1PUaGYub
XC5TglMpomdv/LTHsSmZ6i77B39ghruvAKQhUp/lVXAHgIM+G+7WPVLZnCvZXCUI7WCEeOX+e5OA
8GeJLNRqVRawD6N+2+B8Wa2g/OvhZpd3pHbotgHkuYJalxnwIOubELXtj7hV7p9oftuteY+V8mkL
1R95isvoUuvIfHUC/WESTgoAHDjFIXxDI7PWQ9Wu+tBsZYRww8qJ9dVnuRqK54gCLlrIswwe6uBa
nfz2ElHx6K9o8vG0gYk6Cyd/nrbiyYCHtfEvQU8zwAh7XzD9bz4F+mUcdn6VroIyJmiIjo36+inv
sCRCY/C9PrGHypcMXI/6t822n0ELoyd0Vh0UZkyYOZm5i57RB8FJYpu0lM6T/a/HkCaI/v6fui1y
DUsq6hmiSzE8uhCZlM8NF+o81Fd2XrotwP4PQiVQx+UWtuH7UqXjnxAvf/2zYPtylwkaNABf5p2f
pa5WMOh4rM+wk5xGRYXurdTTkCIEOzomlK2bmFj2JQB2udd1+04LpSTRC/6fh1Es7ZEdulHmcJ+p
8RUdcF5uiSLmfi6TV/a2pTlyH1imMVZyICsRxCKOlmhdYw039syJes7a8te1amxYpdVpsWr7jW9M
PlzJVRfJumgo7fwIDQB4m/ZapmLkz1GzD2j5Gb6iwWKF24VPdxXLlWzbVn4AaOE4KzrD/IwBPkUr
7webjRRPtrzzvsQqQqHjaMRtu2rGu8HE6EWeiwF6sS+pF8xCkiC1OZnq5HF0CAyDSAqvT1LxDtB8
JA29qKS28aM0fHa+qkMf0tUVNmM/N+NnDuNfi85egmw9cswlcHT3YnKx+Pmklv1ohkQr6D+us1IT
0d7gDzSOPvQUF3sI5twBURVuWBiAMNMtA5kyZ6E7b+BLBLzqxc0gr2P30tCLMiwcLsbn8pm9cj9f
TDyonxZmTKM8PHGmWNbISZGr3wrdy6o2lQ4uiQPWnioZAkJBUcovzDH+38tJ0whSwZq4AOgNTJk5
7TNfjwSb6ff0+dWE+bcKY3Q4Rbnrof5h+E3UuhQhJZGp7a9zoUiO90TQxnivc7Bnd0n2FD+oC5H8
wzj/vUYUD5P33+mFJdD2hS77Lb5gIVXak9y4cjg22nT0+P5c/ucIU64XsWD3HTfRUCPBoaGOl7EH
oIp+NcvRJVkr5UjetN4dfEPRsK5aNXHWpO2dWFIr/wHDJQgmVFGaz056yvUBCm1Ni2GworPb7yNO
S5yFtfMqOnxsIk2r6lrXLMmDaeg8YOrkHxO4aA4ygMPAz1i6e5lgE0rkn+5iZbrQNVvFSkB8bZIQ
ei/9EPZkLDhOIpaDOD8fOd0woRW7Roqn9IGjgVGaw6ZzJmlyLuTM19l6mKnKWQSIc4wJ+F+RHwUu
wemuC0UMF8yv3OhGCXdASvbb6HlAu3yvUUSZp5sXIgkS8ROsY+1fQvXLgmVL+J91QzcmFHxkDgo9
vRW5fxkY35RrrSq3vTxQomLS3VCH8h0KBmoY299Ei4SGkaN6PQr56UgLJTHI/9VC0mk4LVcjypkk
OU97rHeYrZetw1xLKamasoYiHQR+sVHi4dGVsecIqzm88nkKKfJN0yC4dly/fqsb5lLtAYq7p8KQ
9Xsw16X42Hp5/Zl9hiwanFvQz80aADLQm7pef4XHYOZ5qa/1QfF30aTDk4ticSD4ZruQGiGZpM3A
4MobdDLmtPIziBpwlesou3xOYhbxW5AI7jTHr9fVqUhvMCBIDUFgr1i0lg1as0n1uom5khIhiXCr
+BNBpMkfNMDhnCaCkDMNjA9AWbwcsvpGiCU7LCGGjCth1W1kiFMKhwm1cgxZ1PDbP0cGps5VoFbz
XGTe0wAAudSCBbz63HB5bDsi81aS0fJGCXLxUsOevAaGlwFpPQ30rfkXaRoHgKRvkEo6YM4fWBtf
+iCIAMxrwwzyZ5en+bbdByqRhpsWmqn5NiIQGO8cSjuce6x+lb9fs2JjjIvwi/ud17LKNXQcnSZU
YqwAxJkOE91eVdbmwJopcQY4JzKn3PHt9XKHz4Kf7u2UH7TuDHUE1mU+bbY+U1/4ipDTCZYKp/r7
2kyWJH1Xg02ABZZT4sCFcWZXQ2PkdCl20OGbkPnE6T5uZVXv/e/B9Oo8lmuWq9gbCSMgbDY2P43+
Ks+o7bcWGefCfIXAIp4pU/ofjwbY3AI+JEG23NS1MT4x9Cqo6AtvlY/fekmwNuJe/N9k0+NmMU43
S8xT7hXxhUWVJB8hYm/grSUgPTmUqjisQBHQwE8RhSgcFKJIZ8wHX8cDZVt1Sx7/G3qir0wuhbf4
aMigA5bPXvesWEHnIuRFyLoddxI7DUxxwhG34+CpD+UPb01v7QN6bqDhO/Paybxr/f+yCYB6GIWn
Bv0HFMfi87/benEoSAzr87igwiBbLQ7dLoOOBBtOKc76KCNjixgtsP+JHDIQZXpPSyfsJFV0rg4F
BV4dDFc9F1PPc9Hr4Uzuie3xm06pQvvnrQ6shr8AjX6Dz1iqeJtUdtqWY9vOa9X/pv9ZIUqrSvpx
vOncvp3XRKXvahYRO8k/72yXfDFuHESqxeJPPOaVLCoHoxw2sp8QLjirui7AFD9eAcKpIgZom1/f
64t38AWiJdf4Tcu37RqhIAkfMuhYF/hUQoHtaOa6hokp7amtNCkIqF6ILD3tTiHkd8K2tV4p1CLR
BoKRVz+JCg5U6IxOPRtnb2DTzK/oHWQDWdMk5Sa8AbaVJNi+ZyXwj7I/P9w9ty9G9FTED25x6DEM
FqnpXaxcZzKtUQF1hR9+fRiHp/KxqMSD/5oyXfFb8NnwelAd/Fk/Upbq0XxM37Vj/vv0NKNGz3RF
rnw/w5XhE8ALxTYjaLOzYT05nAP9y6VwtEf2IWi3I2ir/Ml6T57tX9dUbSbrTrbAv7s2Sccr41fp
tTgl4ABBlA23VkzUvB9I67qbMQl7h7Xvbcsz1yfg54azAp6JKNTV9XGGlkEWtyVBeEKLkRmyt2Yy
2dgzeNB4xpmZt0Ka13ldqLlKzhk7NzXQxH3cPZjUSUXwr3jb2vufM2U0pkGk9TqJJ7fKhxTOmo6w
Z4g8HoNITW3gW8/LPX1kzySurJysIPo5zHsIbk8ms0WbJUrCQR0GLo7nEhp4R25jwl62eEdrZLCE
9PTwdHWbFsqAzpbAu9fRRe0xHXdwbiKmcuq9+zLYSJb315IuZ5hDvnwGBchxGrkwPm4nMHUjqQDU
x+p3bxsLWi8qMmISCdIRDGIdLPSb2/D3yyZLTZ335rEa+HB9Z1Ic/E+S/yKOdFKTAWjebvY1ZWA7
kbFC4qQMiaOyjDkbKUHwnaVU0BNni3vPLbbKzkIPoT4P2MFg5wxooxmUDmx7CmWo9EV97LLnTc3x
WDa/hYQtV43x/ddMlfBOvQNdoJX4+wG8GJYHUHsTFjKcbPjZwmb2XaifQsZNz4kzRuaDGAbYBzFn
LAUbpre5Z1qEfSD/IQboQGO99yzDFghThlmt0xelb+SXJiWj8JcvmpjZ9dfj2z38nDE7u0JZUhuf
hRUOSSSNEvKFUDUaUhCfWd9L8MAeTezhDjN5C1NHhlhV6ox0tlsy+ks/j8y/km02kS1k08rrc/TM
Nq3K0r0Mz4Xvz/M9vpMSoohQZBWeLFkZLDfyPOcbjbvIMAZq6ZVOxPpSfp9+wGqkyFD3nUIuMLaq
k7N/h9OtNKWKinn/Ua2v583KzteypxtI5qIWuakj1pSXBqtpCA0++RYQoHCpBeHYfvYPj/dFZTkv
+tt+xZF5yF3dgL7cITcp9ezJXHNiK4oZvpEFBr6ujfJ5c/zDlOZb5ed/jSulwADyRHna9+31B6Xq
ll0prbATb0j2tXDcwg6a8pvqHr+zYoGm/bbulhb7GrYteuXsqvBVVZxQmBfpZWXCKGLeLETabfTc
LqfTVT0gt+PPlfadAq/0n0ZJ3n6wF8+UEqEWQyPX9PyIfEUz54cOz+y/LEqqRXMSfy7uGuZqHbp3
EP6v12NBapzinjzs7VmNsFe9zE9vqwVTdIDY9DZPCPldaPiG9MulHuFgpbvQQmdPcv8UqTIbW86r
ewv0m1SeRNo4FnA3Pxoruj3FIx7LLn1qGI8CuNu/6CKXjt0UqLhATYIWiGHRjojt/WTyfMFV6U87
gA4SCtMJlBg9CbzX3TW8fz91Xf4HSWUYNVHkVpalMgcl0odcyncAznFi42YHRoEA8c00YKD8RjrV
QcBYat4HQ3eATBjiKXZ/lq8qpbAUqfYGo3jKJYvBOuBLP6K62fDaFtFdI7TRlTTPwYnk/0c+IpMa
SxxMpjcYntopHqxcnm+wjz3sw3pqaUqWPyTDFmgGECZr/NsiGHspaCs53YzxRbe503/zuRv5cxSd
lSov+bXEzLDIeKbX+Kdntj8yOjEvK9UeyZvQi3dyGadnF855tvyju1Jx4coi7ZyQHflh2Gw1zwzo
IS0szHKlQ2zqMbN5YV11t8urgTkZkU8zIHk13dCaCzpUFPAowVY9SC00KylGNLjHx5aNVSm5O/tZ
JJ82nrnDrvsWB74ZnAG7x5j/bKqjobVtAz7jn86RpaqgiirwZpCx0jKvZ7CQG55TNi3fHjkRWTZ7
PsP7iewq984hSXF3WZhmyqT9uPAGrzo2C4IfBUhncddKPaYJLIynhO1ws2eYCW3GXiVx6oUqFnIv
mYRSJddBnYwNPSBnPTNXmM6PQjnozVCafqr8NnimyVR6WSc+nWYwBzGGf1PCRNxRaO168p3iGtea
ZjPkxe34yJ5pwVeOc9eEMwT8OVCAF5ROTu22JAC7bVcUPsJYwhijqr08BSsxv8vP0QaR3eXPgneq
d7m4jxfvUhEFNx9ED5g1uLAXoDh7eSutkzI5Yz/QCQ7KnuG3EUJ8kIdXqmh+9B/slpMhfbjNBAyu
+gNfdDtFPHbX1c+QJhV7+udtjUB444fcC75HOZN3cqCljKwEDMPgOxd2g6ype7KvBV+9nlmB8VKA
HJKAGYWyIxmNsXd5WF1ADSjWV249MDmHfR/w6aBPeP9qTOdZ4jK5OS7DcQsa9IumZxPAdHi+QzGJ
fzGbT7j+4RMmgqNNghsiRiHvj7SlvgXmHEHJC7h7Y3tKuOFlxyG0YhSLzy5cN6rvFESt4RsPTC4d
7zafVGJpqpg0B6SYWCdA1p9dIPqp/NMHeSK7g7ncPQY+dr765/g2kIOi0u7BN97QIslZNCAZkHr4
5eGIu9sADmzG2Rd2ZbxQcQ9mtZNbwC2leCULVwA2zmQfaMl9DZvtn7yPrdaLRdNeZdS/byduQ8x7
49YhnrAlyTHtVwPLs5UvNesXcyGuhbxhcDgau5MVFrgPHd8c5CsP/Y9tsBu+ZsdC6Kb1fWe0gUkx
5XOVrIAxeXUuVl2dh+GfCeQvbIak2eUvKRY9fmkdpla4mw97oHC1sE3WWsMHGpm8YC1Be10TG2m0
LipQLQNkB2AmgrY53SgH/naBv9Z8srYc69+wdolyvfKixTa9sVnTWyy3dQ+mtKm+xY9giCrYr9I3
LAdNBi2dkXEFteqdY1ROwaUFHapTJR3VD+2kGH0iT5mhNYGkh3ZfkfBJnxLSK9e9qkwiMjDqO8JN
/6mMIq4XVCoavk/+rqLYpQt5WZuCZfUCmFU4XFhysJmQUl/zZWdpc6WvBHO3ZSMyb/dXRuQY9WS+
hDL6F53MT4ng8qSgC8YVvHdCctqVKDp1wllLIt1Zb15XKQXDL1Rv4VyC7m9rD/AySQPd62jXBeXQ
JBSf6Jp6ngEs0Fzmi8vEVyAWfpwkU2PbEbBmYqn0FdNhmwmugztZwQUbFhjsSUnYzwFM1IxzHW3O
bx7psxZ3fD25+D1QlUqLSZ4lGu7fSTyePjZgk74LW1DbmxpKmhQ+ovdY8anc42RhF1HFt0TquadB
aQhONCmWJbqBTbrjyC31Yd8u7L0XF7n8BbT9uV330Aq7Vph2j4V0Ksroew34uilBSp8/bbvjxjq+
wvTwcXaBrJ6WBi2pJe+5Df1gXXQuFSCpt4pk5xkAps6xiCTXHax3iik1h93UHfMUG1TPq8WLNrz3
d0hRnO7/VabqBmcxrKQ5IDgQiX6sAYqSaqN5xU9R7SuUZuN/fi2/iXI5hY5lgIVLAmt7eOIZbTOQ
fXYPenSTUqreYGgRpuj34FlrJZRwOe6Jg5m26BGbBcl2JFkb3miVIMCYodmvqr+lE245JHrU6nX8
3KvIE0Q8RtaET/tBb7Oqa7mnqijlLNUNo+W/y+ZmzgmhZOZrPDhxbtBU1XjFnbOczBwoS3RoNXr3
xsSt/g/FPyospRbtX+Xt0xchHDyPsXuXF0RzTXZX3wdNE72GM9JBGF2OB3BFwgiRLCpbHNyvdaki
us0sWKvJ69HOQ8/vWFsxWoY1PZyr0lzbvEqesA7cHhFIPmbBfPJpCPmWGP56t4SlJLbMqPsf3E2F
BrIEsFKxL90B/LGvRwOmrxeLlt4v/IvURq8bKPInYPesKBFJkXGl1KMLzqFIyGpoLfSIml6xN9vA
J4xuCz8BJ7dla9e4eXLzyC6nMWuWuJ24CDuOxbbIaOsRRpoyoF1xPq5ygAbRKK5FUmD7TumwSODP
b/hdaOFmHHtJ9XHBU3eocMckhCwhBluQJdyu0pj2uADEM77dFlZTdHYEnQvk8CqpJ/ooFftUvGu9
39M4EUe1AyLtPsKjnX83Ia8ZYfTeFYIpg+H5n35ZGNWFdh26xf/Zi0RO9SMjObgbbU45A4DY5S97
8p6BXDWtn8AwLlQPrBdKUsdV6qTXucIVPk9L51ikDDEUOZdFX9+AYFoKNPKRXrIBoK6XINd2dw0w
VaM5DRn4Fm+ak+0TaYNpIsOk+UbXhLVRI0xu7/qWFiva2KgM8YBrKasSUjCMQvcQdKsBaUwZClxJ
sWAmwOkns75etdJws/oCB9HoktoRrKxlgEMRrj3Tv1Lz9MsA1gSga7Kk1tsY5YTtzKi8qTfumhbe
WAkVcYNJrJlKzKG7TdqqzecgwWtyZsCz86SJvgvzVanC/ObDO57YyBJFKONHlLxXtowW4u+/Jb69
JKsoFPUvcIKhkGWDj/9SH7jKYvtlKUNordkr5rFlSeyO99en+tIKOWBGwV+shMJfO7Yp30Z2Wa+A
such8guaVmhx1XB92J6RMi6/t3M60DHdjflczubwCroY91/bXqiMDgLklOFaOrdU3zcDdO+SPZFs
0168jMCIvgePTTAf835gQ+WR5+SEDPFPX2xY/q/VyhzKfWs0XtBHeIOu65ZboaDhxS0u2nLXT1ek
DIj535hphAyDmvO/t+Feyz0jOEr2e0OJ6XsU0kvcbgHpEnEagKYYt6BSY4OLSeROet2hulD1Y6zA
vwtq/aKT9NoY+aPeQxxlHIgcLKCK6p8UPalyneRhjlJ5fg09OnNPtXT1bZz1V2c3Cc4uogP68/l9
JDD5uM3tovCHa6ANpAqf5pGqiXUEC2BxcAsglQJSe1Y9m1u/ZYotzuu5T8fYewz4Mq0QDqM1fS/5
JrjTA+JYJ5sPW9DtcsJzRQc/YrE4pm6SQ/hGx82OfYA155hAYkpS7xZ2JFtemPXYpdKWPaQEbuKs
cvwtr+Um/uERShFfuslrhwv/LatmdffaqpCKfFZz1hQN84C8IUWG49G1hdFCQ0pZxqaaEROjI6cN
GrCom4rW1U8qCtt4cB2jh7lcOKCcWi5+mJKsSEkgW58dqcr7Nb+xFUU3Z5WWD+DL2PozRJ1+u7hv
0TkQZ4jjb2ia5rthBZtznk/FC6pVvgq7Jk1ErvUoA2NrqWwrM+Qaqf4WlOtdIlanqkoFqeR4TCos
XoeRqItWwMUcfq+fzwXHQjzEanX0mIwpcCf+L54k8c+M0i4mPfsYxdCsL9a0rp1Jh1T1X7+99kbL
KOyl4BlOUaHfexwT1zIm53AZQV7LST7FpiIvkxjK4gv/3EiKOTosYRi3zQitecvXxeVBNZ1jOt2s
PCUMKePdedb+blPRkUm07m3NEKddvG3FcgO7zw0zlleoW29Gleu6LRQhAbE6t7MqrLcx18NhyjEg
iLf/Q5En49kkXL47zBB25AWPfVXLlNKyxXMWiHYhTYdcQkWUtUgcW8wGdit0n2TVqeiPJKV32vTp
geC/kJybytJtPII3JRrVPh+GZe0vFQaIaQZv/VXeu35tCgyHcpG9iiFwMH/HoSq+cZ8n3MIyi4tq
61Tb4hQnHnyfhSyveO1WO0jeIu+CaCrf5s/nFeXH0Ozb0ddpE2+N9J7wJ90HkBz1dMoqXfX/L084
d0/YRxHVErKEG9J6r9AIgkSP2cJXBkd/OlfW5/7P616mkwtjjsL2coOWCJUfZWkoyKicDeyxm/qA
t/KWK9fjSRHbhkh9bZQjInfa2Quc8m6mwst6ig9fQ1uwvAkpM8HtE0YaJPhFvKkxFpW8Zo3w8YLH
PiZ+/EBQO6I0ERcfmJ4jpE4ym4wHNyTK4Kfy2jRhwD0IA6mXpl9g0W+kb+tjfVwZFB5DSTl6mN9D
4ELV8cOmQAM0HnmDmVRuphbqeSCp5KkdbQf5zvSjoO05hOqemdS0fT4Px5h2wBhbFOuYe6RL5LS9
AyCBRwYNAG0AtSSkLM34bPZvLaA3Rt/a3Tfu3cbSuQKXlmdvTrK5csW5rMycMflzWFS0ypBrYA4v
pcxh9hyvPwNSBfHA28qTzB3CcEMtWj5DCPl2ilgC1bJkj9G1c3kegxOdIZq7+mSzPi6ZQv1Gs88C
60QiCK8tIflvlVvW2WOp3n4McPFXB2/YTztDmwp5kmX8rr3n+YJV/S7ggbgKVmIfzkxWQ7YW1vNC
MB1ROFvMi+waYUM1hIVdhBvGUGgqs1aC6ZdvvkN7kPQw03Bip9LEmSvdsoNdR+hi4QhbLtQgY9Ck
OyHBohfTxdChVLQRVwLO08CcWa4372+053x91QNDz0APvX8x1PhYm0ZfnSQ1snlZNWbnvSxNrC6L
sbmrS3hO6BqpT/4ltVywwDrzyxGEZO0oCDuAXBps4aAanary26fU4MPSErObtNZ1wqiMmKTI5i5y
tQ0dZoya+UHDVhq2qzAqx+zXjxSTE1eTjc35uLvj6tkvamV1kLz3vBBXlw2uclz5vvTLQPbuCrBV
Z2/B6zwwU7crTdy0S58+Udfuf21vDLElz2Djjq0Z1vzj3Z7Zn6hiZ9h2c83qyNpaVVJ/ATs+BCSP
SNkGK2J7PeCdX/8C+H5VAUwgEB0jZPAu8WufeP3WGziP9P1+yOzucY6P2iytdN0eCxN/k0hYCwlv
5IWWZKXu6EHXjx0Eenk7SA/+VJNCymOmdt+WxyyNtRSlOpC2KJTePV84PGWetv4XJLduqkFp+rbB
JkQUZrXBPXlKazGZmCi5BPWek1QuDQQ74loXPXVyqoANQbDkew5qiZvMO4as6E3UCFFDYDpXAFMp
edVJ4P31BSMpbpGgcmCa2hk33RWOf5rTU8z+FP9RcJfhqfOKZLKw2OVP7UGzeYRUo3F/+RrVa+Sa
sDDHH11q6POfOipQsiuorkzbPDfLO1M3emAE8RzXHBTgF8HFBUuW5rz3GgJhVZWnxAYq+/3qtzNt
nfcSO9aZsHMRxjFjHaJTvof+UUIeYvs7sQ3E4PL8cp6+4GJ4F13kukfMfBdpjyAEZOuN/72lCFYT
oxg5AIptf0XkUPcE2bJ8vI7BFFBzwYeuCO3p7tFU7P3GN0hDdFZ2Pedtm2Ukae3zLtmlMd/l20t9
3MGWMp7TpXUFsQO2aW4X0ZPQxDZUJzpoDPjBL9x6Dm5T2l0cp9G00YlLX3fxv+zCRKltCDKHl62B
9Dns/T7jPs2CgQY741m0IwxsLcR9Lbq88wyvhiAdpIXdFnGbCtmEMDviOOMffV7D5DSoBVDWBE6F
Qyd254XRgi9Hn9BB+RfCEb/AeAhyVHr3yyQNdyaESdDombp+wZu28IFsMtU7/akmO5j23+gwUuSL
UJNG6/FLOgxpHZjXl3yonLuzORLxk/AiC71hOhInreAtQ3MzeAapyJfvAxzfQ/MDq3zN0DoyxgKT
BFRbTZ+TRoT/TvBJ5ql4CxCzV7UEP3Q/VMXXJTOTdulqVB9hvoVxzW2ebZ5QQBRRTuRuceARAz4u
F4wxFcBQfOOv0hmLgI6sQH3dJKR80ErRZQTcQucQC+OPNRAYUZRHhlqL5HVGX6uNjCpNAhjizuvM
AlT861s6CZDIfqURmm02uDkODssLkTlAQ2IsZn91ND2wSfHb10ZVrc4tqJLIztogjLF7LoCu4g7k
sEwwVo2SSvR67/fv/lvN8oE/L6b9Pvs3LqL1H9+lyTDcE41ymSgl6xdH323LRAj/h4rlpr7X8twV
2B8DZ0Z6hzRcER+UBBDYy0/pZqmcZd7s95z+THlJXxLEYJgNJNi/LNFz1CYPgKxJf6YakZTx420+
94NlZ6BelyxCo64R1Sa9iTXvyNMyqORZV5MiMAVvjfvS5eZ9VGX/8tk6bim3cjRiVI8VSOFfATX1
nhs4O8Uu9VsF53FTrm93p+iRlkJD3FyukaqULOfNQG1BUr+YgqQm8nou6SE7VRqIzwX0WfMa3tmM
TPvqpwvRlDBryGSroTGjn5rkisCoQ+DVHEPqxUj7HaxdQ/nqGeU+O/IFtP+DAYQIXXN8ZKJe3jFy
wz/RPGOVCe6GvTS2fsEY657vhQnPevbKdts8mDYKE4EAZjPBV+Qr72e6o5G8cAvUMWZKqdUib/Rq
O/A55gPrHI22wWiqdNKQ70MNK5YWlzX0Xrfh5J9pe6fLVcYggBGG7NyyLSicNaMl4qEcQFTfMl/Q
8Fz2P7Zzyrg44HUp0G4L/evssP8haITKz12yZh3iTskLfKg/mDpsDqUbWFQ4utcAZeA0oyq+9YRM
7yaaNQcO+wWIoODo2g4rdjWgfYSGLdPpSqgcbG1OpHgXFDTa0yBCmeatVK5On8rb8mE507r80nS1
mBtYsqbbifW7UgjO8XCOLugaXx9/KQNKZlbLjOxfNM7GFSfNI1owHtwJPQh/qcHKfGN77mOzVcYT
tGpmJv29qcx5peutwjd9gcdAvhST7KXmjgJYEJ+Hc/VscyYk+AzemlBuLDHQ/yHbms1Dg7IVaK+Y
oE5htbwUWNaDX+oPJh3oBjf+Y9/AbXvebHPUZReQSt5pNq95gag4G9/zCq+EGy5Gly4/APwTPznW
+c/S/DhAm0/c8rKa9F9vc4F8TSK2xkA/UimbDCJocZxSzG6XkT2OdP/gB6yOCqWbMqXyBpOTqX0I
VgazDs4SDPwV4JR5quhf1CmpXGOWsH/8FekT2ubMVydtYQWnuS19LswlCnxgXzUHI3Gdv8hBjGSZ
KjDBQmqqXQZnZp/b6fdCpKG3VIgyU9I6Y0Br3ATeVqm6xMOtmS00Q5Lqf0jj2E3YiLsDETHPgbTw
425BiCUDA2+8GTllSW9C/rVVH3R1nYFRN9aqP+u2C8KrUUOnUHUMNGrrXkkXAZI7NvLE74auXnMB
bqZMDNBR3eN60ZVpOAumoEJwSy9uI4QnCIKwFLzPzMcV3he6MjDr2xdatXYFK7/ROFdBTXzuLaRc
6TgX3qmmG5qgsrkLyDCxh/HyxsCUhnlnLSrJ2zPKwIRR2ffB8AaPXP2njNUpOS6bRk6KbyuuI7Lb
8C+ND8lPO6bgxayL6j+bcQxWKvKE085EIRofbLu7nGBAMhEjyKX/QOsTmQA1NhtoTS8Wk3sszJQ3
WgTyggG9kqjKQ5OX2/UEDnxLzFRnWm2TssnJYDD5Nv5o42XIp5Q7NbFB3MkuvLSJrw0UTjJyghna
M2C5SpZrd+t38NnwFHkwyI+Ha7kHg8H29bw7lmBT8AWEKKd6xgrXM2Vdn6eRqjEP0ArtV/6AsOLm
Vrcc7RWzZqaGIHnBmHc4rsGwP0C/7sNcaPeUP7ctFNsE3Dymsb7d7VOHnurc0SG56CESFBKuysok
aBcICtzmbRYNYsmq/8ZN9F+9qfk7EDJU/BgNx+PFDnmQgrxEOQlfe1w83Q7gZvI1D7RO7UD719qJ
pZI/OBdWqjNGNnfkj8YImT2gErWff+e9MKe9+UveRwl4M2mgvCqnv7g1CnNe8V9XzuFzZlJMYXuX
TdqWYHdU6Ikue2IP1HQGbJJOHC4hoi0HzKQzjfflgFCQhFbEfgQzflQ7RRDyhSkEMOTkw7vB1aAo
M+szOaHx/2ts17iddWIKk70tuXzz8tpCYOO+l6JEcvteAyc0sKXHpGlm15zKG/bfggKx/ZhXIgyQ
u7wZpzsbemarMHGUTyG44X1nnKQ6y0yDYQQpcFxrzTeI9uvVy7fbjSsE0D9sOEbKdeNgZ0oCmozB
0eVotAFSapaHLVxerQfYYu1ZOcO7XIlIXDyp12+94A7fx/cYhPYjjKhCkeTBvdXGlZvWTfR1xVd+
EKpN4RzI+QuYMH0Pjtyc9vJK7a9rSL8YcMShfYtiD6i5gSFXSaViRKYF3uAXNCMyf4Wn2TrF/iK0
5uUsnB2/bkl623Wr7puRVRgNMytqpZwydwuNueWGZ0h9SzBVL19lxnqbG8U8N7u/hk7MSq/RCXHZ
WvXQUqhhUaVjTRQYfRG9k0d7+Q6i6cIMYFl27k0nGc8EoZ3UoBMurhH3bZCfYEw3KvyxLXuuFuGZ
Drt/fwGYuMQeBCzSnLtyGZJPBvjMK2xPoFlGij9pUwLBvZyvUVTB1bNMUMUuCTqdewc/qTTMnMnu
0bJfpBEB3u0GE0ozaDsE9G8P1QGvyJhbSGxk2AtCzB8yIjDXhNN9Sfp2fJMF2izUI7XCMm1YFkbw
whLNk5vOpW57kKuknaw3KDMvN+xQH9IlKlh5KGkL8fAioc8WNzTQlIcdb/KW30wlqUpVk5b92rKq
JjNjqoW2/ABeWzcPItADsoC9Q47fjLMN2tE/EhUg4pAvG39Jl9bN1sL6aR3rscdeQ5of8eR3hif2
7Td9sRxIcJF9md/5LMC8qhdE4ERZygViNvSXNpwknLuLy98y8PNuemxZzOa0TBYZ8ERBC/KgrX1G
SD3N+xbxGpnBa2zIh0E8124rI6NrVu3g0cIsSWMtXGZKwOpl5oiDHy1vkVcXM7FAtlL4yHu4lDz+
3WuwKnVr2J25j/8rDDUL4cAAyMl3rV1+nfc5gEzi1NFRAXpFgLXG36R3fTQAJl3Vj0ca7Qd5tAIa
AV2Zq1bK7km/OBKutYcg9zQ3qf0CCXd17HfrEdTzblijjNAuPO/+quBnaXtgCz8bwfSRwsLJcslZ
wImPnkQ/ZZUB5eEEsJQhXXlcT7p6oNeRFJMgFbSVE0rpdSabYecmjjGgbhz6kUjY1v+Onw0ANBpQ
Hz5jHLJpjSZj6p3j3OciGkctP5fvXzzTNKv169VlBWLsYhihL1LYk0Th840ouDM3El5/esNnUy6h
ej4apMZCxgUVv6BiU9fmn4TbvEKIDhBqT+WjGcEC9caTXDFZ0nKM/GAN8HWrt0eCK0Lf74zG/iRz
0BaJBRGjX7y+zwlHz/XG2YkcnS/ZItIVlxuyJqvbP3JaRLMVBVZwx1aw3nPKLgz8oIALxTFP0TRa
2NjLSkDcn3FPKhYsnyGEQy7ybuuodpoGAtx3l8/Ph9lmAh1sY7SkI+oGt+9C0PlPfQpeT5maTjhw
DRdnn1yWtCj1xYhAkYIMYRqfM0KbZzvtsVqC5tMmJbA0SFd83wGBaVDGVsK9GghuVCLBY/CFnIgf
nd/1ARk7cF6nc0HGlAvxUuz22S+QFz4ERmSJ5pP369hlBfiYu+L9wZ8e23DtHnzk7wtUFiOGToch
ByzzCTFNvyKE7/DZEFYF/SWysHxxpjSfG9BHOE+fh0X3Q3KQy7Mw6dHLxg0poCa/n50FUWZY3DvH
GcWEKCMwK6G/C2ahruu53KXiHwLZxKP1e9QVlS0pIxOUF4cfKFisNM90nohB+AwXaRuAoErDXHC8
ya583ESbcT7WllA8brxOwy7gzhFhTZPmATkKNR7KHmir6oluhWuYb7QD1AmYMH9ZHMwklekKxMDw
ekavetkteH5QKszeS5IiuJFfAGNwMb6b/N5GEWr41NFv3n4n1T227LnPp2Z6ORwghSsMokN7GMeQ
rpOrxOfc2grtkNSErPGY5408077kmr8Jf/Ng1g2V9/T5KYNLLEMewazUQjSUb65sCvklJ8xOUlnJ
oE9oUcEfo7iSTH2EoJRfGQAUrhe2UXXef3LuDX0XH/ySQKlX+pGNZZazWd9r+EP4IV2OmkPuETHf
xmCGcZaNb1LFlWNRsvBYbh4qwaT+JISarHciNQoiTOtjeizbr0wvwkfkolDxvhXb2GElw/ymq+eH
RgDKzvtYpzkEM5G6L+uVJYMRVuqQvqpNPyhVNbT/QqcQtlbPvZwyu8s31vOkApDyno9engmighEP
XtA2nh12ZmVlpRGf2bUYxMx1ePJnBHBtu56VGBlfzJRrZL5MmMAKhIW+LDqK1qw1E1GeQyFEjSLn
p37ZBEY51dS5PrB9zhL3VmnmAWxeDaX1UnBiOu2hBkObpgsnaOm9b5+RanC+7I5LmsBt4+SIFIpE
SuGIXH9OcS2mUiA+voeQCaMRYiLB0pwaTup9TTg/UEX3Q375p0Z8PowZo9Kfgj4YbnhDu9guL+tl
MURq+hRx4eBtkB4abLi3Jujgekv6cWf3Ch+HeXBAj65hHEjTsAKRS7U+gthriHoo9m6vZCvaFd5l
1qLe2JtFfEiekSwAu8Yw2hnz/cQ0Z9uM4BWxgov7VtHR+da/I8+54DTdTxNT6JrmBSFioVEi3cBA
IBr1Y144DovPacUedG9RPQ4txZGDDaJ3MTQzk2FFvnfdxLgyNPefg5Wh91xKakZ8+JCZFpXbCDU1
Q7zp3790hDkcmERGOQy9bitdYhu5bl14UOL8r81zze6or07eOIxKErhpVM9TExvUarXExzpFB+24
NckNXunM8zKgWRcfu2tNJCQO1iTsYQHwSyBZfpYSNrxkrNiJGy+YYLql6XX5L54GKqakaWqTpKyz
nWvOadlHGkSeqDi9mRLJc6ZYPxmG5accfMfkg367MrJA3J6HafuH2Ezy0oCwQ2dRjGT4dG7vq+d4
+yC0xPJvmHd1SqPNelfJwsejf1oPfJ9XbaOYu4ITpwdEyV57LwWt5Af1Nzo0hUJxNEfCRPkokJNm
9su9I3bjqP9hJ9pyS/c44d6mS+jVFojhi+Xi0kPUzSVpPYCWf0FbmKIFUn/IKFR8k46GxScKjZ8A
zQNCYIk4GfwdSnxm1LaU+T2YHD2hLn3p/I41fdZNC+SyQ0uXGxhtFkW5/CtuyJmo2picyhyosrja
ALU0IviHUCNppFJhqWSHqhPzPbDL0rbABHIfOMcoJwI+qmAF2zs16XATls4ZJIwAy3urf2zj6ZHl
+Dja6t1RGJ1VrLS4f4SAMp9nujCn/TXJIlQT9QnMSVf4nLuY4RNseJ0nsj3KfQ9c2JODCa8WiJyf
1j1AitZcBvBkBoDaptG+XL7GvszOLmfbwyvI5axZDPUYHefoP1XvvitW/wXrGL2EhTRe4jwbcN1U
6kkMZqGB6jelywZV5xyBoEEWvEDoGJPZYYtXY+iHzZV87VhRD/4SjUEiw44Hl1indKVNNKBWTnLJ
i2kEuihgoDngtRq/g48AuIXL9ob8UiPKet5BaVYLzL5tHKJIGK3fm3zp/coPSIJddEt5+OKKYRx5
osl3qCTLwXNB/JP8FP603YnHx2OczLo3YWvPPst+ohP9xev3HuC098wQzUPVaqWFo3dBOHfxMfCb
BCfDVw3ujEDEUBe8XgNw6s6QOo3U3VsvjBB7Gyg4uxvL3zO2z+LoOCu389I+k+6t0iwvMIyfjXkv
3r71f7HObIQU1J7vgHXJBiD9a9DPtZX4NnLeqZLVkCOzPbExQXmzMyMWK33GmpvNMwaVrUn5J96N
JY+Myaitj2vFo3PT2aDJgRIv/DdX3aVXQTxGH40Ej2/j0i1tH8cH8W/LSiW6zAz8Xu23gacXkBRO
yz2Vw3IsqICX2RPJhntsJlvSybxL2v/owR27Uvp/AJvxT0wj9YP8afsSmmXOWXVoCzz2oIHvYWJ5
jFu2ssmESZikf+19dhgDGccdksT26M+CUl9M8AFt4Zso6/epo9UeYVQF5L6oIKoVdCWrAyhOjt61
tM9BDKIy/+lD/L/AGMLW/btMNAKSP4FguvqCxU+QDJJJTt91vx8sG3bRfZECa8rwhzH2pFyUSnN1
yD/Z/ZBtTmAI7Lt39CipbOggmSVbORrRTVpuSqGCIISOL5lQ6M42guuHpxgnWMkE2EIdrKIp9a/b
ZJoHwqSr0KyAK3ofRivH5/USZC5u73VU8QJIwuMM5BznuZeAlWnNehC/62OA4loPr0sEp6QeequE
tJgFYIfGoFHbbFzJ1CEC9xZKhxxe9YdrBRv+1j9xLkcDgPMHlYAv3+/SL/KQBYFsxxMBkQ2401sl
5y47AdIDSKLEb93PAoDO3kn+JR7FYqXgk2SEFAGMziIcQ0OnOWe22Rxc8xLgwcsJx2ZXGI4v+1ME
aZ/tHEJ9WcQ+VYFg76PAWw2lj5vI+6a+4z4O4O/xZVseZqZ70S9fca4krU7XDWcEDwMnpr9I+wdS
VCb8tXLCjwU+8T8kP69ppy2zCZIlmfWpojxZJjojFR+MT/SqtikIek5Yr6Kah3HFgcMR0TUQggOw
uU+SP0ge15P2bgqesm1GGGZjQ3ALBWGzbA1NHw7MSyHdspxLE4F69EL4OEC/eCc0ezsiJ4Bbx4Hc
4uZKUoxxsQpMsppTHqZS+wJeS3kVmn/BrGATh3KqyA2VgB+j+AVRFSOVdkOXNlmnFjIb+iL2cuQl
WBNdc1xThNGJgnWvpKdSdKd/53lrZNaf/ors1BdvE1mnzLTESWB0SbMUmQqG6v003sqsFmAhy5fM
ISJau2wbuf6r2388FwMs/Rs9BjyMXG6nszGjlyW7+PFfAedi4smy1mTcoyY3JDF7IsKz4kjoHZx/
o53WMxAX5tYERyDhb3lQ9Ibe/M6zMZzvad5YCv6lc6G0jkMEdqfJNVwZNYnNxyWdEQxt3UWXZ1hZ
1VaX/tZEN96J5JWzk1VAuLH/uWq1v2ahyxIFatxooTiRPxg1U5cP+DuppoKAwWiHjaN5DVgPvQNK
js5wkAuFJubEINuPazO86aDAdJK0seetS79ybayu2twzcglMCW8bA2Jd9MNiLMUVshKkFAauaPr3
hDJoo2xKuQXRD5AEQZ6tkwWij8AHhvYmDyuJlJt3wn4VeYJy2NazXsKJ6d3rGb5knA3FqhIm6m9Y
GONRJryq2R9UsyZb11PDNuPj60Cmmg5fSajUCf8r0+nXGNmCDlS9H1Kxc7K0lbR6TW7PuA9riwg7
bxMT2d6Lg7xYwMRbJI3s8S7dC28UfkiGnQN6t0bemY6hqoqsw0SpLS/6SMXGjzOI7R1xRxeu3iVe
yZ5JhlcxOVpcRlDFe79b/11WBlvhbbLVHwBinQnsHmLt0+wkB7RtWvPsNyrv7mx5R2jpdPilpxc5
e5IjkxjSX2MmPE7Q+2Y9LfaG6DP7UdY0w+48fK1MKmiWbTfethNSl6PooNgPxk0Yq4/74I1G5e3G
Mn6lVbBARFvYVSQywD2WBz67j2koSkYOTfhLo7zy6pzggGWP9TheyMAAWIJmFyBmqbomomDUytru
XvfT1wfK5aUAXEqRUN9sRKMzwdBKzkRdR3NkirceRlF9UnjTeTqDwGot4pnnDZVElkW/McGNzEr8
E0c6o231WxPiIYPuZK9Ky2/r5I8PUu36jwQHOeJeOogVGODu11EhzjJNOMIZPZT+gIMnedQG67ru
w8enEw5TGF00zAG94+i/oT9g4IfK74NXEcTJmOBti0mJebUcC6PUX7C8vGG2MKM2MDAwnZl+b8NU
EgCdai8RLxX8lQ4eDZxrRmY9fswYGyvTOlJNbuxJ0Jpivdr1ZJXSbyVAx8mSf5FtAQxut3qVl1ko
CZ5345ThXskgHur2sxepy7Fftvi1v5cjCfUSQjBm181yn9aiwYaSBHJpxColzWj4y6v/mpeEcQ66
FurzJFuOXMbRMrowgsIKf4UsWa3EtYxq5PpZuiIM+z4mHoUAJvN75+v5LpWfFauY+WszDVlV6Y9N
4gHjJM/wzf3VrYPPJ/YIg/rah2IlKHXmXVLRcpmvzbB5YmWdr3YKdNaCoquVNhaTqUueLx+Xz7Oq
BHggoat2RuGBm5pVYedywbjgFN7S7vNMa+hz0ljt6L+plG7Cij1+5QzpwL3RXc1r86BlxUyCKrP3
KYHSwOYzWvxl5kkQedO1An7iXC8rQYXVR5GCAGceFPVcwYKzoeooqepb0Rx9AF6/6OIJPwZkQ/Fo
xqK7oLwnAjPDcmmq3tX0q2IDB2jL0UGpFGv8nLgFLwDN3kiqQ87cIMe4+CGc65HcPDPLKJUuskCc
t2qjKGXUDvHNksWg5w6HbtXQzbjYP+cGRg51R8LGb+DmJM9dREmFreWCcpOwhGvQxzcdKCa3xvVm
+IILVp+VG2GlRO5D4Z8k9EjQeggABEKRP9LktdNvrgB5LwRnzBK9gv+IO38cOoJCn1tIJd4R0sM6
yd4f/uXxPakDXkWcH2diHOMuAEFDHsbnEVLO2lOIMEOLwVrZvZ/w97nD0l4qot56XUHaNgi+s0Ev
PP1DAEdtizTLgiKIjWoNTRe7+JXzFsTh4A9h474ucgAHWkNUdigHn6CueUHvUF1WeaCZaihOWUxL
fiGVJkNH35buErw+zKaPj7EBoePr94WCYiwC2VzoFK3EsSoHxq/UX1IeIlIgOI0IvjHw0yJ9UBUX
8PiTXXqxoKNbt9nfvFZnb7cRRX+gF7zn7d1BzxMeRerFS91IVQcfTNeAnRqID/PPA+51W4ah1XAv
Ywjo445qbU6Vx1wAMuqDUUbGl/t8Jqsx4SzC6QWj0Y7ZJ5NCFuwW/wLfylzp3cItqdA3Tgha0DeH
UjOdafyi3KEJ9YDbGbQEY924L178yxlERJsJjIl0a5KvRzZ5uvUaDA3eyGsznYLyvFZfXYrR7/Sj
wwUdCMY0ufiGh/Gz9OFY4QuNHnc6Z0Ls4H6SWKnvHcw7/z/Okh/sFa8R2udkBcACpPj59kPmPlMe
mr2rQJQYqh9XvLppOjQ0ArHL6oLVPCqjBqRQDj13ZzsabfsR1RWwAeEbjNUB5es6KrfX5ImM7CDr
C32XLg8okjI3xe5FlmOdGgzuWOWrcTy2YeaQt2BBjD2tab8v2Lnx+EwausEnIFJ/x1mv3oDposoB
eUzm1matwqYT87w6EOrpVUo+/AN6T2WNUP+ZmkZdLbK4NM9joWDmGvLjYB05SmXpg7jl4b3tl1wb
7Hh0HiDVgqMYztsKKfLYkNlR45ey4oONgcz4errsbiM6LlepJ/R4S4eLdednzfKyIhjeI6fdu/Ea
dawCCkd9kDHMYWEOnWfeiUl1yXF6u9tXJsxrfgVycZY0b4FK6ls/J+vLAM1PFhj1YJ5uYNfgvEVt
RWbLCPrxkC4cncic56EJ5xHGzuyiUO2K3TRRClESExqj6H1KUiR2sJQ1uwhVsr9uuDNwgqIxI4x6
ZJOINpwoFtp0LLr0vIcc21yMn0oAoFFFlS1KwKsuYtsYjmie2VwhRgXYMvSRcsTbh5u/CrDoZzER
AH70cwf3QIjFOePOEjVVhqqfFJjrYVolurZjQHTewxAfVhLHiSUVFjimdrh6BkwfGFyxcNGbXbdr
aM4/FaXHevAQSM/9ZdE+CELLSrZVMzPNdbCh56ty1OhG0LMs6RAdAOdxxI9O4p7S7K9qKD+DG8dQ
lwZa9wQlS4XiOZu0TIeGaJOa51GoceeCwnO7vMJL6S2OoyfygQyWZVAyTptoFy8gTfw6pMcVsE1L
GRVoVJxEteBwLIPWIly9Rew8JOGBMAzEsBNSVe4pmg8LZTkd9S0QMmtEZOKfYRsf3o7Plf+wpBP7
H7oVlFXF1+jNQ36R6rQYIzEQIb0AKYD9xDlW5acdf+tcUVOIKPJgfht7AxuJftNpXtRv1kR5w+Oc
VJaOoPX3x+vHShkUj7Aex10WWqD+Yk1juuCv5e5yfA7skBwX0rG9DFRIH6ADjE9EiHIQa+yTkD+4
kXAY2qA0KtjWzLZPp8uk0iwjqrxt4Y5XfIaONhoiJV7RJLCFAjnEFMLszQDa1ynvSjlm9SzMd1s2
Rkg7bLyVgz7/20w0Yj8m3dNIDT9brmAdzdAy4EyYRyRf+aQl8LLg/+d6z+Eutrbud7FA/7MgXW9Z
s6paDdv6+bZJKoksLdu1d1P/LxkfZ6/9rcUbsTTus1HU7nMaiD1psjtpIlGKabYv34KUMuCPWB/a
IJRwzM/9tIPXUsOATIOgQ3Kczzg3pz2QXGAR5QDG5Wr5JNWnJ6LQIxXS8hjQYsKpq+TtEnx+sa2s
Tb1xSM+sceZ6AbG8omBi56yLgZ/YxJuVdbmz7YCdhx1khyemhFwmniO4Z6oAgzBGteMfuHzY2I+C
KPnQBFUiTTKqRJeN+NM4UqLereHVEjGtFFJx6IvPOZOQiCFSgeU85W/0Jmp7iLMUa0EWjSwNUFZ/
2iZzrUpCbqAQ3e2v+rWtG2TqIJEko7gDAU39ywjq39ukvp/wTk48iRl8pIv0JrBvkz1zobEZ+LAk
b0yY0agNeQkYNrStqyt57kwF//+lqB7m6sTEw1EV+Y2LsokiB77qzDjfEReiEt0z25EOZeMZ7QY6
6KH/P00lyyCibEexxLeY9gDc7IWKtAZVs6n95PcEpST51ur0K69igAfxnnYLXyc4HK8+hCVSt8Y2
bdku8U7rZeMcdQphHIbeCRh6V8P5JIYMPkFu4NhWd8EkG8A9VoSpc7zvjTwpeqK6SrSQuI79gHdD
LHnQ7Z/p/APSeZ2McMiz8vjr09s/l5b6K9bq/rkIlo+AoVHP4nlH6lFQNjWvIyJCqutqVG5oh1JR
eZZH5z06L9DtBgadZ7/vlg5XB2eRiAC1kyPiZI0kHUpgnO26hMSaTGeW32raBqdRAZWYzgjWzHwh
Rkt4oOFIjmIn3/B63DgKsZwXDNAfobRwEL449FHiAKUGPWKu5/vEQ9+QnUactyGsP1bodOtZjwVi
6lx9AS07Kexnr6t8SrLa4waUOZt6pZ+8OOPMaNuTxj5dYxkHidRClMpgqSK3gSdaAU0GFbW6ofaC
9/BVPQrrsSLabG37XfVlSSCb53zPML5H3qcN06VUo1QleiSdz6hO0M7V83LnQ9gBV6C9QGfMohRw
cLQR8bdCpNIYN304mFd+ig/qVxK5UmJGqZ6oXxUNhhDlzE+zgmn9G6MTN27bFIRcp60ZSeHvGVTb
I1A1/pnS8e03hpietWJ7bg4Sm11aCtB08XtzJOuJjqqgOzTwFKH0eRxP0f+/fj108xBhbrLqjx9M
wbavOJbkLn/aBOcv7GzHRDc9f5GOwudlQ9wuC3WGBo+svFMIxJ+eNlXv4+TLdLD0QsYctn1t301W
Kso7aRaUNSkwXmpo5BEyJjXBZvas8t5PXs/AM7uVNDaXYJiUwME3oemdzivu8rKnak0lP0zu3L5F
1lKHonKJMphXdfyBxQ1/1QFu/TR9yk6EhcQmWj68kXEAMzPc0Cg/u+xDOEb7HgDKoTQ1WAIymZnC
Ms8Q805HiNmKM4LiQUyOPeuQpYXA8yY6+kQuO5/6dAYcTHz/n4zR/6wVgBu1tpHAg2+cmfJvQNP/
TgZIkzFe9lFILl/MqW9ETJmPOnkAxpsirBfEs4ByGaO8ODmgmUzLPMaXPrz17Ux9Hpv82gTLpDUy
JkFHh6cabwPS4qST0ILzKJdE52EA2B5ew3c4lsyKT5TesRk0SXYHsvgHhCD4ZhHdilRStKAXmlhK
v/3Bx8inE5yPs9OB95aY/Ug+S307/LGllxHATjrqrShKbED/yrAnO0w+tFEd3ZpRgdZf/uh3guD2
JT6tabk0h+PW/kNMvy69iu/RHGU3laZIYpiLX3dde4fr4H1Wmficavnf6fij295mrbJz3eDm9yOU
0jfpHpMD67aCef07+yRIiL1aQFbAsxrJSyApVzns7I4hmTVHuV4QCcU1WtEhvqu4NpNTEVMGxLMr
2nXXsvMFG+16Xt7t82XgKI0yFqUTbh+SFUfx0LYqHDc/4hqs63YahedXbLPlameqpeWGQu0osB4v
9tv1o9Nbtz7VGedsHxmZJhpL8ZVBA/HpLBEbbgWXBgdMKcIe+83lEfhVFApWoT3Ip1Avo4f5whe8
zHWzm0FzBvtoS2mHbL9DCxcj85PZpywtCa+/tX5haUf2/9yGbqxb1rBN5t7x18mHvsYN5H+lQkXP
pygU4/BR9C4InXwuGFjm2iDEbrEp/tfePfQ8kTD9dii4TCaWSDm1MJBNXbeXKA5Bh6HCfOISg7NI
tdLCFQ1zCLyELUtJ2VyN7kzEdwqZIEytcq+GXEczEAJYjMm4073Toh4/CfvpV4Yo0miLAs2zCQ0A
/89ESMBOjtV009YebO70/pT9s9mVLXqfZfE/bXmPI+B47PcoEM5k8s1SGAylZ0uqCEgWgsgZF+h6
ZLCziH4LMH/kTQMB8ZfxGfwmtw2mRVx2VohwW/LoRx7eBbTiyGOjkmgSQCyhhJUOMVmsEPP36ENH
74F+5pGSd9xFn6uuY855Ww+4DzV+PkJBLoMi7aXEU9lzdS3rjWR2/PA0//6AUFU40jxLB/RQxLuu
DyL+7HxLv3xjLqg1We/99QmUv/cpcgMYbxdMcKTKk8Kotklb51Hv3QvM0mjpOkN3Ku8Ri439IkG3
9eiYcg08Tsi4rEKstepvko8CY0TQa2EKphCQ4O6p4Amwb5/jAjfv7/+pBXiTLG1uLf6CNgSAg/CJ
Jv0Kz/IFIsmh4e76GSK+BdPeUXgy802AOii2D7CokdwNIaA52yoBjHWBPQ+Y32qjRaiqVMwnKUlW
BV4kBTllbFy3B+2mZYJPJEFIZ7CdWHcu0fphgwVTW8rnZdpEURswbk/o1XE79/I6h4+C4cn9c/w5
RchGuwNxyec79PGBwM8MdMHnhkrIqDCoB5eE8wql77cdXiw2pi8zuEbWEBpBvInKI8mXZfHpXwsA
PTqnsTySPuhd+2qDiefK7LPtQJUAJhnMecrO3znEacnmEeHUO+GU0Fy64y9z9VAI+wz9W8JY9zsw
Nmh4ClkGhdTZwOkpgA3z7hJajdrjopP/22Jc1m1v0zQ2LU+NIv5BIfXvv4TGjOSz/bc8HU8Zp3qD
ZzxAv1y6j3atm8SRCchgTwGEl8fZhoZ4hQcwu9LEU8hoOdoYTLauOcxXOVlBIy1+q0E52IeZZZQx
6nv63k6Ns3p1aDq/CRLIv+E4GTqjmLLdcchRMhbboaeCGjttyM7phWEQRhmhhFRI0On3eQcDOXdv
h/gBEnVaSDIm5JPBcWJlY0IHN+tQCikbbljySmAO6xXHIiuoQSl5NeW+6TFNuO4yMM8GhnzB/dQj
kzVkU2L5yAJIFEGv0j3S/M1E7EuOD8OC18PXLmAvSsIy7EYjseXXUbS2BZJxTkY4rWffYyE5adaQ
IVwGrRmyJViYwwrHLR88/QnPhfz8Wnd+/AoAtnKnQmkvVCJ8EdfEVCkDE0zFgzxlNRysNiBepgOM
urOCwChVgBH0JXtYvSDjB9omTntXyQLity+SAwfbM1WpXeqcG2q5XSd0f/mjAqphX/AcahksQLGh
cb+z3JwCIhhdRbP2wFlYQAb+fqpnH/2LVBdSNf8mt+Zjk7+d7qwXcCz1PThDiMhPZH2wmoIrSf7Q
cWK6qeVkKZuXWmwqyC0Y7PMdABx86Niuv/m4LslnTHYr+YciUHmS6VchkHg6Q0AdR13cAlbnwUcs
K4bhVPchGUnuEb0f1mAVVrIwAFYp5O7zdfyhfsZIKVRusTyJD7ja7Tr2h2PPE40SvhHcO6DOYq1k
4q9VpT0HBxOT4g44GkpOpcmbnCT91cIoihdBWnUqDgBQdEr71kaAYrQ7VJRe/1ogWGOx+CpDO0X3
N2SiwDshC5l10m5rAKPfkldrzJv3OmYB8Y+v9mQoepUJLY+/Lr6S5rJ4sG4L+hXPbX8HHijExXGR
1xBUrySvAv8bV5CwzU/gfs2KzZjrfER2bmWyRRHrm2MJbTKHjg7tvIrI5CKLPQIBxEvfLrJZZmMN
1i5t7Dt6eSOV/QDDv0SnsolyoUXDVXfBJItpYZ4zeEYoos8l2/Fjskebfw55633oXaz7VhSQBwSd
AawC0gwxCpJUVl8D+u37yCaleu/L/ZSm8IuC8gtUekf6NizHPVoZn5dz/iZTenSmoswGQCtwQapU
aoh3EjFX6y1L4PDPMJ6mOWVcCwi5/2bPOKlNT2Kpk2yQoXnpLpMbvx5y+Vwa4mrf3GqaT+0KYG8l
+GDh/PMt8Rc4h0t5EFw5IiXwhSHblMw7RRn7tQIZKOUk2/ywUNslm3tnBsTZxaLd6G5Bfx3utBWg
F1tnr0QbBsP0CmLP5eXLOYfHqSzSOKWaP8LXxkk5klhanvj4M3Rw1BS+FJEKkwv0rF+FbCEHIWOO
0GQ/vFsYFq73+pUk4/8YlmeiRst75Q7+zb/9monJ4+DEMVOVT056Yo7M/BXORt72f1lFJtJmaO7w
02qd5M+OwOtlu3Xsoe57rTPKzmnYys6swDaX5Oxm/q68I2GiZsXi2FGXVsud/+wo5WBM5vrlEFP0
yApQdWrOY8KgRV71foApABNyN17bdM7F8VnUf7wagobqF2k/92++EI0bLzrcSCseP42MelWe2CYo
yWbv/gcQ+h4l6e+eAAjOBAv9h3SS8Hiylb45unC4m5NS0CjeLc83xhVgoBTZpdcGaBGCSt2OTDjy
T5AyQiS8JeB4GcU2uyQbvbZf5BdajK+q4ZvDgE+rlbovppMMsia3fwkYfsBpIUdjUXam4kNvd5el
ak8juzr0z03pNihZitI6ZLa3zSKAyRkI38SpdQHqdBMzX6ts47s82WcWcnSVB+qgSGNDLMQS9mqA
XgZv6kiXVIa6Kpn3M6m9oPAcT5jBqmE8IO+ThVEB2DvqM1j1XxNBmrJwb8pWve/Mp3ExwmwvzK/f
4OKS9BPWttOSM9bXN4iqsd0H0SDURIybQJiPtSiF/8Ms44csFgXkA8BHL3QvCPnC4q9cL4HlajX6
XFDNDdBBAZe7tgT9zXPCoRhHL7tMJemmb0eeH5w2bZy6TepnGAitsII4t2A3/nczN2d3GJWucr8P
VRn4a2iowUru2U/Mu48s2KU/hj2vXrLsP2J/s4pFgwQC29bt8SmHQ53EWA/TAvBvXA2a+DSOlIm1
+555fXz7uK8JS+cvAyLbaz2jEiKnv1fcEiKijrmrcjgUURqhXKetggOkHc3HRDRniOfuAkaardoL
2OSyDwZHU/7yrCKaHG3JWKijm/gOszGw2oBlYkKzII9YVwskFSxwnnRBN/ufA2+Nd0tkfXexO5lO
WM6cXGekrPa5sQU1tH7uF37XFQyVwGFCdjuasKODxS7KdVQ4r2FHY7Dj49I+x+ppjcxeX0e0qjJA
0uqek6ybTB3Nx3fbiiJcd1WZ4CWSRpW/drAeHvYRXkfvZKKMjIrG7E41/C4zBAPK4abI+65YFJV6
puqoKrQ9N0QLAjRbgvhPd0vs+hCxZnrl+2JAISrVUJKi1NJNIekGx9TcwmOO+B6GgEhgG5rzt2sv
I+uHNMpLbPo1LY170hBkpumYEEZ0BbhoAgPK2VHqHit6DLXL4+Hw7hQf2de8ddpEpoVlz2XcGe5U
PmYhRBtyfiigCXdOIEDugXTeFU7N18/BtzaoNbpqkUjRGX6LSZVGmxDtoI3bQj5oSSyq9QgIAecl
JnrYtZDJvzUYb67P+KcvRsDB1Yt4L16j4Bqm4P0HVtkN8UQOYtszq0YT23A7zfZVK+6MUyNrDXeQ
kF/Pi0Rg/GvgG4hMyHRq77u4LKoIUbKrocjaAdz1z79BH6THXEKGO384JzpjPvg6VSxYPzOXT+w0
IQEodrSb/awF9Gtkrr9xUObXcy2g22DZpiCJFj0si8omtWi6M0MH28qKZMIJsCVtk0LW6yvCqGbz
odUo+NrqURK3+dRBGsLYhoptLwbPBw+KfC+w28xdOLaW4ywPW2J5sXLocK1/q42jr4M0qq01QHbk
Uap6qa7uED6vPgOMKcPXbFWzQtBg0m3szkMP1oRZay4SJdVuZ7Gs8j6X6m0g+LfQX9V4VMmclqXR
MJoBqJZJa4JvrzvPHAdyidI/E7uKySfmTThfrMcS/M6vq+QnkprE1F/nS5u8Ksl8wZz25tSepr6N
YRXgQrpuMDVttrCDMMT79Hq5rlk+7saiXsQHTKny0r+jWR162Z5oJh1y4VfOJ/xn8UqDmFQMj2UY
JnkV2cbNDFB8aLZKOVLL7AoeAeHebKi6KIgeKLLWJxxdD21DUwLdT2toyz4wVCAXJjYVysi5eM/u
B03QkJAY8KkxyCqa1k8xL2KraMNauFnmiP+y7u0hXSGBR8i3z3A9CRBkY9NwiERFcjJ0EssuS34H
zJ6v0ZQECDa1ziYWxP7gJ2SR91au1bYsEUWoKKP7DCBcHbSHAfMmjpdSrBLlGIbBKi26kvIOIFpP
n6oYsV3FDrv5xaoyIwU9hCYhgUKXuhEFIJQHIS2w0C43UTXCEihB1ZB8bp7wdkls9f/4jJsj+sXL
H1GDQhvC/RGj2fdokTbM7VDmtJIhMJjG3WY8TKLdfIFsu0zAeyaxx5p+y52ntjlbNdxBiVCneoMW
g4n8k303/cMV4ABBN3YeUUQCWyueWvQ2dq1BysiF2gtTmWn7lOuBDm1q9lWQAxn0ZOnqw0jKHhn6
1TCc0f4zYhQ+s/esSZEE7REU+qEbwUzgq9IgvcczKdtCH3C3dD/Ay8MPRKeqiD+QmNo94qiV2XyC
OjGb1062vT+i2HkRx1VU+MuVws3JoJy4LzeR5x1UuoywHdg98CQfsnT/c4Mm700CknvmXXiZ7j2Q
7WRNOz06zuMyk23pz96aODSj9E+sX8c7ApWTesDFakJcH6SulzvHldtJzozEiZ6+gFTc8gv7fY1c
YR36h8mQPFtVW4xS279e6EwGx59WAnyrsd+z8ck0JyWaI9YuRFEDS+DAc53jxtZkeHhVrdljdpv9
SkSt8RUBqFvLhmUj81W+NbUcA1UY1ZtUFCe2XAs762/xtT+KHJBXJ7VDuaHxpJRsYwxN/qFtjqzx
NNzX8jsxki+rsHIfaf/iXY1Lf8ly+0EchUlp2NTnN74xHtQjZJNlYHWGI1hmgOKuiLZ8Dlo047ir
jnRkd6TGxH4c/J0wlMkoGvI0/P7y/7lVAoqf26swQFPWwauTPe2thHDw/0MqyAOjh28FS68vjMXp
cnIMiK7BOBO+xzaOtjnD2wIUsC/g63Wf2pJ8e0qoLFlkbjK2tYq9neYRazKMfp8U0opHyTyxZimK
qbKZWsT+i7TvPgZkFlJ2G3fD/6sAGTDHUYuuWA6ewQ6B+TRVCnqDx1+VmwmU09d7z90/pZVSJkC5
IOA3z0uXGqT0cG/JtyAEs+bKhuhg0z2sum+eb83WLCj92D4tUKmX6ooF3DoAAfDlR8QaDTJC9Jxz
lTmw+PKPSM7tm88ZACy5kS3uhwmMWeWKV8ZrGt4tZ/MYosjDHt5GpAWWkKYAGjAGVKKv8VQcd3Bv
6LlWUfhHv4lYMaWjFHpZ60BH1xZNjUc6UzSKDC33moE/aew+DqIM6G6BbygaPhpr8vpaADN4iDBu
Kym8SPLkGiNtA394TjgrlrBP9AVBaIPzGnii5DZc/ECtE847l3+xl2AWIZ+vI+BQCvhG+JBNxaWU
ki7dMAknosboQu1tq7idLL/OYlwYPgRRUhBjZ2RN94hzXfq5dSEoUy1ds/CwW7Z+9sDm1DY9JLlq
lI3eo/iVyAXYwuK9O0yMJ5XdJqqQiMPHgh4Y7fHqDFgre9+e3RyWbsvuvfeKyucyDF7ZfOMTQqFF
pxkVFsmhRrNba2kYhjuHOB7LyDwqzMxBTnREgZN/Bg2JtCHc1fKgxvKIKb+IGIiAPxVzdXbSY4D7
HdIe9tTXtiRvzw8VxHee+yHATY3AXBkuhwtHXEp4BjrDCufh2XG3l+tsLYGUGecQiFD+RRlqpYli
7E64gUzO3ayhMC+n6kMTy28XVRcYTgxsWRNw+Fd+i2UKoAQegTQpbh5N+vKp6kyE0bRfYUyVT/wW
bJxgEXRb1K+Ib3My6gim5u0LHxm6bUxHsZTlC/Royq4FKsrB9HhLlCAP7tBZApzs0b3nJvJX+R17
KPoJaiTGJCJ0V7J0VIbde74zU3E0Vet+9g458fFO7QSftvOAkBCXSLmybzQ7Y+eNT7vbI8GhUFlh
c8iMNZa0pE9OOPtg80ywef3QGWLkSzF9C3XllsF/Ij9qXiyxkckpPDz8lft4x9jRTytfwY3HD7Ek
v8/nmb83+VEP8O+c4otRGgr5vc9euuz/JBkZRLIZUW46a9s8UJ2DaD2PEDQgvghs8NinGPbc/nsM
wmxSNAVzuvqaO2827TzSHe32u3fGpLDXkohYG8DWttYL65aNjeppjqz8+lmJ67Hg+QYL+/cIUnWS
2v7Gq5y7ewR39d9HuXQutkexlnvPVNO9IhqDQFySeq2gZ8XBbAFQw3lptdSyh4hRAaYXgvUd4NuW
abOlm16YcCDfD2vAy2T4UG19KA31H059/KayhfkZcO8pKQx66rC5LYqx6bbArGO1TCclO7uIR1Dn
P09EFCsFxk/EwMoIZNK3NeOsqSEJRk3NleC5LVraQ4wqUXE1EyUHqww0EbIxuPxE72xRXpW+cVoP
T1+WDDY15a1gbSS1/M8v/zhRN0vguPcfkpWdgu8HSMmQ+iFHunxHIB+8EXNBPgXBZ3QT/bxcdLJv
snx4wFY7c7gtWtyYX9SHrLuCO6Agb6OcbOdPyAgJ0CWgsJNe/yh7T0oLTpYGjmV4tkYKTXFlE9kO
1tNEUP62FwVj7pWPt8hVNhip1xLeAYKGKqAND1jUTzff5YkNDIJKLYETd+2034x7R50SwcqDvk90
e13UdkA6qkuUvvbodGDreGA7uSxj+r5jIf0bOwgresMkW2Q7YnfZUOXRxhukODWoqts0qlbYIf1T
qTHc3Q8jwIFf8qrDBY54ihYyq6+zwXxd4hAZqz20nGMNDi9th3JgGlhlaNIe3BpoiysfcPy8fLBE
16K5kEtxj31yzIGgss7M0IkFk1g6zeOp1G8SAasYFHf6MtaBk/24DKiHMDoprHuiW15JqrQJbmTO
yl/QdEH9pYaj7aOKGRtQTkHxuB1u1+huigmbzoLcryMhEUCoGxFDiXaEza+5ZO/mEvnu+H1QAbQs
kmmpfGWcV0cw5I18jpZVqdwqRI9kFknJfH8B0ee8/Ud+MA1coWpazdHvBCcVjqxcnSBOUB/OHVSf
w6lr1eS/3KLWP3x294ddZJTo/HEHogY3N3GLANJKGQqJk2+qMzLNAdEaup0ltMZ+Qg5xIN2io2Zz
uiQhx51msP0zjzmIF+xfgO41qvxLOVXq+73N2bHZzIb3zdDEzY8iOq3PXX2CR6u23U8lliDd0wOu
MdYCtvziXfDBl55ofMoJsz7gxWTECQM6VG8XsiXbDNjcfBQAqustxL8mBmGcRyTdWFEobXho4qh5
5SwIWzDxob3AwjOdiwT6yVQMTzdg4Bzd47hen/s/+ouaRWHYE+BBN0qvfXK4HRzRX5SNUAvJHgt3
zZFjHc/JExoQyynDRzLK+bB6M0ji1SkVzS87cVqSJ6nwhTySmTLGnoHY2QHiy8QyYqX8YUTAMotN
SwzXLzMk8oc+saKlyN3GICKy4KnC/19imktcRGn/uzlOLnGjeimXtgdprBR/kHIJrRxtKKXxhRHR
TTIMwLHbVsFRkkmUtvHFFNwZN6HMqa/UgGeOZvRzsPDzawfC6nCraMs9TJDjkiRX4iwVz0NFG+gr
39ICgBqJJ2ZJ+y73QC3lQovZHRJE4NaBqXryPCQ6h/sc3/YDbLlLhp3PA1ryoiqBKGeLInFx+dP/
3ExSPaxjCdKfDmiN+/SPSXrAcKpV9+7yx3Yfovr2sIL1d/wsdAxdVx13Z7ZPcIj2nSo7RAeuJJU7
lNcgn+ZtR6OFH/bX+upEdBaSeuM6JhwsmDP4Bn2zvYURYQy7+9ln2TYVOZTePwmzPmgiocTmKH5n
v+oi8Vqm0Szi8j4luq7u/UO3F5Y+FmEm8zI+izZLaszI3jNJeX1Fn9+wWeIW6/GFGWbP0TMMaNpT
kAlBQQa8k656OR0sOWAgFT5osH+l+L3RYqn8xD9zCKT+wMk88JGv/dRLwidWHMpHfE0yqBnaUVyl
LNUZXrQhuKQaG3kILGlhrIs1Y50n+Cpem5W94KAmqTZF4osUqjsFR93CEAV/G9PfpPSe7ZNKttFb
Xg3Nn+M4/fzBLR+0UyblyI9eQlfMakrVACni4Dw/xkewSynTWV3Q9QN9YahudjwfLpoyjcZxOhCe
uhwitiOmCxUvVP/SKxn5dpwOcrCbyGG9ID8/KHO65A5egna8RaB2l/cktXk0sLlq4RPHji5dg8Mn
PSkOjRvGCVEiru9X0HQZxmVXDS8tIwR1TfVwiWjiAhf1vFD8VnQ709KV7JoGHOvgmb3Xp80KJP47
SftpW6mX2hoVRmjbul7ymfqlUlhhBC4VBwt2dyTTrBe0uyH1ujyeFCXVQMpl7iXyK/vqhu/GPpuV
Es195RJe8i3HnL0BSThujN+bRg+WaVwC3J9mDXo/BOkQr0OWjFm0k9mMbthx+peRN80vlsimVoNS
hYuw1AEn/6QZUsBqRPujkuyM48xHNa0DQS8TSaKNYhuyFaU4LriYw+T6OmggqL7Z7VPM+wPvD/6g
xX6boUNzItGJAxnKlUl3DViXf7IyN2M/YGS+RwI2/wRnK1CIxYRQzVYlJLMVHIhd+mFIuAZJK5IP
OgASxoo9aIfxsxR0PRl0wCJzbpBxGYzlescufq0BtSTMm9iiks7FHR6NgdfMDcCE0IP+SHMVP/K/
/NBWm7w+C+WoE5ZG5XXLq2ZPKgIQvHHoV86DfyMVnV+rWmScex6ZcA/XbTVbY5xYX+EMM5y7vJkR
FHZaNvflI0I+9hD9goH+k4Ahxflnh62BdWokt08zu/tHei0RiqKGGNZ1WPYOuJgGCcteLb+olqkf
b/QXuaEBozkKtWoWeyVPZ9tSYfRba0nwi5UxrToIjEiXcvUzHEPalW98trJ6nBY6g0wURxZa6MNT
xYAvyPeRonbTEKpwi5edxUHeBwVf9ONH854z1lABeJVD2zrnMcrR4r4nl9TJF5IAdQ31mwe1C0ox
WnECOVhmAn1uzjdFxtsouqnM6JwU0YbkVyoLjlA6118+pd5YhFYpmYHysNIlCVKVCrJOiFYo2Dnc
PD8Pm0X/1ONRYLc6m1v42pCNn9xHgF4E2NKWgAh2aARNUJESRwrZ1eq8GGkqQWi/zWCqzIYsqMfa
9O9xadnGmTF7IjexjdDiolnXKgGLoVxy2VVr+5t9qd3lHxdt51jnjRByFwFqujep0AkO3QFE4fQY
3L9du34UxDDp59yLIcGsY9mdyapd/07tUUIedINP/JwIxG5oTCBpyGDAr2xJC4Q0EivSBW71VAsp
m45BeYOKTMBumtz2biv/nmgCc9RvfkGZkv0RCweAwbsHPngRI0o6fISLfhyGFFmeHXfyv9eSZ4Nq
lTZEYVKGxhwgjGdxrSsC7a/FTBSHsoo/Q3MfSqAKYcH/H5qDJke++YLjNILjUtCGtpm5Vg1nNJPr
PPr2TjJ7CJtTD7RHySAfEpp52EIsygttF4ME+S7OC6liI54Az2xDaxgUnbB0FcXEgDxEnX1FJz6V
Zq4I5VMfx7pvUigLv1SU0Yi00k/YHc2/4951U/uGGtWfmlwhgWDdY+/e31scb8gRJjoiH8YdsBzC
bfcOG+q28brpgAg96z5kvyQxphLaDWMSx6un8sEy5yH0REOx16zmbUutDlqLqAWN0gVpd61EE4mM
eQp8THI+Ckhfvmh7kV6A2xbmoOxWofgpp92GirSeSQVuquuHWcFKKoLQHxhSyXdBWfDedZA+Yrt4
xwEJyeSA3P1cR7tEWEIkZRcgOEHyZjzUw1C0eHI75cGbyWHvu8YOlJd43pEbS2yFw7jFU8D/FSVQ
GBhwAWUC3kpJOASspvAxfYCR8rRqaK/CyE6JjPbNgsiS4fiENl/wLfIWcygF5hiDjYZkrc/9jLz5
pxFazri41UVpvDwtzUnmGUCr+VKXxSiNQzRq88f6iqwxecDKZKSaRvZayzuBXtbuIGar9+65NRy8
UpPjj9l40B4M/GM1X1IHvB64vrZKXF9gsQUV9T3ePWr3N70t+s8wEm5LG4+9wEyRPbu7+QZzEkqv
cuo6Y21bFqyk/lHeu1uRMTg/nUwkwBSQq470C85wql9u1LRYvgKZSmK3vVZwHRNgAMHWlACcXnbV
MVd6Raq9T4bBT+EG3QbCmWP/nmkgbKEb7mdNGmrenkVkhIKX2JDXsGq8WgTFiZDR4BovQLCU//Wz
6yS8hl7e8vwxp32qr8yLho3JBqmNJUgjB0Hc55e9jowBJCRzZ+C5fkZypCkKnhAyKovtSVYmfiBN
Ky77XSbDASexMlkO5OXmagVuPqdkukVxVkRXHCF2WtzvVTJQmWumuaL2ktvrOEFOJEraymLIiiYZ
kndFBnL/2r2TRjmKllRZRPcMrRrhJEzf3p+e4YZvMc4phoZgUOz5MSArpUAhVcImq00OoGHb9me0
jfJFwv9BzmkEAgtX3ORVnuvjOWtXFBmFY1c0KRflEedQrltt9ej3GfIyU0NkfHnMh6kpXKMFCrv1
8gonZYKlYbzeMuDROY9sFSLUs4NmBG67wYIYWK5wfrAibPJl/8Uq9BRL6M9AXm/jVYmEfgyiQ70a
vcBAXO5h6O/yqDogbNrznwvAszepKYAALmoASM8ghKZDBaHa6ANGfHodnbvijZVLfJ+BNcCl/URr
xU3rpqt6S2qZpG9kLUN1ifggRShfOnY9XKmlG5xmzBtdSqtTNTUvCJvuMO9y7Uskd6L1VxOb5+aC
KRls4eJpz/Vl01ykQpGuJCsa/BoKD6Uen3EFXJaFZeNaPsO1IeKD++36ypX/TQJeUCIVAbI2+J0I
alQdUtVjSBqYZ3HHHtDMGi4BOIjcw4Bf0QUj7LAj7M6SB2aRdx0cxnVvZuUawzo/WPM8Apexre3k
DaEXDe/GGI8Sxo2iEoZrw8iKp8XM20oPWo+LL+QJ5PqpUlb5z18bnAPr9s3hqnp23wao9CsFIyd9
qni5yn7XpdUuVSgVLLIKAAUvUSFGr6j/7v8XnXhHxFJCat9NtPCRm2wT7SFJ+LbXfrWFbJo1lJ5K
Ti5bOmw0fcq7E1Lo1haEPzZf+lu5+7KTCO9Sdu5NmDkytdxNhgGiKfGfyB6u9scaqyitqC1F/7Mn
8VujStIPLdFfTmJdEqip4p0OnGwRnp9eicW0YQ8ic0OIps/dREB1bBSO8Al3tRF0KxqqCs5PNlnm
JSP527V/oLY5U+BFdAnbBI+FQAbgOsuUn76as3bg1e4EtURB5V2Sd4Q+BM6pj0SOzcLgVOqlj6/y
NrZ1KXYUPkte/TM6a3IrgNZuX0ud/AeqDK5CbeRVV33FADoWIS6gZrcZTLSWiHW24WtTw4oSnQrU
2zU5GHH8FAQWfWYZWReUMRg90p2pS14HwMFlzZVKAtMrbnsNXHTbs5wTbkE/ceA2m5iJGxbLBDwP
4BbCfX2CQewnaABwNAz/A2IEY8YaVtskZBimaDYvdzBNzLvj5c8Tqail91U3pYKsOXt0FsJc5wXi
mX+6fFtu1JlMs0foDHnMyAWbnQSx+/9c1iKb5drBnA++DLkaIhXcK5ib+m+2dfyX3xQn2mE00FW+
oa3faDT+MHZ8ceylSl8gxPvj3CgRU7BRgrJosf9EMDs/gWwtA1wf4wwShXhfnqUff/Lt0RFekiCm
q90Cin9q13fyChqTfOkHFdVWov1cA3p2drx5qgGLCVJh81ZIyGIGFI4NifQqZAUAmPFDD+7P+wz1
99KDvEqUrnEjZM+ZPv3Qd9k/yQb974ksYPWDop0ZBu4rcJXsPdckE/PcMI6l8eWG0NdZbE1aFnMm
+J7LEnCaWMurjlkturdsHVlQqPekCn2akj/aM1KU+SfoA3MzKhK0w5mKqDm3A/4/WqqsbHVlnVNb
IrzmQicM1pD+BIqgxwLN1OdWFBbgqj5hIsVueHSE6u/KPmavBWSO8QHGNI3bSoKyqK91kgfdxqwk
rMPmxXtOSoJ3diULP53AMdVJorb43SoNfai/o+pF/D2nkoiTwGJqaOzP5hcz8Gt504N1ftotu8XP
toR43bHATFoIrXhyOIWqaWjmBPavasQruy5rRQGZFtv0FOsORLF0y5zGp9wiEd1jHuzk/V6TDpzY
W0phKsDxX/QKOoUYJ878oV6NiA0FZEDM0zQeXWrBWzcy45GJUWYqcD81W1SVJ97Jqm3BuTVGRGI2
+CS7o/EIJGo27ziFZ0w5E8qgIgbOTrir74S6WlpKd7mh8EJLXmdk3k1r3wgrADOdQklCusrNv4mG
Of6XT/mKUG0RH++x5UMtbe4jmcP8Dip/NowwnfP6ScFPxkgvbmoHx3qAmWHyAmrpxY/ejnnndyFO
pZ72NZfNYrkSIUB5lXScHwVcw0BBLMv1xDv+TgqbG7azTxJTkwBidf6aPloFP4yIvrot9x7C0/jF
BdQEozbNW4juoDD+mqLCq/7PRCRMVFNZrzIC7pMClJvw6NX5ZxIyalD/iiuAAGXL5BV4cdfUSZe2
u0Fo9W//lsFTK7UGkMKrrDC/MEcIUITZ1q3xHZ++CHO7lNcOCnH0831aeyEo5y+ksjjwsJSD8WXz
HYWq1591GBFTovCuGI6yalTYLuEpUnvS5Phj9IbDR2R5+ncnDxs3fmMoSg9f98nURZVqRoY7dYwF
uU3TCqqT6Ns78jCKX2A5L0YcXxPRAknppHJ3qw4tQMfr7E3INCROVrL88QrpgglhIIEK06RMZmWF
ALqUzL4e7Kna4oKUF2gJrAxqYBFfqox6/dMkjhWjmYaPg8cR4sx5MODovdJJDA/aZMI07BtX3hhK
IQcXF/6fZjV9/IcIQWq61TbP3KIl18ipztxix4P3YaJv1VsfqBgfSMTQbs+hEiKN5giSFYKSF1Lb
8kfcuDwrKWHNdrEJ8LHurf/Z5M52p7GhRN9RIxui7c8BG5pLPNbM0XHJuezwuaFdq2x8GnkC/Eyq
N2VFC94qh4Ek2P3otwcaBgzi5tRbV7Odn7jhDFk5JuzTWhYrvsQjOkZhkfXa30T0oPYiC8ezez/K
JC/woVObaLOqHL1ZV32YgXPg4XsNFWSxeY3oDDI2cPr620iJZhxSCPEKnOSHheXF1jKdz13vm7oM
Ay+aMEOywMPrA4uoD8IXwD/a0gpif8B7C5uZ9lJ3TpMD2fdOlsyLZDQX3PuBquhY5sA727Adcy/F
Vw3KRPIz8BwLYLSkEM581A9uoI2EppwR3ISjnMLqCB8MGokcIlfSJlOxd7gHQ1M6sngVIBYs3fwU
lsPDx6fQjcxSSm1jljBhGPffl2IJP/iExBP7FE0nVEtGBFNTERmfsvr37Rbu9GtMLMMn+ciDP3JI
W1EUDNUxJPxCjjvU/mz9FAUjbPM7FfInewCvFs4g5MWU2TnvHOLYfHPxe3YqRzNlqFeAvk3Zm5Tp
WvVxJWT92stGIwOZ4Wbd6tuGGL5xzI3ARzdeS8eR6DfluGZAJl6a8ZySohHozA8ZQxj/B7SgdaGl
B+OWLEi+MGbhwL+asvyBQVRI0tUIFQc1txB25KrhP/ruk98WIukmyklNbDsnR17oExdRjaZ9xB4O
raxttADWYMEGNERwbyu95+Bah15E+Kib+aOFs6z9dOFaHJ392CkQo9TlzjuEqCjfc2S+OqjPx3lH
WApS1AmYusw6H7hGSy4x38PlXypdv10X1OWUyAIkuWQBMDM5/lZ4O9cMIbuIBM8ja6zOUiaSqHYZ
vGF7tEe7V/b2UWxgM6UGljsjcRMpa+x7fw1YuI0dmpkQAjaokhq6M3fG+46SvQyzXh9fhhpJeBNE
72qist92e+A0Am+cKcdc4KYa5kT8I+8FzT1E8X4VGCJudoY/c5m7U+UCL9Nce9K3DMPo0mZYlaJt
6a5d9tqnZdGRr9PFI7EgrFx2iNKGbbRZ8W60DAxHmBXuH3R2tl55gWyF8kz9Ts2SC4oejYrVUzQM
8MhJz+MaO1/YJXu0mSjXaE49M6Lfyn7KAt1YSOGZOKusv0IJhuIe7mKP82tStnbNyWcQ0uSBEyUp
7syvtakeRj+6lOn8q297u7aaQ5bWjj7/SvJXYimAMZS9i7SrYmCsz/1+QmLZr5OR4GcBQCO6d+IL
Xjix7wYIUe+eV0Vmgho6QjvgdRhjt0BKtvU+SxBUPwUkEWOHKoopKg/zZQwrfNmb/yuw768AiLar
tlvC/1etiiQiWEV1LXx33HoHn8PUAUuVgusL8lJl5fKPZBv81wy8rIU8jBech26qGIL+i9mhxBxT
apqnSR1WQgELTaOsiAqAQH4mIppHs7SiV9Bq3/b8qTrYJs2JALG7Xv1bo2k7RrH/AWdhI+jetzIa
JAZbDq8GRh3FlVQfkUUUN/1wydnQZ2u7XVxa0uF+aCP90pXvjPEMxi9bnMSRwyhlAvtlh0n+UXBw
wPR0/l/oWOf4af0r9LUXx1l7Xj5D0MPoQduMWVq7QPqJ5k+MRuVRkMeR0Ig939lj1wVEZZnoYUDi
9N//2tSZL9NAAH+YbNizy8vI7QiJ8IvVK7ALu1VgRt5PAXKv8M/RWD2MI01bGTxA5TVot7eUbkwr
W6JsOmnErrb/tu6j87+srz4cD2IMBt11y39cBchBVmjsDST1PudfLCoI+vVWAjbSfvjz8lplLSoD
liflu5wgjbp2O6nJ9y1CMII8GQjQp+jvfBWj8hA31Hm80w9LuUizd/KfDfRFe0FpaAxdz1g4meMc
S/qmCwpKHPg9mma8Kwd9nQOwXR1Ub2dykeV03wcbGI7jrQTE5iCQeoL3RjWgSD9GoZXwJ0pJrkPC
VqQ2W+iE+nvvgBCvFH6FeP9XPrxHtNWp59uaVTSbVfx3R/K11k7pgGrZOqWRknl5UeoPSqhjsAm2
0PsQnl5N8xL97M9a8STLMe8Qs75yhcMdBQHJUMLFltmrSQefPbaHA6R6z+g/b/4pJXJ8nrBowK2p
ssnsONi4bYxCcGRCnFU/x33UvlwNBUPqoDw2OJ34WMQsvz1sEnV2p9HT3K4Vgjsozpasol6Pz859
G5Yck6u7vEyjGD0fmbumWVwZ7u2h2NW/TG46EN1WnA5BOB4kcDYD8bm2kTEtDyz2itcWOD3mk5Uz
Q4vpDNnJi4zpXAk1N805D0cTSg5lPctGCGsos7GWddAUyyTjSelWP/6wTQcsFxZK6M9T7OELWVqt
dcRbeWBd9CsWZsdKZMmzKPg9FmzgrNMnDzRYIeEbwuEiYSaSNBSl/WnhYWZgnaaiFhhzZy4l5nNc
8cSEQwPl/7HoOWGlliViyOZVCEJLHu0V0RJK06MLb8u9IN1dn4hNyIhrDUIe4dHNNfW4r1CSBcyQ
+3QXQcHO6ov3pI+uHQygJb0yCVwdSoN1oO4jgTbgb8PdNDk/oDO3XRDO8ZmsNZUMHpkDtrCwLRnu
xIvuaWzTKKzJItwSAdA1o6bJhbTugXAJ9OFsdQDqLMAIkw4VxfrUI00Y1qAFqWHgd4AHLgkIXdGT
4uCpyDtNRKxlOr30jMeBWch3Bv/v53tGnCjUo+pKpeRJ9W2fmDM8a6JMWqLhfEEtNIhLgTD4lgSn
pFpc2Kx6CeVwUjUWtmoW1bR12/QmR7GvmpwtrHjZz9qQc43NejKj4D/zX4Cc/CEWLPE9zxUEooEd
gIRvGbIFWHnuPzIG6P6o+DtzOBlotH49KTl/J3vTslMYXMs0BFn2ZYa0oVuyToxWXUCaY75uk2Rz
gOPqddVtmd686dycfezd8znRJPiCOu5yM3F9qHJGXra2bVd1cbzvbS+VGCqctq4uw2X7chWBNnQR
wN8e6slYrWCovrOERExLE2ynV2A8zxr0cuFLzsWzv9NQ20UGujQUV51ufrxmLli5E6W8vJJC+2eQ
h+IAVfyuugB/yLxL4baZMdsAJk0a7quyQ2zjfht0O9hR8SOCzvVuUsTmuHLd/xn8deOFyj/qr9wS
sruLoX9bWQSPAlNRb6LmzPqCb9D8HG/xjoSS7mhAcqgsO18cXABeACaAvtb9WF60e/A4Se0VGKF/
QvGGeTEssRx+V2a070ZuPq8mAsd+hqrSORRETkSbHZulL28ujhlC+k3RY5btcqi0K562tztS7l0v
tiExPq3nuNA61iqiwHIiX3vqfqSzBiCsy1Ecl68bGzKGPiuw5U8qh7TPAH/1P0xvW22MJ2E24QfG
xMjqNAJTrZfFpGp7dxavJQE1sojHv15iqQ4+Fz8YMHxaIFlak/qEVuMl/hvZixQIB8GrsvGZOoRk
O3KWPEp2uxw2zFV8inKvP5jzvlyjow8fSxIuq8MatEVUOMVb/YoWJaRL6ompKdH/fYUmkz3VWJhA
DoCG/KkVrE9aENzUMaQ4W0AAVXd6jIF7X9kq+0XPilM5PpU2L6Y8me/1mQGox+zUO2rVopz1YpHA
PjWMlkeVOoHUb8IVS/Ov+Yt1uh65izgcZ5NA7+EhT5v3bbNDHkt/n8aO8sO4YXo4SoxFPDoqMRzT
VoZ9fglk6qD2dAewTXPbjhOv3jD1WAMtF/g8YJlXClM5KkAn5qQ4h1J5OvquBPbuCPFw+dqjup8l
cBO8tS1fKhEN/peSelR7MSiUzyFBZJG7zN+VDGX60JWjckcU276RVjruN+lwjKCEZ0y7LTu7f2wZ
mxUuMAPDh02Ss9awrru1wNcEojdlQnD1jxNtwDrodHc73dBloZaQK0UM3EzsXA/qe912QUhs3Gti
3FFPgYbLa3WOeoq5DS4Nw7mwvC42hwii3eD8v8RtomhZF2iChgfnUGx0Pmmlov0dZzpkfi+icYsf
IUntPJOlvEGvQC7sSZBEXvATqpie3u0ti9bS6ueo60zIFx9u7GJ9a26zcmWDemdJ+wAsDqLeVPNU
hSKlGyTkbW5rxOUld2gf7SbGZJ3fJ/EpLnQJ/e+ccX4sZxd6wlZ7a1g1+IOtBrXtAbv36H3H9x/5
4iTBaEdDxwq5DrmHPTbM1cu/S6u+mz4vLk6NvnSBUuZTlpj2hNhCMxmeuF0ZeLdyePGEF3l3NgCF
ySLBqu4JwozUSJKcWtM5bAdXZr6qaaPqSEqBwPwA7kkV0NtYp2BRPsRyDoWJOmCTn6IgU0nDgCSu
VXeyiUDXUVBYKIEw34A0rHNTdBi3Hee6qy/WJvrs82J7EYmVhNW/MZgVzS7LL+086pIsZ/O3GA5o
QgBTUaVMTWG26q2WThXPfz/G5Hyfd4xMsOS35bwT1d20J4xwbvn9QxlXUaGYMRsLp69B/lq67hf/
dJOwmr9ZIfUmgmLD+Eim6IvOWSwAHzIKGD/V/ONhD3thEbYvq9W93VPKDKLJdxVWWjFPDCsONZQ0
XBUhmfXKZ8q+iQGaoV/lZzsi79BQkgy6u/CLpYberyfU9VK8hSI8TTedseSzXTMdXTKPK311UWtL
OkSz5hvAcccSl327I/NKcUPSw4CPqfRD56ETaVOuwwCiHxlOf1vso0MjaAmmw2rU3wZj4GIUBuhN
yDENQaHMUAsCBSB8bzZdWE9vr+6R9tWdB8Tb0ZxGAYfO8f6DdlqbO4cBZlA9N2nkgxl7bo60E+cY
dM0fQZ0e8FAxRw0bksJwDnU3SGtU3VKxSrP+wrBJgZcVl7ZZ3KkqPtMgRLUncs79NYJu8ZzYQ4ka
7l4007Z/02lXFwboeIfqiU2LukCcFtDf7L4KD9MxSjH8MFsF6oIthTfbjfE4CXMyg7adwamVvY7r
HhhzbN3Gz+pK8nsyyEWHHonDjIR5+EyrvEOm8+OYnr+yzh3RIsvnnhWt4z03ASqnGTCMe1JXarcT
MgTcZBFi1AcQaK7JNkclebmh7HApb8s53th9G3BM0cXaG1hMAETTbHMaivpNJWAOfsxcT+kUSZdb
vvkBbwLuXyAEwxzkkFrkc1mx7UZfydy0wVemx0SqanL0rVFVrNl+7RWUG/LEVxzMAYgIMwZFGSTc
lefA4BMuzCB19ZzInUUaBELqrRD7xqXO5gweZFyRazCfjkvgFYIRa3vz58VFR6rm5aSkoQK8n0sS
x/TAL7/Iml6Vy3rov62epzWbiEybv1tPA4uqpXiXv0VjO4ytjD46H59FSOTrPESeH++rmKKWFHtk
TZ5JLxeG59fJNpX3CsRROZbHXbyPeB+wjlVUw0t8IEOmFw6iSJppBZFrmRU0YuIhAjfx97RxBGcT
hZGdzmaoDvH/fHmyAet/2/0j8UDYoXHnuwpl0wrH7LpZ/iynwAY+ZitzgWnXZHa9/8+bGWfKQrFs
0L92JdAsG1G1jpMdGhil1JGuXTHkyqdAf9lN4JSJ8iFJhKKlL24GXdK52nCs7l9y4TLYAduDwlvQ
RVS+BwgvZSLLfbTBx1VmnJYwsd9H7CeZMSl3p9KuB+42d6OpWwHpSI4KxuJrwNJ+tBQTm7kcJI5e
q9UZTlvAyFSBu/SlsLQ/BB97We7ccaX16QFa4S3oUDMVCNRvSmcZydnvpQ2FQ9lqYIuNaQEVAmP8
r1TcT90USRK+Y00znsTDvNarSp1brcOqSo9K2ciERyWqsWAcpcGhXDbv11g9AOHhYRIo3Ft/Avco
4dMh/8ud33WksrXAwsrS2DUcawtmZu83P7f/Em3nWTbn4tkGxHGV7bFobniPxNYdYsiXcXasAnTi
dUXtVS0MrXA4J5KpqZhfrJETFZdvYcvjt7O1whp9aq3t/R2QTGZbz3vYQ2lo216B0K8eRnW0x3Rm
N4/UH61kniZ9SKXco+K2gtMkgksb2c9k/GaRl1XzuxN/rRlqp88vo14Bt+HG55+R92I13JNicIaX
XG/h7CgL2dT9QoaRtLtxxbGDDDk+K85eNwKuudHUD4AVCdrOIo7cZyi53eBUJMIWd4yWpRimCT5D
M6VvZIRT9YmKvmYD+RdxRyBqmsKARVdfPv4RLuUTBBM9TUVWkmApswcYhm7mTFWwLpD7wLrzSiqU
+0axjzMD8U2PzenMek5W8U8Dy4wQKLpdkOC0lXwlYFqZDGmgxSAsQzhLlc/RGcWHPG1ZuJNq5zDP
1jtsNx4PByi/HsoVXYTtFQL8AVGRI4sfBzN8aDWLFy6RpRW+LWBdkuotuYfB2r4dMWXNtd5AfwcA
5RPUcLOUwir3XqiRopayBJbzJjVwmPaOVneDqkKyScmMy0BTs/LqpvYHrAICM29+K/U2Htxr8Xhf
ZlANTYy5qiQk/JUyxnbD355MjQ5muwJ++K9hjnUuMIJ6DVwnhwQl55umAPA0z5HYCsGSU4dL++Yp
KHUloS0el1CzddO8M6xaTHbT5b6CsMcSzmU3GTCG2Pcz6aeGROLdfrRast23ok/4jNUX/293UINe
yeQMIXGpDqzxuqdFiRVPzFRfcGr2Du6CKdneUYWoxdwEMJR7RnEOTukv0vM5cghznqI/H9rOHeAz
5WpxaZZn0ok2WxEte8a39OYdaFjpDsJrZFmNBhLq/Mpj0IjeeT5Rv/7HRGHfCYK8VZStWqgqfwMq
yFyEexw3tTcj6B7ZqlAMBkeabhsr+h6kT40iyehWceUD9RkIFlCUUEjr5SHkk68Q6ajwfu8MGBY5
X3cdpfB3D71XmPo4QziKaWHqAxE2c8TREF3jPHuRylRo1uCBSQpbnqkp2K9PQhRROh8KAYE3d4xi
cz9ea2oJPs5ADb6TyupqmT1oyIAAkP+zSYdNaXrk+rSkMClV9ExxoX/INwHZjupdatVG/2Lj1X72
sojXpsu48+ekcCQWjXe/LBeQKL1Z+vkwacDvVv/weJT7pT8jQnTbUGFxtCUTPOmuVjKVRqWJLf7P
xvy4L40f3au6B63YkHPQDOfsE685j7ojeL0185zS/2SGFhehv01eVCZ0/DdmVEbcr/xx1wYAwzwZ
ylQf26JRXhA9l3ZkLkFyS649+r+Y0tjBbyxRao9nCllhWK6bqWCNKENgGDBP9xhu72tstUcV4Tuv
5clnXiRi0EuJ2ZI10+/T8xrL47dIvAQ7cNCysKtAZ9im7K3B5c9vAeq4xSGTQsiD960swUR6CWej
xZw8+B7nhDBiOrO/NLEO6cdd5+Veosap5L++o5+wr8zkBNMmn+2KfzhrtJgw140/E7hCvfmN+HL8
IhLs6ulcV3+2VZ921QfPAcKv2u+LpRN+andx1BYYr09ib4Dd9vScBU+4WQekgkJXU0IUtmm9eHKh
mdnhfbDd9UBRSb3VMpGQ+Ci/rU4SWDOWEX2GML1hMdlt35JexDM03wW2YgDDI/Icm5+cgsMiIy53
yTK2zNbkmF/D2e+UpTKaVMI0Tsn26USzW44bt6+rA/RvY6HXvVuuSC4d1nsSe0Ya26cJcJHcTYeU
tBbAHjUcDPqZDFPGfm9vKgVuV0G6Hehr1lY7ZLb4exGGMYqtudkTGihVQD4Kz+zc3zG7Eqxre6nO
fyOkJCzVjKaoDEa7kjNninXC1Gy/YfVyvnEyPi/PrRaxlnBrSsrkCKoQEN7dtJaUkUuSLZeyY4TK
x4ilvEICgszoGEHE/oko/3x8oz/8gLxGNQFvRXCHZ1lrdm0/DETgp3ih7PwNSf0qmjy/hNa033Lx
9mBtZ/f+ZgqYT8KO/O68/6CsxcvJNISbjC4pAxRV18pHFwKUISUuWLXAdcMXgaEJ6izHbK784Fkc
TS7p2WhgYM90X/FuzNuVLZ+iUp5HYUeTgJOA+lQge6800VihRsThXaXCcGeYivZ35tkMQgda53yn
iVVO9qLy4Tkw9xSecxa9dKKtzRRBNc0dvaRV48eD5XNPOFqHx/2ZOh5BQMt7AyLY2cK8XZSIfFbZ
QYocWvmcMK98H+gra/Jz8eXbgChY/7gobB+ur1aQ6BQFP9TPKNnOZOa818yTH6PwJ8qEPmPZ3bEH
jweowJWHaz7cCT3c5WTpP6NC/9dQoOk9LwxYbA2ns+L6iNnJD7Uk65TzuFjddYgDlV/fT8w+0daA
k7Gw5uJtnn7Vnb9fqfwTe+lj0uL9H82wASEukqotxEpdyquTzEsR5Nq2RRhnEAVprSwixfisdcqa
QdT1KDkR/qGijLUjV79J3Z/UKDLiv8M7RgbOO2JmGWnZUSYIjryLUWXJbeFgC9BYKnJjVZPBac2S
UeilvQadMwSCa4MEBr0FNgr7tjIXJP+FesVABYf+3JnM+ZuvPaOxMMWxmzps8fxy5wDhxFxCDMEf
Q7XJ4WIKr0QSkFWt4zxTD9oE1gYekW3vpvsrVzoFDLPV7Xuw8fhfcJ6RzYkm7TUUM8EUFKpKUiSB
sQqJhaQ9ZnGqVCdS5AqtWxKBjLmf6KL7+25lybkpjgfWlNxt3FfipgsDYRl6rFv5lF9ClnPcM6Y/
7zoQDfaH/5P/V04rprktsi6KyJeZwLmTv46kFpBdQOssifN8rKStd1vraroXx2QH78eKZeLIKxLb
9yMdqD5FICJZsZ8T4t6bZ2JAntizGm/Jj0xyJFPEtq7wfNXIGOYNY78emx63mVqEcMjP+ByBHxIF
cLlgMRvo9jZUef9YWiqcwCPAQDFbltG1W0oJDDJ0KApPJfxVd1XR7PAq2uJUPzoBoWPbhUKaKe9Y
ZyEht909YvOkDlOuuGAQA5L6noj2hZlJiEbMfKSZyPey1K2NxP3F9HSq/lcdSyFGQWxghtyk6FoX
fb8RU6KbM/a1FRYbS1ACzr1vmKl5SuUsqEQYj2i188dAg1QGow++MuFs+SdoHr1XSZpUAst68qc7
RpnwnF3rO5TeoQObEZmM/AlDIyP7waH89I2KqWFSWT3dkiAFef6VM+mKCoNwF6IDXPCthkQtyFEr
2LmdHIQqa2QQsNqj8EGOJkEFAL4KAwfWQx3intPdZKH6uI+of1HqE4gvE/qWutqDxNJ3A3/fHZEU
gtrQ4rmLmOcmvJwfNzpxsifEgq1dHwOL265TKwJ/DvL4Pig34Zr+jPBFhIh7lVZqemf/o/QuK1Aq
bFN6tKm9B3umwNo8IcJHDDiqFFvabdh21m8AGqsruvEBYruA7Cy7rwAFLIRRhvIMIbZp9ip4QQ7x
e5JbvaWR0mH+Dp62MTWNa2W+qU94hjZ6qjvT+fHFOOfUITRW/0SY5iDfc6O2SGeYbpIKdmGGDwlC
AMqLRb3p6hUG4J224ttAqMnn8KV0Dq8BmG9u5HwaH14qMD9rwQ96k/esTtfeqmAR7iASAL7tVHrz
ODpcAZfGrQTMI7wOLkCuDarAv+1z3uVXCrl5lQzBcNj+OBh73a3CTV37JvpDsLZ6q2JSlLrFKkDV
sKlfL/3DoYJcY20x69uQoQWMAh0YG8cNqMOoKOQ3hiPeX0QcZ1O+H9rpfClZLEk6qltHjGsFiZY0
BMPslKt+hhgwpVrT5faLKzvQ3q7vTm7i/eGCJzWcVFGeemAFNlc1Ee3ZU6t2uP5aFierVQaJJeAp
xgHiYwcYkd2/2iyom+O4fs0QfLId+tfS9TDCtrGD239T4i2ekLRgETvad+8uSl14irFgPqCU7UYn
NQcH00eR1NjcfkdE0Z4cwStzrWWnK329WyaXtHlIUj4iCwxuuKK9RxHTZKmi3pauR3LPWjXXbDWe
vTYHgI5MVTGqDX9uGY++1JKv7V/9dBEd9tieOMfGZzVHCpbw2+1kMQqVaOm2DyLK16U60/iRq5KR
1FTMhKsRgwcG0hfYS/RmownudL1V0w0GUgapO4NND/hsYz6BEOBNJ0gJtFXi1zRNKvVJq+qe6fln
yQxM/eJCJBlYvD+FS0QD6oAUF+E779xBuCVIkVwFdDvmfu+SfeNMJW0L2qQgE7zZb1Q0u8aJqAUd
i2gHPePTiaN5RlFrHhc5sRoz2Xf26y1ukbazzjXo+38gq5kv7eMUM7ROHBoR2j4WRo81JO/hTC1F
s7JY8+ORGeBWzFKqabMG2WRbmYmngYgvKC6ctyLBQjj+kRvz8XIq2gtiUAh4Qlp1wXrU/59jsBlU
Oj+Z0usaJ+yUFDC+nMroSsMiENJAJeXtyJSt9buICQlHy944iels9ZXRFkSnTCxXNq0tM8begI3k
MM3ne7JNz/rblQwh4Os2yeSi5AQXy1KcxsNL56jFUpyMx101M+D8TRZKwLXbMHbWEqZgTf3wTOwS
Fn9oD4186QRU2inxt6RiIQ0h1qVd7ydGkUixhlm6T8KdvEue/V+IsnIjPlriRWKdfU9hCCrIkxan
V2DFJOYNqBNzkkzd9bQ0FVSCdnorJIOdmjmvYfRy2Tou8cfPmyqjiBwa1uw/qlTqMk/vnJVWgkkh
W93LDnMr0GteZEZzlRWAvX8j8jjTdl967E1Y9TUjS+ajtz4kM+67EjTh84ejk96PIbe4t9p1ea8Z
iOhu0w5Y9kpF44JOaxCd4D6fzjpqMQABkvf033HJ7QadbAT67LbZlmeUuBkfj76yi3xbAOYJw7DR
XLE9eg4K5uwPPz/qbLEGYrA7kaRzZzJlC3rM0MQLZjOT+aBR7t0m9apKuvVTmJ6Nwm5u/HOeArzu
7v9Ha1a95S3rDUtow0PdJGRaZyN6lcSsgloKV8Ro3mCHcM1Bs9FsqMQ8Nueo9Cc8O/RbRjFtTVuG
xfaqFstJ66FPKP32LEYa0XQbdC4O7a0GPeitLdyiS4clHi5vIWlYp6wcxvEqGxF2CqD9ROXYO/Y/
x37xs+FkZhwe097dUlNqU6gBQDMc5Z23BJu1hRqhAmZD2qYjlHqoQWkqG3CD8nM3Xfkyg0QcaBbj
tCyElKUkJqiKt+gsbOqUduc84bMoero8oZz2JUueH6CU+Xi9EPFzxmXI+cOX6u5eA2yh7m+m6rdv
k+bfaS40zl0RQP5uIEe/HkQ5j9eVPptZwY2kHPzqAncKuGoQHvoxqwF9RMELjnKe39s7yeoEQ/+k
mmFFrwub3qFztqw7p9Cs1zsB8zevLVLuOc07jz0e7Ha65T9eaPzHhbSLTehxZ0KUhlhZyDFgi/Gz
pVZwrHE5dH5mEDJHKynzzczRpr7rknhgFk+cnVBXBa4LaS+LcgVNMlGWhIkIpVYfhxwvBbh3rzNh
P49N2PzX/bsQ/11z9WkEi7wF/lTlYpZDZIdEVvFfSoywMIn9dHuYcZOg4nHvnnLvJahaCfvADDbD
faT7zKE/ie0UlDHO3CUSBK3Dl1q/muqErNvvwxUMziLfNww6V4/u5oYKgCrkjRd/vzJ230q2DtaP
qFTtqiSeNFNgSCKUsLvRZXpwFne5obu5R09XJfZspY+1mXKkvj8AGNN8TRfBe16A94ftpdA+mhxY
uxGFrfRh6Y8MY4P209vGvmCPJM39UwLbNVrB+JnUp4UOjWvkdHV6DsC+0bbDPRrYrakmO7LsbYB4
D3vbGu2kUa6y3+2nEHARHBCEgn/PGHW678mzNbnue7W/3T5+l0w2vwluHTNxsOc1ys8P6Q95duVf
fv09hECmB4h9Pvx3lByus1dv9cseHvb/wqx2YQoJP3h+mBs3VkOPTqVVLMuTfsqsIGBdz4bvW/P8
UOvBY9BDV4c22ddttABK2uWl7nEZs/d5nBWOUyQwvzLNAN1foOOatljoa48d30VMjIaY4KqvVF1/
hR48rny2fJWQ8kV6EQ2n2Zip0yGI0Whlck1dlg9G/CtupCymKFHiLmhHbdAi6QY5ZqDe6xMOC+fU
xJ0YleZj59Bw8gnH7aqnoaIgA3ysOHt3RJp3bRee/5ELuU6znpLK3/jup8w+4WPoCqyS+9Xh8l0P
oLzZCNeh+627zK5nh7cG0UUqs60LKgzZrojBpOs/1eERC2ADdu3gdhfYsAvfUOsyDNIzdwZU3day
7mIDTjF3Pbip26wKoT7WbSa617hIp0pg8pyC8bIsodOrHAbQWBjJ7phFEDOgsjQRtnljrOHQsh5e
whdJDEFspI76/1lcvtca4ztirpXvKpjrKPeI454FKgS4KH8Re4vPGCn3pOcuP/uHOpbcs1r/Y5jD
3kcQKYWnGePOZfU/1LrZv4FnD0EmG/IN7o5q54h7D2dak+Wv/bQHFXlcDo9TEU5gu7qLBb4VX5NX
R742zr9ZNPnCbInMV99Hno+J2bSzhamg9LqRK+A9LpQhmk57jiVWFD0d75pleqQgs3demrFN/A8z
vvwN7ZuglCCpiVXK9fk5AOO5rvChBDnpju/wDbFMaRfAD19QMmekfzrkWNMoMKCN4hBurBSygbFs
8/UPXx4/U/R4VTCKV5JrgcLAUyzS2+doMFytMOINnf96MBp6EetD+t6i18Z+XPUXRNRyccNIWZDM
euVQYYX84iATOzTLMitKZ2J3g+5dF9emDjYsBkv3nz688maElCv7S1MzZjr3N79EzGGlSEdhJwHB
NyWsjU4MWnseMC8AHra3zal1OCQmoUeMhjBhrk0d7xRBugOTbIGz9ULyWVZ/rsN/9IZWhQXnlkVe
LTtVZwwT0aF4nIdKZvnLa3XEBjDDZ4QzKN/dQbDmWjDVt9zB1yb2eHeuBTb/ErOWLcVG2YeYVOYh
VFiX+o8F/xH7RkjLKszzJ8X5DUxquwfhkGtJIu0AnwUgRVMKVL0y1eoQJ4wHGMApqhiB1D0QsWoM
1L0bF4tHhclpOqkpzkEnYBcGYePtI3baW3T4+DoF/2S+5hXaQPVhw1crHqs9gpJtgYFHw6Fw0TP4
E2dKuirwLP83HvSSjR9K91JmXY1HmcE4Zlh0tUmqimo1kc86b3RXznAPNPIqsqeiyS8hkP0bB+iP
MraSDTLSRNvRu1mS3Y5hwLDZDlrWejtlowY1qhSe9Id633s28zbru8Cd8jrtpPRqRSNYqXdeun4+
FVi2Fa5yqiDlmI77MD2T7yUKa1bY11A4eQb9wj9RGe6vgJ+L3UPKXaRi40tx7ly9zu2+pFNnQsms
M2OdUeRs7x1Cf+JGuN+nyVXmOy7C6G8oBFPC3AXA4KEXZoWQuUETptMrv+6XrNrRTZgV47vrLmLu
TsfLquw5EFjJzEuDljvlJjnwHbWm7KoD1k9lfr+Uh86q0ePpf+fz6shCb9iQCpzgGegwcwKMHySA
jcJDYJyNkdalIx+eAYWU3KYuGXpSmiSQs0HN+rHtJay/s0QLlZIn+BwLqK6KnuTp+ZNWoTaKk14L
H8Q1T9WyfyoWlIFlrK3dckTAoGD6vXqRRYZ9Ctrk/+Qts4OexgYmWrwnZ0/854AwcxiNZU19w6PQ
Utqal0acGExzqDRzbwA39FHuj1k5QL7BvjyO7lA6xwY8BTfr1Ck1MBPc7dSh/sjGRFXL9fLNbY+Q
FXDvDwZhvQFd352mwXPJqPwtZaBlq5yYeo1jK0z3IQNGe7ZoG3QcC8NpTKdK67/KGTj1g8T9ezBx
mu0mj9NdcZuPhSCpi3HP0eYDYG5G2SVwH0kQzKTRr0g4dbeFRIBs8MnAbJPqeUl5NzelDbu+BwrK
bBarl/iHbynCHEZHSnpSc8hWQ3HcJarbmE6lKznffn7sW6joa/6SquFZc/1VRrRxFVI7AlaEAwvs
sR4PiU2YRI/3pStl/FcHevcqoOaFMvoxypoTJOViLVTzP7ZrnZfWnQ8fM1eqEKAbXmmEfUqo22tB
+LnIxXJOyDrtGg8uWA0PXhyHXSe0TybD3nfsCrl6t/e3xOy3T1dIJYrnKhcQZBg6T3xliPZrQ+QV
hPspeQBRDQy+6baPhMmq66gQCxJBd2Nl4Vm1Af9HrXZtwY2GJswYpdZ06oCSjyhmIz/p08FHSCul
QOHMKb+LhAMHDfMZTuzl2sLS2YN1rCElMNupcOQuH7wWIRHW3a1JX6KeGeID5ePUo5xXXv6tC1+r
4GqnJXSVL9SYO0cDDZAiUBL5oBg/vUzAepq5ptTTWpScFpvIvVxO+5uCHUXFmwAJF3P9VB8edgQa
dJc3WBEq0EjsdnET0tj0exhDKHPUc0GFPUWOa89c3RG9NMfLb+RXspfHneMhrfp/U7bJh3eUmqkH
EPwyTXIE18S5gVSe6wEPi1SmOSYbgoCxF9kL4z9484ruTW9yVUaJNrxOMPNaOu8PEnEVyymOMz/J
pWT4PqSzHFU+BrWxWnQlnCh1JaQbPGBfctgohy5UfsPW4ZpABnljMXyUHiXotdtyxXkQJPDhYp3E
mkzcoJZ+6EE07IlGrm9ebn9orUp9vrEOAAK3P+L88tDiQrrWaP8HCwc2p8GBdhkUYmQsMfsobdrW
Mr+gSvtRhkpvaK81HMyEXrGfDtxGIogsmJUmsQl8oTowt8M0KMIzZ5MgZuv157YxYKjahIAd6Wny
QSh6r4x8t00i7gr7rYlrDvY44BorUzRxFgBTsxdz4dmaaZ3qMQzQALof/HbG3o1DkmGztRfcX+dT
/wPCbBVevlCGqfDL+6EnWFJdTeDZW93AwTWF9FY6tcm9x57/JtXdQ80kInUR0HjAwrVxtAD0JeCm
+DG+JbwJzU01PLNOCYQoggK6yqJp+VT+DhbOuWsFcIISH+nYS1U8KuuX944LJ8znLL+MzbCwr1QO
UEqpWLZGREFPkZu362BWrn17wuuoeof120/rKD0LrjW1G6PujNORpgDuZPK06px6Y+vAAsLORapk
0yaVoMsYESIMJe9rKuN947LnecVtzCuQB4ldOv7pSGLwuAZI3Giuc9VQCBwL984k84b4CB6EealI
Yq2KpbnTwSbycPtgAmrWk39aT6vlLo4YhP+GWSpf2veUBs/EOH2U0BSQDirHuklxfIIB96AVz57A
W5ipw23Jd+uHCll+99JwC65Dsg91pnlHLpQcIGYRmNqxfOEhuIklPdiO3qgSHDgAArjjgLIxFzyd
ZPfdBglJII5SBHY9Vsnz4P1dHFfF//TvehUEkXd+n4rafAny0dd2DRan2pDuRkq9NospOw8gGyOI
ZpU0uvsQBaQqsaBnPHyjiuWxqwMdWTwW82drYellyQRInBTHgD39cm7fSm38xw9Ani3wMUlYFDLj
36MlzF0anUGLzIosh0A6l1nv+k7v49KeW/O24DQ3Q3G87PvGaCWvFoXho6eHhLOAihyYV/eYKwEO
88R53V964wvlyjRSsSsOcGg5HDAyjz8geKz6ht375gpKEYNJXs2jK/VdELG/yMnqkvjjmlIECS4F
wOyQr6JOcPlMOup0d0Xha/jBXftQP20bTxhonxv363J+XW3foVZ7wADZqRL6U6/FcxkEb7J4+ib3
VzGT+TVdDlQz5Zp4HVJx4124RYN4UCmYn5PUjXT3Ti7ce5TxSS2MDjRXIaTGltZM/KhMStnSptAA
vq+yqvGvYjyXoJJDQWNQ/pbvU3Ux6Zf42n5x15y6Y//pJz3x3fExd3huNhr0ufK7HzKJJ/2uBnKQ
Q0maYzvwD9C0PNSrtU7D8oenAoXqlVLQCOKbNBLFC1WeFRGwQNiCMu1T1I/YsWKj1ow+/8wNxbnC
RUcgus2acVvVndj+SpwB+V2Mdx5NqSsgskhEeH+68TAMVDwZEBBQ+fdRgVp1UtJ5u//uEskmbHKG
XntRiMFrtHGQjBNgnm4nEPuSqFIi64HrBg9iQ/ImyUAJUDksZ2BLC1RzI5Zsp8b8kuT+5Qq3bp7v
F3CN16+t8YvP7RLalACgOIJ0u5caPT9PNJDju3rex86bWpaV6ggJtarnzSFNtac+4ulVVF2t8d90
R2SiqL2W0bLvEDDQ7ubVDza6l0F5uNjgnK+A1hUjip4PKoZnhaXWgBTudEqPs4o/O41x7/jc/n9f
zNurMZ7QvzwNJioT0nepaj+bryOhQmDR4/+P0YsV6UWduWjCehoqvRJ1oBRZcNeBsl5uNVj8mttf
qIJkMLaQhwOg3lae0+C99fYiTRV18RV6WQWn0vCF4joJ8v3qKDj9mnXjJWBZemfNxDDQfjRirC1c
BzTjw6hIberJ87TNnbs4hhq//mhL2ItgWZcTgPogpyCbOHyXVSPBdvkLKstsPfKIA/SsSHeW8u2A
xi8nnr0prHLLwFdd/cvvqBp4MNWNzRrJ8mDPEFxlXiS0BN+wqWvZRXp9bQK9zRARjDVQhpqsJ3mr
HVV40b2uSJGhTIp8piKWzw7fBf6oHTmGu4JXzPVyjan1P0yWAsk8h1aXw6y08JKihWBBt+d0bUIX
Um2t7f2Y8oIIu+TfrGKpaHH6ksK+w3UUVBxm1C+mqcLtaX6+KGPtYp4g7Fd2+KuE8ZBilt9ygg+Q
24u1QgHE06x7MGuslmwh9dWqt7iFVMicCPcAWCJOrMIIO5v0811xUBGGYozAUlWO3bf+wnTqQNzC
t+x5KM21mKn+uz8Mxa5DYY9YcI6FP9yHB6yQQO6QVU1r5Y8pI0zKNv7/9+7n1zlTLYDPfaKQsvBe
9GoGRBWDE6UehgqkPMtYXLa6k3lVTSzUvYcXbKOumsmy7DcXOxYB3jANx5hJqtLMAHe+mQuYoR1r
jKWgjz/ArqUacwqPb4PSF4pTacyEK53Am/he2m24dAv7lf0xvz1BK6zH8amVE+I1DJ+zEmceqz9N
FLfWl9cabf/Z2aUgIkdzg3tte+Y3RCzYQgnRLpqGCRkFZwOcn9p3QfIGahFqreFmewb+O3hwfv1T
XOt1do45yi1a1t9c/y5s4dUcoPea39XK711uFnWqrsTXNhovBmCup6AW/4K8XYU3zi5jVFJa5kJF
/gCMn3JG2HfRcdVZMpbQUN2iFOKJrxT3ItqZ/9paf39v6rkj87WHD8VnlN/IeGcDCL1eWhlyx4Gg
SsElQVd+ev7iNa0JFvzZvyiaBaDMobgh6y3zxoFqbbNwfAQek9lRByZngP+2FfJm6j3L7kKAjIZB
rESDX8QP/oc+lpnMI/9gpKh1sviUcnHZJP094wrp9aJJ52qqNIvNbggnYnbvEwvUkvH9Se2JoMYI
LPnHhs3lOh3ZuWyRPkZ4GlDrmiJRmPikKPm9RX8c+bH9LmRs5SPQ6OLryo86XyEOis+KJMQvMgw/
25z2Xu6Yuf26DTHghEc1HQcAM5lSbn08/700tUz0Uj3xEzTkD8ypcb9ZwVOY0yXvI5uh1yOf7/2q
aQ+GKJpNX6nYu6aFSWBX8WoMQ5Scm6vN6VR5vq/BAQKsBe5Leh5jZUimsxhk7YHISvxW42x6COb7
pIHd8asAZZeNGKA8VkbCjopRBB19RXEidRybZfyrffZS+jBDfcFomB3Sk6Z3RaN/wZX/oCaXUL4h
uMzz1YS4XEnbCRjIesLdlMqpXqbltTysb+HHjmyQaasHRStFG31iJa6oL5DCVnXAmS0gCp6vGHKa
vVEG1cWRyf4RmrCb6+VkC+B16zxDIdbo/oFgxoSMDDYDE243XeO3GLy/QK0QVeX85GUJT6KLyJc5
hAz2obaHIoimiycwHTMhzERpqQlr5WLudxrxUQb+fXZbJTFA1CXfoeCFSvdJFq52mfnX/mAa4Vof
t9F9PV+2d7clheSQ/cIItedrg24IJbZlH2qxMJ2Nf89NhFs7Wqdqcs2A58bS13dXkAOvh8dQfJMp
S+86gDvOk9+cIxf3vqHZ5J44YokdrRZZxIkDxFZcLF9e8ZDNN3n8QkJc1ELZwt37t24mgp2ssLVh
2jqAeG4frM7H+c9J8FK8k3d6ceLv/cOgkjMGXeE7gyD3j5BjSMAqraIBEculG3f2xYfHKsbWAVdn
pK2h6qnHHjqPZiZu+oOetlCGEsK6LXZxMESluRRilffI7/rRJHkNfzcXPPEKrh99Ej+DVRH01FgK
deMfkykD0SEzTQcLq/69oumNyWPqv+OHHtvsw5pUk/JAOyCERNK8hWNkhlg9FoLu9z4xW92xnzD1
aZ2glmwgcnu66mbZyGO3HikA9MNbmh9oQVn4h5A6qKigatD3KMhA658fI3q0AD2xSae4u6geNx2U
m4PMLHNGFmo96uuYYljea8MUsiCvio3whRf5qXX7GQVBTR8g8IV9Gg9xUNVABSX5bRHD437j0blr
9+Xfwwe4ANT1wM/wpXqjZ/Ur1kUFDDLo8naTHdkpL6FergjrPaTy8cEUgnawS+9ccuhQGsJQo3Wa
u4pNd4x+vqrWrjzT3P8pj2I5pR35fpiTp82YA8OVusvjG1BdA1EJ5xsAUmQ9H1aTHMN92YDhbK/x
MjUsKhSjjmwwD7ZHgh/MBvdvQhV6u/KSddMhYRIIwY0atHf6JpVxqmVEQHYLbVP0i+xHVr4LiH/n
Sz6U3or3YLqNPSKnAHu2DiIh4WLGyJhMwdxrDBpltYOgUPFe3QQMpdB9MHUdc6xckwz2nlTdIG0Z
n83v9aZkH+pkedhgTLRNZa/B0SfZDsTpgx5hsPk9OvPGKbCb1tP3mI2Kxpcsr7u2yrDKjInI9d6I
xlku277ucpnFVdRYHcpsH07p4JdE4tbHuJoNtBqs+jME07Xr2Hg6dqn/57m03SZnqpZEKODhgjeZ
6BDzcmSYC5JeENI5dYnupwti8vLnkRZkkh4yjvNaraajWPQM1AJTZSdSmoq0tSUOP3xdGH3aQIt+
gAQdj0hWjgjOfLwwbsdabBPYiBmoQ//klHG9AEo+vx6wxd6BE0Gx4vvereWaW6xtBOub1H11apJo
sQR24s2ua/wXWanu8K02nlN5m2LRmHTIkkLxpGIp/xLDYuDnxRSFcrco81HmKIEyaxIhWkw7RhIB
ezUGzqedxMpUWmbMEzBMfMtDzV9IcsWCp3j9V6Hg1C5RnqwvcLDejSa6SEQQtiEkzQAAnLGgCQJc
6pjBEm0bQoSjWouNAgG2ZYNLgHKO5rye/Grp8QXc/HhIg9K0/xt/8nVpQCvpRRAHJyyJoGXdImx/
P2vXkwMV5sI24YtYotaQOuiyiON8z/NqqQYQbR5AOIl5zwQ7JSc/Wdnf4HX74Jpvxfx+lp8ZVY4k
XPQWR13WE1K6vC9Q8EzuNEvXky1XZtT8vDJM5AuEm/yb253JA4vG+hud8Sm5myX6XZHE4m8lu/BN
NNSkP5oM9PTudVqySFKrTwZwy+1N5okgslx9yw8RWKS4Sm5oZgZZydcUdn9pDSperDpERoWBRoS8
jcsE6RUTkg3RJr9rOh6lxxsjaqN/SBAnkG6R5Z7wSrOWRileaUBKk2nTPvNoYDoM/VMVTGfwR5K2
+rRM6OEtfQjbBfWu3E63+N+O/knSlF5YWTTONEMvTZ4LWkp/W61DUkas3YS4bufskui2kKMr5kDU
YiDUoV3Pxc2QaT83QGKiZETL10OIzqw7MD4HEQVprjbN9/q5tx9+KqcDlhmtOY9LnKS7aP0T+1ea
d3f4zAZUaXIHVBvAIffFbTCePKqansUqxlsTB2x1oAh6GTQ6HxwRDBWIq3klkLjsX3KDUu9zpJYW
Rmv7u0m8ioGCAt6guREXt+kohWlGw3WTPHcm29eWloCj76VDjgg4L89Y6uCDe/W/OzDgZbRgjSrG
YOiZJHRYWkJtHl6teZnt983J4y5dhwqsg75WBfkjvICwQtIjkh6gFzSbihA1udyEE6uLQDYr/VL7
WFMTM2vUgYXRewwo2EILbsDf4ccLEPtXRQzWlpXInRudNVey2WuvLOjtJzLJKo+egRrSaNEJ1eMp
QKN5M1WErqureW4xsr03Me+x+ur1aEEFFTcJNjfDw5Iuwr8f1W7j24BNL0USAzkue23Pntltgf4C
ka8k3/BjyIKCCnXAhHnWz7W4MGAkUDM9x2QPCU/3Tc0zZmrwyphD/QRoGTWYX9EEg82esrjaV1wC
7nyYtVB29MemYYgC19taniYDta+r7jrfdHoP1XvfFL1FudmcimlPAaEUowt15Tyem17wBfWtOo6Q
8nV+dMW7jQBZa2qQrPqf5lgOv1Yiw/wnFsKs27XauiGmtDgI4VxSbR/rBF801CkUR5xyBtqFV0E5
rcJbvaoePUUl4sq07MzTz5P8Dp95M49Awaf6osEMw+Tl7rVV09aCcBIeVxHsi/LDWSrfUUBUxc35
B9hHsTqlKqc469iV4oC9Po7Vj9/UfeNAk9LXscn5rp3w9QzqwL43GYzG3BJ5mo6I30Stb4L6NGBU
qs2i+fIdcV0Y9M9KerN8Ao67mE0vfhmS1dxypVcDPzl4QLx6NmBXQJK/XhpzTjGakS8w818RrNSB
Zg3mPbR3aGLkKiHMFGxTHVVghaNYHPtNtd/MfvblSTTxZ+3/YAV+LmRvcDKNRRb3dv0d1o7p0OCX
eril2FfWeeYhoDUsNAvKmr8AcTS8txT4N7MB1HOVPr765Y3zsFY+ccXx9DrBQP0WgSdFNJ6PRVpr
kZZIrNL5S2qyAL+iL48Ry3YbSzM5doCd2e780sYXGgt0SbUSYZc5byGgC+axF+B3+zrstV+UUNnI
4pN8ZfPi+zdK/nvChFUL5PVkk7mtsgO5XT3uX2es4QiWgzlpGZkMFQAM8XreNjFugT4CH417w0T0
d9PkmBLbySxgmP0RA6Kmfjj3aN6lBmuqThE/xbt4nuk8TT868CFP7Lpzl6PsH5rGdIYqFbWcV4mF
3UbEMNvRSUObv0yS23IxVXtsj/OuCGh4ILflZHqY5FGiWzqKXQzXbqFdZgXRd2Qh0JsLRF5VcgZS
r7gtL+SjWuNjMKXj1nyzS/rXwb98b3U9bhTa9KAS+gy0lk4EJzKVg/NH9bbJfumRxK/gocSLRNXz
INlh/jTb/cBcTb0bIacLqy5Q+SR5HYzv2Ni0clcrzXejiBVwqyE7hK4NEdZtk2tZ9PJMP/NUpeo0
njNeklskVJZBUu4jksIK7E16k7UCGamg0XyY3kLDZBAHF0/8WF/lhFFCYc87faJKYt2l40uH00NN
g5u54ll3T3GuGdd0V3ouLrSmWZ8y1FU+GadMUqJnXh3iEVQFG+iz/TyaNExH8gregooMUDdfZ1Ob
2gobx8TZAsnfmaoD1fWnPjzZWyShE8nhNsAAMeA1yC3cAgUVAGK+KxqZpKqy9iJHYSonaFENk2Q2
Lwy4LsB+19+8ffFRY0XHhgxr1/fZSfUyiZt1D67oKwJmxZHT3FFzA6S9KWIrFrS2uv2lq+oOSsE0
5vwEN/htHTIlfiaYELvXDW6YQE8WHZZcIfiLosM5VD9ud8gQKJocYWvNVRLnrTy3tnaV5Fz4kELA
bhpmPMRdJfMjMW6jILHNJWpmbRivhHZZ+FSj6hyj24tlKCubQWssCnMEUPKoY6wFaFZ6iXXTE/hZ
r9DcRwWkb2eNPmOCnckLE04/OpycnmQWVYOMjv+DB7cwZukoKLssusmqqgnqz4FnTemDdA2UQU+w
p9AE7C3oorVuF754Wf+gXFU5ptWPs3QZdSA1rCQYQerCRPKNZjSsM+U78hfUTZ0ZPuL0vE2sOLI+
ZP+vX1ms1a/D8ekTZR9NaNW7xIGslUSb1I6G8lSlERPN6C7h5dRVC1q0K0l2wjU1vw7eSlOSYW8q
mPwBaBMNlyvolpp2bFbalCxciTGO1eOITFIx1fb0t7M5KlDCdYbDiU9PGDo6LUzU6C6XppdcKRTN
zstUVv86Dl2SOxsAxNzRoltmUDVfmrhSFrtjjifumc9Shhq00spel7yaL9ISp50X1lGFu/Q9u6jE
mA8UY7EV1OSzybFFVZ37HJvJq50FOHCij4EaNgTNl19MVY+uGTyVG4zhwHp5/5bgnADr3wDGf06x
dfGeGc2+rt+Hy04llSg+KFVDLyRR8y+hiYQwq0nVKnuRG/mbRwHrWf3rQkihB/W22eser85w1n6E
aBDeygs7Q0N+6SYec3nvbxoKgqmGswdNfO45v5sRywFf6XXga1xhJuaV7XiJddJVYLkaTDTQjI/H
sQG9Z2LuWy7pvHlgRDrvhL1x19iSD7qiuIV8+zVIoeiV51vOCOI92s9N8cizQyeuatKovGjWbmNO
dxgE5E9V1yr7Mx5Bypo/DXQebCJGcAgP5QTsvkzfR5xZWecBo7LiIhGh9wTmx7rNaG4FFpvoJ77x
RtpNPDwnS2JDeGABZ5B0gft+YK6ulEqWnQCoKtKsGrZEFIUqBz6iIYbXZQsEKNIFDRdZlMm4j+JS
uNR429nDrZL/D6jwoOcezyC4xKnkCR8TJ8F+ckF+onjlrX8gcQHeOxrSiDYict0WfERAa+Pu4lFX
Z5AbuEGbHU1RuMghw9P7MNaHIk075xyGgSBvLWV20jgINCzJknUtRaV7Ya38yFRwikUK/R/RSSZS
rL8QAK+gC9XOTVCjlBxdhV+T2Z38/cbqLt3dV6QQwMefAIDhJrCzppYP2z6UBX3YbkwjlFuja63q
uE6iE8tOMIz1XEDHBo+MqL94TGCyudABMxX7HwS0MxAplygKWJusZeVzb4CiwaC41JjnNeY1gnOl
zUmIkV+MWkNf88VzELe3ROrDQx/4VPjfTTUICgOnrq54bpKiqIyxUxdIEFT1tmKn52vtCllqUABh
Fhgl9hkIoYSzVxIdE+CsuCQGmjhWp2M6uFJtsgRCmCPsmx+hz1PzuoaCOuH3Oqx2CbrSPJNjuxf2
n0tBIxqJSpVBCCmLZ0r9sx4p5cNNCYNE/jhM+gZgGR8rKdioN9baxkOCYCx879f73+gEJdl8b3A4
+B0E9FHn8QrglIawHHn3xmDjZjx0cErmr6KmJ6QIz7HU5R6JNfIR+Y2sjbtQsAccomvd7JQ5gCQR
pXUC8NXHoODBQahzdP+J8Ku2lBj+VPg6grRnt2eKaLfhh1/ZHNrAoLrWq0bWVNWCwEzYOmpNa42c
0VI+jepC36/K89sX2NO6LFJcVD/kxgxEreiUszBdZmRcPTC/NrfSfNrqSfOcGfQSCH4jvpHsKcso
LqJoDpH90+4gRJTZZOrM03KexG9NHekaagrEE1j5MNqMtJ36ZGVSIulVrjYFH1Nso+iD1yVzoSoM
JPhn/cM8yxPkOxpuqNY+QOx4N9X+4mf19oBug6FesNhNIFBqMY7UiLBRfJcx7TQ+4CNiExfEw+P+
I/o5FMNSRomppn9ZAI1v5EpXvNEQZo2TvU82J7iJrndeXUPuKahw4HUEOiySSwWODMRgvtwRy1cp
4+etCKcQp9Cdb1pV75KgFsiPaf16q+fzxMZHEPc/FCNw3pavnWtFGSajb/dkG4MkKaeAUO8Jh3Fo
icErMn857JTFJ8CcP+IjgFUEHgE+Syj0pgQlwkCtOFdCXWT7W7aF03WTLAgBhyGPZR1hlb9qTnN0
+pu1Sg1+gwXpJsl5nSws9fFvK4hzPt68Fa3qOcTnozr9pYkVyfZse5bmTLgG8Fwz1TLk7FkXOdTb
R2Fhy1Hct/aWMCP4Viqz4Zx2gqABqfoMUPzIhwFb7PeDtHfewX37nzVnO+a2RQ4zznJBxl2y9wXZ
yVRj9zbgvJ0bovV3vnygxUVlyv09TwwZ/28yX2oZkaXD1Dlhicdz6S8fR4ukO5M7aXwc3t2GEuDC
xfS7s5TMBzqn3N/cEr/EA7+r+aoHqbTKPsG1kxDDEsJFxUQwuvresuFxaSTiRe50ubS2HtBib7MO
ZDcsdURc80ju0qR/FoYvo3y4fzcHPK1TzB41sy6G8KDeOavk5lX7n9hVb58iSmU3q6NBMoJNeEus
VVJQ9c962//UgykKaXmopoE9RkF9NEupAz1zdut9QkOhqVblh90Hu0c3XlBq0RqmRg3poMvi1Ink
D8PnU/Vjbg8aj2dTXG0dlhXx7o4L942E+cI8cWAcXVm7cFZ79qboC2Vp6FMiVS8NIPfPveZgoqcl
IP+QAxs2khOQbps4y2Y0hcIOyI7YKVSc8NKWKdsxmyYrBiCTC1kRFiv9Y5FTkWa/Dy8k5tGajwBE
+sv74Oz8zNXROLtB78fem7MImFHgIDRI1r2qg5OMKB+ff03SMjUeYux9QinBEg7FtqCzUBjp0q4p
qA5SwOsiz9cCmtcuLjLPMX8NEEUOtzAwzddzl04XaVfDq/5jtzQBCJG7Wwz5hofxq+Y/OWFSLV+t
YDZXMxjiW28yCHRuM3rcSmQJHGxVn69nbM7QLB/mmXMbB+8e4rgEb1LrMDm9ldSpvKakLAOPVYB2
T2hMw38jeqtADWfFMrp2r2/Waxq8GqlvEyxS0UVMVP8qgHaMsBiN+k5RCoOGE/eDWkHUW2xwk7u3
oMwr3zPNdow0Anubq+tlEeH0MnjgAUDpWAqaOurl9OPmC0fO7UksZizSypRJqOQL/BbyvVwS3NDU
+dFcNZ8R+QhIDqjSPNzDb+6r5EOF4Cl2nHIL1N0TikiEPB0E1+C7sgnQSwMOjtFQKjx1Bsbolahg
lOr3MMACOjffenPmCq60sWyTllbfL2hL0RcJUE4pPIvQ6mrd77fVC8qXQyYipn2dMIb31nH2Fr3e
BpROruNhK5O/gNohf91xE2iyINmwej6V1EbPm1G2SJdP16YKpD4qB9+alVxF/rSGhzOs8ES2OCDb
Qdt3inZvP+Bv487tg5mlA4NSqh0TgwjFvMFb0GuFmghdC6mZmXB8v4SbVSvqrM6JLwy0mKpsId8s
B1jXFU0thq7XEL3nwMmZYs5lYnrFCoutQ1BtgECEyWz+OP7sib7BS931KGwV7jNa9r4VkSHGC19I
qnT1Mt7I7KCs+1zl/8wMFjKFOuqFk8G9gZUOBpfpBfPUX/nb8NohYVCjOsb2EqRTKCOHryUnEqwu
9dZQxcv6Kk7SXNaJSxE0LgnIs3AFKY70lkwhfwAC6U7TEZVzWV/Uy4Pj1JLss21Bmzz9ybgTbppj
MhcvRYXwzjX5+h9VAeQ8FYscFODc6tcs02MF83itle6jURwrnuxkQwVay5KRFYTPLsgkVhwKflGR
QOKPGqXX51gx/RecDrI7gD5yr1hTihHQgyKm9PFneZIOHjIbFkZe0QSvK68u2zRw41YblPW7XJbX
A7AqJrUsA6ZFAlL0sSkr1qiAQGSTLu2soKfSdz/48oweTyq1IlikWfZHaFgJO4FfaKkkp62igf1G
xTHrWv41A2tR+UHG6+v3rxR6i69AhDCWmXc8GAe0J7dsBlED1kG7mIQnCU+BIXE/ecULPRZv9aW4
nkTavCvkZN+PBLtCXZMMTVTEOlji3SHeO6CSLwaTX29PeIBx07rVl4L6Tgs1eQ3HPYm8klU3wWft
ROE7MJLLB5+EnwtoGTz/erQZ9ELSgtBmLM2Y9Gc386m9Nax1d3borD0HerJNB+bkEVBEQFzqXASf
NpGOMCUmmMKYjd9N0g0Id81CaRU2utTDeiOs0XzkFG1bot2TRmuIoQMA5ZLwG4cZuWqJH6XeSJMw
iFAosXux3KfvbqnrW7s+41qaA40vhPtwuxmTA1n04S/xm13rm7G7axckmx1KRPmC5dVtCmVnLoZQ
+7/a6NdBSfsG5qPSbLeZFZzn12yhddji0E3EXrxQuMgIhU75NhgdW0TLDLyvaqqRJHVqgSHlj/30
39i6v/rTwjvGFYi1XyLYByiEsJ96Uy098ddzS2HTDga7P9fgvpA9gSxJwzs27qiL5vd6ZCw4yO1O
Vs8a3vGHrLz51f64rKmT0W5/MTg0RUXabFZ928PMmdPUT0lmEgDma6OFGKjKHMuTSbsyx2QU+4Ro
5i5xQd/YQIvVmOeO+JvGbdyQuWA0X6YEDntJQB2Q4X7dUNcrt45cWwaOpF2RJLaXozd05CJPbf+J
zPF0Od+CAsAJTe3T1i6jcuDijrNZvGrC8OB9ZfOSjnSUbmEuzQ95qeVBHgXSPEIEfCD/73I/q4C0
tZlvguorgO2tSqd9j1owbxBgm00PFGrBdpQ9Xf58mDaLAXeWsT4063AAQNibRIzGNwlqx12mXc6A
+fWsfWiPgdKLL67guFf1ki28cqBJn31DcDn+Z/fsSO7efYN9Ho4lEfotbL8kGku28iYZ/rqSNs01
S5SzForbNrt3QIoPQA7WP+Kokos4z9NwatXowo23kPb2MLK+F5VCzJc519e/mil5UgFz6ZFRZofy
f6v0mDa4tyigMa2zZz3UUEzxNOetZhIl+4YmWHVWcuGhfgUSq2ubiejw2jVeN3q0fF/Wks7PQfYy
F+0B52htRQ+j1cXtBzhtERXSVPWhRjO05X5oyCO1TtFaoUcnN5e/hxEbbZAAegIKZlqVoWBSX2v3
pqVuOgb3+MJaxc8CKU/+JbZwFJOpsoVZR3z99V6VlN7YUzRwa/92apmqJehTdlvTNRcbMRrW1kFO
qpM+D3V4lVPC+I1PrV1sUPq9cCmar2S7frxV9m9ltvjoGEu84IwqwVjOApya9OLDDE+mW1WYL5yc
KDn7NAXxtRIoneKKH294p7HjpKpsn70D+8MLTQoClTE2M6Ip4z8dMfO/8khV3mNDwKsqsS/qof4k
4cuz55LdJk0ZP2yQsbg4RleQXAs9iV1exA+3ICndA9YVnVJbNjpCOHikrGAJm+xg4LMftToSWKKJ
xyUJ91W6/Sjp08xoFxboiskeWXNWfnG50As5Em8NSQe4XPXxu4i6zJ/juhzg17bQXpAefEM5g1IG
uXuGMjfVklDLhFGkPJp2uLbAaHIGiy+ZM5FHXs7qulAqylHOnH/IXsRw1JQFjN5aSeQKT5zPLdIg
xtw+Dxpw26T+5p1BdpC/yWtH6CtO1z+umHWqRyidjUFt+5fLx6r+/olu5sLm30p8uBWV5dZFclGs
Z2/b2+DkV1Oe/elzCc4ZJe7Iq2D3eoTZPgCQ2A3forx5WHAJP5B91ao6Rb+k+8pxPpixGjdbL4/Y
2EZkMmB7qaBDxvb+iODGZI9ZQ3U/0JJHTZLvifLI5CgVcHoGY5u+AZLeiFdG+n/ao+YLDuefygVK
nI3aHKADfNvG26NYSa4Czf55v2YY5YgjVHb5czNLikBCsqpgANWuw0BOW/3RPohb4+tUGIzCWJQu
Qe0mJyEzzbKb2yaOTPs7tQD4+HuAZ87tlKp7ktrrFhfRteH41k0KK0FSjlOIjBAx0NMHNFZefLKq
Q4xhzkTVKTuHbo/ylVQgIxuis+9U7u+hzAk2pXgVJ/+UeLiJgl1wzOOvKFBR0X3ihSLv9K9/W+KQ
GK/kB3H1xvjk0rCHe3hgIvlgiKPsglfCzi3XNt1N0wDJw11VXnQHxHEXgxa7seXzjsUDao6AHIjv
fhUwwF+Gz9gULvrEN+Z3FUMwLIP1BfeLgMQFaT9mwvyFatQ5TyQk3CU7GzkFZxNcGo25/uzgprBM
pjFDojFRVbyMzBLfwwP8ur/8Trer88THakLUYs73NQJwq+RyuK3f0A/czbjAvkAQGKyoHkjoPoY/
cJe6PSHoeOR9RpWGd9Sj+khpIm9h7g3oExSK4NZnZGBMKgt/beC5xoKGjUqaBAeNJk6bCUSTaBbW
U9LCkdrN4FYOPD9UjL0T3ybGW3+xMf4f88CoX9LIr5KwF0MQBLNyK9EOKfYO/VJ93yTzVel50/Yf
iJXR9+5nyPRD+7Uyb1G5R6YFo97U7bQH6/hj2sPRjDyOIWFXMLDa1OGDwf3d7SJnf/8wjyhDZslv
rcySKus15uq2sB9cEttwtPP/wb1dNn4fbTPrlWT+1wM0Ty/UMBMPDLyng2BCwNuCSRB8DSJ/fMh5
P9pcPdTdrG/f5RCWw6fDPS7SmXMQ2jpxRwH9W90Ylsr6fp39XCZm1ziFaPQ8RUZIC4Y0NfThqyQC
ZpQK7IPk4YrnTQAYfu4XdOnt5Iafa/VggHHG5hZyyNBhmoHO0U4oUj+PDJbL5qQc3MMTP23u0Cfx
vekgZGPVh+bwD1qnUOJ5LUFIqcyPs7VeSL77Hrye7ml+8AHnf3TanKi1bqDHuXdQN6Gmn41s4mSE
NUhMlTe0r7pEmaolPOJL1H2IroLPgAPcGs9PnFSq/MhC2020IzlkxR6/gn8aYpUrheI9+qvP6FC1
zj/2rEhPrhPIxN5ddtN5P7mABd5996fE9PtgGSnREvrpMeSRRtgLb1kV0bUe5nIhb3YyZ07zbVLa
3QgPru5Bc6TTqJVhAZ9NP3ya/jWj+upKpn4LtLL3Xcahlc6yekRsiITJ2veCflT3oiAjiAzb9Vg3
UhhSf+6Ay6+LpcFwxjKFpB+A3MIU0zP3wl+cInNzNZEAU1ozjytneleImxr9NMQSgXDOLSPvyXPM
btLXe49jocmpIieDJr7HoTsuiOubBqluf8txTUIdZIzYjD/EYZJ8YKFdBUe1sEeSNHaC60/dK/g5
EWdGFqhbcaNnKifHk7fIcKcQ6mkAEigcNuowg/AoDPpOk+mkysxs/E20fD09krxzvxBEuEXt+XTf
GmK2PNNaeHNJ8PbzvFm+2JpZcoGU4l/ILH+OrpEdDXDKhVxbeUbeQF4mOLOl9Y+hSb4IcO7NTkZi
4Yg2QsuZtvfx5Aj/cKDRdeGciROtIOn495TMqwr7HpjaGJd+yHFdHIfihC0HiWU60iQCd/hx0AXM
0r1Thv66W6xUGxD+BWxPDVhvlfwoyzhPd5bU9AkG/W4vXr/x6XN+qucSTm99U4YsLRm9ZWUypue8
PI+712fvFa06+nNE2Qv1NU2IIIcTfw92gRSG86cU2taTA6X0mgUSUiMIZthsjqy9gAMEKMcGvfh1
YBWRhdvImjtN0HtUVwpW0vwmKV/p+7s92VKiSPIu2QJv56Go9kpApVSi1B0qwRPbd6HnlFXf2tjq
oZERRbFBWFpChWcJ976xRE8rmHH2mqlx0KSQxZjC1fcne4/aSQZgDoOkAQrwJZYlhV1iiy0vfyw5
/JXm92lR+McNBBEz++6XeFf3acAI5lvwdW8l6sMneIcWzKzB372tZexMsQBwo9/GEZzF8DmGK9p2
NqmvqOD1NbRhtMIcVli8sfZTRzduPRz35HAlKsgkD7hnXBV/HKI8VctQFBAyrsLgRY5Q9OFLN/Iu
LJLvtKKQnI5H4ivQ8Lo97SSsgFlpxHvqIFPScPPSOguMeDpN/jtU0aPkpHBfl25+q/vPZjFygTz1
D0U6q/gMxn3RqT0hKLXpSY69y7dl7bOdiO51JgyI5zOX8V/JGzV7x2OE8rJAV2im9drF9ZshYBhf
1zJuOXLg0puUZKdrMucbgJ6CFGNFTWIwxVNsboAasl6ERHWtsQUeMR3U2ERkO7wmwauKzpAUle7v
7hztoGwp+kJIkrjTTox5rYvwwHBv9qrEYIbE4bxB3j+t69h9NuIgEHjisE/0SmcGrGjUiIQbdU9m
+3mYGsSfUxz+eXFWkXNspXmWep5C45hF6qNN4fclmgT5o0H0y+bViECqKdAxfaoBbkhNiKhnx6zh
IQidVVXJneF2KfWHpkzLeKRCFEtkFHML8O57xOYJt/4ZwpQZF5BJgfeQEc8NLXouwlIcfu/UI4m3
2rOmdXsspbRBCRwVwE8s//hMM2VmljGZ5NRRztuz31xldL/BUhbHr37zcTrE/hLWfQ0oZuMSjHKl
Rgi6i8QawgeEI9bkwgfpwuraVesKcQeW7VVg9oJSoUVqY4nVMBlGtAx37fqL0VmPs6+TILG6mDFb
qfzdJQsVD+u+irZ6NFFuauaA/wcvYkr9AchbrioS34JCLwskzApRt1KcxWNGrYLl6J3TpJLpYAKa
Wcrknd8JhTrVwLUgh2jYrelZ1xTP5esYJluMFSjw14kQ8ODIRcyCALVBEB5aswZE0K/FORb5rxL3
qzg/xrE7Q8T5Qrix9eo6eJjSt1SlcQt+NpKVi/4nANTEkwXLrxziKRaPd/Ari5WVVeYjd9ucWVyd
+VElp7qrY1VWuWPuW/Cpy/9Js4NNm2OrcWKUuinu0DZAoAwMRWAosmGmssOf1WeRAP3dfhkdoUOm
aWn2UD8ALhsjPd3LU5BWejbw+cRIEP4fXsHx61TLKWvKWeUaylpgAkaMFCQMctlYklf59pnMWu8V
DwVEZfOftxAXoLlwIVz+wmuctJL5zMAnwr7+s30JYYZb2JNJIjn1x+2EL0QW/9q1VigdCYOFDf+c
h31odsWTiZm1ANG/DstmTbX5FNln9VM5RmxPeH4/5rxlHz+NuIKn47IsQzLVeMbBrBWuw1uebJRU
kmzb3J3jVqIWhvP5WOxkktPo+683kSMAjYFOIMXJ3OCgF63o3xrATbg9hyXora1wBzNn1C7qU4n/
jcJWSg4XSpZC7hquHN9lt9O12e/kVSCHqbPdADG+HbQPwrPLzSyIJQtSQxhtYlthXce/mzp6pe1f
Rq7DLy9ZY2caIdogbO7CRFEXX8ZEB+dg8e025xT+BVCNFhKkXUx7DRvEhmXlt38cHJNRBfhiQuLn
Xi6zqGr+N9n71/ICQU52h0ADMGgrrq19g075Ip98PHPNgj8t2UWIF2rKKacYNtifG6iH8utuQ0jN
yMSAPK7mcTqUKkemy48cPqebFNo8wCmVxVFB7SOYjXiUVscQtO5Ze6mFrJhGKuybQghGVRjhvIib
ofeI7121FJ3nbk5MvhXRBI+99uroo3JmmW9ct26bVMbZJNpafKqjhFml/Wvs8EYH35Me9fCmW/xs
gjX0AF+7zGIet9I1FX8L4g4jbxpv3gfig+Yn67GXCd7ppo6X4S/qS3rcFJnALGUB9nNfw3X5pII5
EP5kfk+G9/R2pmzL2AqiSN5ZrqfNWr0+WgycD3rSCTIJEb1OqWQsPVLrGJ98y9gSrsSnf35+AI1j
/p+uGGUWIpB3v3OsQpgQ5rrrTQ/DTU+WMbkc8FqHMYgir5Gq+7S7oFAsSzNW6yK3U0HyTUYOyoO1
pkCFgJq0nOuK/HjQ0G45raYOoOlGD0+uw3LMR0CO0Zz5KHSjRNAB5xMuvJ4SZZCiPk0dEqww2COg
C3X3ScrGhl4K807xA/icTTKOa8P/gLbsBcJEu8EQpYi4n7PF9i+yac30l1XvOxbf/jWy5VcWSiw5
bhFTXdA7jdxRNVXGnfTVGidKYt8TLgJIE/Ta8YLmEs3RrANHGt/EHEI2HrxX4yR2A2rH4eo7SUXM
kqDH7YB5K6QdCPQibRik0rhk20M+29gj2h7EqN4lZJBmLocg01ToaCPMEVUZBLMgZbPr3yfAxjDC
l8kFrScVHhSfvB6CBa0RCN/bTETH95ni92BBdheyDqv2JpBc6zhFXt7jDpStSbxaTe1h3Te6O/NS
cngylhK2E6fhsur70OnW64ZTFV9ZIXhilenZ4HofmOUwBPD7RZjR/uHEez2MX134M9bxH7hBeaQj
rb3TplNroiHkGd71forq7gApYWSEd/3nyw91H7Zx7oQd+KF64udOy/+4Eq5rMqGi6woSeZj7chqO
cGvdQdHJzsHjlKBHqihFjE2mB3jpJkV882mVbRATKQt2VKVb0gDGxM30IUABwtVBK4MrW3yDRF7D
peA5ng1vSk3Mm8IJhNcy7LfNQ2JtbofGolcSoQUj4dIDYp4J/aCHYvlz4AbHcY5Fxdpu32tF6AMB
j1N/M+Wq5TPfObvgM2f0BsdlR7YKo2qqLuUuKuZIdFN/HUeV7gpNr5NLAgiGTEn6L/YWRCbFWuuD
PufGuGOpIZ/okCsPX+wkvjONZ+nC9g0IbF3pZs8u++YP98kaY+Y9R+x0SsTzoHDQFEgrlLo3DnCM
fMhghdYX/3YJrQuMHz9f0/pmozKjjLX7z4dAFDp0IyFKRz7h4eqGgeWRJ49WJpQuiMZQHzUMjesF
T6zsJ5jQ6EFjVrgBeyPXdIzZU2L2iXwhZW09GFYo0YX1VSmoODxL3s1AtccLPrLMQXoOy4U4cfHk
9c64rckryhLwk0zX3coeX7LYkHheK/glI1wOhjFDuPFwJXgr6dW3tRfHlMBrMecohCbvZML9X0Wd
cJP86NyRxW/jTe+lAZfl8C0KmOcj6O9J5COM82E8EQSWKQW+MhaZrYFJ5XZvm6iq9ZGzjxnuvPwj
7FVBdGjN4reMwIkvd61qVcWScLPUij4yleOu166mLgQDG2KqZwaqXtNAXpcYUik+xBmMhbaPxfxf
WgT+Ju4pg/mJpE8hPBbNAr8vItvklbb6ZAT6ZyhYh/8Jzot1I36M+7nWM5Xb6h7WBZ27UAT4EEt4
e8N9NfD1CsTosiYqh1MZy1oXZdtgJ9TTycZWtUj+gL+XN8cYNBMMmBr7IduRto6S259ZNcHp1jHI
kL/+fibvCSG7ZB/9fo2biru2Pmo26TNjsXRbIV1v6nHOWzVAxxVrVMdrK9TePXwE03dCBZlJUG6M
A5Xga4KVOL6itGAGbstBh1MadkF1FQ+YaTzwULCfw3j2uxpOMxjRQ/f2ensw8Iczw2gb6RROHC30
FqzCh9tiakvWi0fgJXLbAxHGHMy/7ZGucDER5YAmTcyiMXz5qeQsDly1Q0t1Y0F5LYQdM0ICS/yK
5jMH4Awsl9Sjl4gn81eJrrQDzrnQtcxxuLpn/21JFwqWvX3aUaWnjIFs1wDGXeZdsiO7O+x4kZtq
BDtYfSPaXUwU3E3aaSjAOgXZ9JAfh+muQuXR9KGhzoDApSrBvtUQKi8kZvPntBoZKda2MUjunOZM
wb8xtLuT2O/8tnMS2pZV45T9HpeCe//Pyc3o14akREc1WGYAWq3k7fh3v+4NAZNRjJlLhjncMIqP
PWBH+R1ts6QgwsuoMDQzKRvdkUY+jRsXZcXk31H85tNG3cYvyJNTaWqnJ+VgNXiEayuKDPcFlEyb
iXkno41CxB28JkXCzEUBOF9ngWtT0sl+2w6XXmnADTdNhgrl63nnlJDuGmIXGV0MXIRMD+iL9ytr
jPk/IV8q+WUp0D4t2wIcxzXry2TEgrBg8HW/fo3gRHymetuLY1y3HkbXY5i3BBJOvFXJR220x1W0
UMXtbCGD3gmPlt6inneZ2rd33jvY0uUri338rCWrC+cm2ST9t0Y9kI/a+r8cWhOvH7YZfVQpByyy
5p1rtraMtGoe0MT6TSfCYBwSN/vF5OUPXve1gxojmLrYAxivsYQmMQpzq5SihG85Ngo8tOdDzM7n
/Ea22QoRjhWW8GkFZzA2nk+PPB5/QWdtSAxFZPFNlvL788NX3t5GlGyXtN47jLKITB/6i5pPRlMl
Y1uyOiC8kiHk7WMfBEJPotcupv1tWepo7/W64eDBx3rrm1FiL8DiE6nP/crLKMxfoVb1BfRMMUFs
67hYlr4nTv0RLhmVsl+C4NCSGb6Z05tXey4He0FgeOfYJwo9DijaJ5KvgX0v8LhZsqvSc/tCovvT
XBHJHtODG+83jZCy2mkN+SyZdYs3Qv30AdYSrNnmpV168jvSO4i7Uj/bMLDa7oLY5gSwdWv650+4
9IiGL9fKDkaNRq0KGLmFivENW0wXJCS0WtfRMl1LrLlLba7mootKoHOf7faH8C1sw1yW0GhYkg5t
shDKB4JxaN3YgUYnYm2b/ekPDZC4XBiTiIx08FlTmuWTXGa4qzo8k629UoJYtnjrOiMbngfLj6/W
IG2sn1MLoqMW5TQn35Y6rmNSYxH+efsrXPQDS0hgaMRnM8kMn1YpoRv9eZzyc2l6IsnFYs9/tw44
ldYaxUJT6vYRghvEPmhniHj7F5cRPUAws6ZQFc1iYozbNeBab+kotS2Wk8eCWt5qzlwO7KbsVPrB
gBjiYCLiPe1TNtMKad9I5czgBKVMdl86hMlEVfv7LWgUzsL+csb2PA6ZnoBvLT5bG5XkXE5zdOFj
vQzFLLn09fJqKFweFBIBZa362dJcpqMZ4ux5Fnrrhi71aJk4NCxjIiaBKODSf+VtfrDWl9nGd1iu
v/KV3149Ri2dkUTp4dQqPjtP04/Y688jF3SVvQfXXIomnAMNHj42YKXdKM7CdYMwuIvtotTDvmf2
84TcCvIkWVHH3PYHlES7DZuXoWcOpcjzq5zItQuBFWg0GJ/okys3M9RWaJUVfhAZNR8fZ4Cru7YF
e8IGoZEqpZTfQ2JZgYQfH5/zG+xjmdxnEZTAZjo9N3UB7br2Nx3WUmwP01IZpfavMBSYT5dDlzXX
8bWzXlGhx9shnd4yPP7icXGN4kj6dzhA7fn+vBfmWJAId24ujq9GxCSiKA+kNFEXCX94jILdvELK
dG5f9mEA0ccMstk6LjMMIuysJg9Yebh6ghU9b1i76R9B61ozlb5KmmwZ14yibZzvr8+lpJGZam1X
CpRO0KuwgN6/0ZikJTrodVNvRRm9vMHekELWsJhkwHqnRnw9E4JboRuEDBf56G5qUwJrbW7llyMe
8bnwbSAoVXAcnc7soB2VWS3VJjGYsZlQuZqueIKCeMpGhHTZ7q/tHdrUw66mD8qTNG4EB8A4ILTn
5RS5ulX4CEnNVnyxd0zc1eEGWaUI+9ZlEm+LC++ALJJ6dyyZtDb2Q+wCWNVU+/aAwyNVjDMBrwJv
cCk6r7X0EvmeyrFOQ+2C8IIbaHXCIvuPyt6YMKZGSz5x5TrZWFGrJvUIfpVpyCGFhI9Kovw64s19
zrlEqvut/rdf/urrsnvjFJhk31m0tlvIHsm+SYI1bO7G6v/jTmThsDRMUvpSmN0yKvQUSE6mOxZi
J+3pOZ3vjfcif+VYN6E8uzweF//9eOfS+NanbMHpDufXvcTKgxrL7LOwmZfw5yKm1ZQkaS+O1MgC
4A09WzPMQJuTArPeKTw7RxCNFPw39OCtLy3UwflbvxEsGfzussSMLNp+iRElWmh6yUWhkZjFDqNk
GxKVF/bipG+YR4PsH9lFp2pfmf4SbPv9s9f8owLFip0mDBmth/xU/cFAOUAt2IcOXHh8l+iGjMVl
2pIijTttK4lDrS5c41uS+Oa7udPkXg0UOqQkV5FBe88lMo9VyduhDOdji1n/zAF6x5yoJKeyLacM
TobHxOUBwewdE2CaoyT4fj8hK7RE7x4PKPqdwRUwmYBYri6K4VxLAiaXiiR5A76ZQPLjHFOJFjeQ
owReTtbpw+24/UiTfKUVbafwhjj4SEiZFd2I3403bcnxvM4PHBrDTULHEcDjKE3bAo0fEUXp8Yu0
YeOwl7nyVXJCPaoMmOpJS4FsPmhgVN0VC/QtoVm0fU8Uet8oFWdLHduhmSSQhFzySPJ3OnL/fZw9
5L+bvxEOfX/SfJR/m/Eb953bKxgwJvPATAkguC7MpVdXGyZozMk7zq/Cg5/9dQscEUIS5RBmbJ/q
/m9r5a3KSKKuWyk+hxqRByaFRrBgkRboifi6QYb/R+Sdyvarp4Jb6HV2wOR6/cu2AnpqnD0Jf7Cc
e7pXVDyLIXdTZgvCLjXdC3g4N64xFsNkvb14ggPR/++sl+G4qxdf+JQddBwEw8dv7FeeZeB59Qk0
TIAe3hvIvej1RjcDmF1hepprXfEl+5F3JALWgN6+Vx8PkMErYJkPsPu5IhbLUdhSaqkkktx5wHwm
wM6alkcCvfdluc1MBg4Bpm8UOzsHoKur4InngFpstvYfCV33t/jarv8rYXIgt33G+B3z2uXbD0bw
FNibs+QX8VnN2Liaj+2w4dMwpAeCWZorQElECByJmBlNOj6DhaWY6O130VicY6Gf9y/BzKJYsogk
CbqvFmsNxh41DLKjJf3CowsE6AflRZMpqIa9tgc3NYRcdps6Tb4vQyRTKjzlEEolN8UzWfILZjki
V2w42DYYmGukSyYOYeGkTo4ive6F7xiV5PYIzt09ZDuv/MehC0ftK9kD8dwvsKXYV614AeH3PtTQ
LTiiaSWB8qfNLyDcEw8BcCJq/EjkmtXPZaZRTioMfksgqNxxQ5Tjiyu3TFxIuIfxUwrA43rDND6X
aHogp6LfWnPkkb0nk4QZ7SqZBCOZN34EtETm+1aJeRvfL7W71Pu2fJjpaCAO4PB9PSk14BtzAYmw
c+KfAe29x6DMj2fTSTsSGpXT4gRBLBlqTkskG61ZLolkEtwFw7RvmvRDxiU0PkeUIAa2PrbB/6nf
hankaoD/W6UbG1zpaGxMPRJgdW8aqBtHMJEy9pGailQBNXCTol6KuwufCLSTpauz3bO0VS1dpYru
rqUK/s3cKyvX1sc9DQ0yVCqWcX/OQBTlpFd9oz5z96lpwq03rCDy7zp27I3fkJMMgLontw/TwVXy
OMGlsSG8OEzlEEKy81Cwe7kaf687Ng3yMgvACtx+Nihd8g/COTP443erlTaYpnY6nRQ59SrK/hUG
430L7CbPVLALc9En3RFuBSraGG5SxBOORN2Xyk0/GZ8FcX4z66gTzVqRdzgN+nvrr6JcjPAPQz7g
bQyeL9Jc2jLn6e1ev73Qn5m0jpLhstaxKUTGrBtociyLT4d7xHGk/Xn+QO+DTwRFi/h7c6BMaFNb
sD54KKom4JJPitADq66/uvgMWh96XuU0DP/nthqDcVkQAdnIgqaSCIPhaKSy62MPEqI3/teNkFj3
pmsEZV1reNroDGAAZgd8V7betGxbEDm89YT1aWfQU1OHfWbzAgKW0bFt/5QPlQu5OdnwqMOHIsWv
Ni4ooZKec7woiLBZP/EAx6ejYBkOl6+S3P1GhZfuUDl5Krv67rQUD+P0736fj9Esw5hK65Q0Pim6
IbV19KT7fkZohD02LB6xyfu6H9uT0XHFskmc1mP47dvvx0qhGNzLp3v8YAQdj+GrdFqbIzDkGiXf
5b+KHaiPlop+Y6GsOo/3KCU4gmWVofQXcqmv0bjTAOEyqlX/TIz0qwogNXFNm2RDrCJFNmpo1HtZ
qm92dkZBzazSBs7n4VUeZFpR3YB9mmAMMDcbXlv1gmsPzapbzvo5zf0xaOM3tNTE3I5LPn7SR9lT
ScJh2joxKzR7y7yHskvlplvQ0kmrJFUagqA3/IZVzCZg8W12zbOIPEAgiUOcQvPfqbNMUNBxP3Ax
3dYGMnks7UDJl5IXYAZ5rbhY1xO8jf3qO5El2vRbjAl9I8wL+ESC/92T+GwDodMeKmmnGslf5/xS
dBcygQFrVMuweT99JKdea9uaFiyDKX7yVLZdgps9052s3VqnDTVxTL+9v6J+f7RVjGwKs9YfOpRC
878aGLcNC97o1bnp+oMwlK8h0dS1RkeItWXJGi+gjzT9KiYYO3HLr1De8jqqq7Nn3KpXfY4J0Gi8
j8kNqjyviiqMW7CGLQEtHMuzZ1FbqTT1r6MRERAo/8bIheEGheb875gP6fnT44DR9o09/feghAl5
nLRK/ihXA8LriO0b7ijRqSJZiwrvBQV6/mgL86YGNMlM6TcwxzD0vM1nG+gzEhDNPmtfu2T4maJM
D6u81fprqT0Kpfbwni+ebWvLRoeRMVC+yqzJfKdrF+XqFasgl7FvV1kXhj0aQWQ3tKUWaUGMzFkN
O6+s2BK39tYvUJjh6/nc4ZuNyqRQgFuJ/ZrujPy9uuJtFGkZt/M3ZqgEk+hkUSPJu6Iiq2bFxRh/
epVqOOxR3PTUpcOjKSyAxHQAcRi00z+sT5Tm+FrXuN6rnxv8v4y2l0ZoxnVH+g6/ilYp7sYfCWx2
aub80rc+qkU7npIybsQxkdlERTaiu3E3SNSCGUgNbXCJ9dUjcSshHbWdcRUmEemeiPk5Q/BVv7Ne
Wm5/zDjC85AiXPbXnQXiYPBfhzcNP7p/IHdlXFz3cYeLlksHKObQ8VUSqT3GYakdSlKn7FUmxm1T
W2cak3tUWceRcj24IrBvorT/T+NrntdSvaPeutxu2ZWwkDlsri9NuOVjdc6+e1+Eztj2p6OGohVq
ATamHsBWG9xmtISfHtxztFww9CjSQAp6N8Rb50BKTCtisIY8OgVGsUeJ1jH9Vl41Yr7POInuRZtw
wZdKOCh5+d5NLk840fy3jEFZ2YuG3TpfM9tNHB8h3Ft/Io67H1AoJJ2/KZc+/NeoqgCRYXWhUIgl
OrFKc0CVjgyLHvJbUTI5n6eAdUSV7bl072WOVg0BSpcdG/tGbqVlhUNBHR1t2hn54ekTwgVdML8I
0jafyvaQ6abJ8PGel6TknUqD2zD4NvMoM/JnGfjpWHkrTzlnBh5BzHWWi/QtmYSsct9sIvzB69ig
5/gd6BPz+AALGNkvqgyMsR2p6PykBU88+hJSbFcVtjb6W2TUpG3u6JjIx+6sWKXB3uqKoMYQNK/b
h07X0atLsbLuCDpKSsl2DscjpsDUuiJcXvS4/Vv3Bw7ysNBZXfuRYGsKElX37Izv5ODJEknsg4lE
qrL3i8qXmuRknkzrE2z2Xy7sYMjnS3kWdgXy2K1jR6mfAFuWV/+VBByrfjZ06xcL4I7+Og+Ur9Tm
1GNpzCB+iNcNet5IpJ9Iavc69ycn0WzxjQFqjiwkKgYC7CsLKAE3zO1Jf5BDUUe0L490y+vBhW4u
2ot4hsIEFOwbJMRbEBiAYc5qf7xIk/el5Sh4ZrOymitafNE0zUO4Bb3Xr8aJ+idWH2R7bzBGQw0N
6T1E+fZSRk2sUxS3n+jOiHWgitqbOCEjOHXRdDouvPLrrxP7GMl2rxTVstmdonrDpr8ZecXrZhec
n0c5uSpuE2f5sKqs6aOy+DRRwUhmvbgNx8CWRtoKiddDVealZzd/vfVFqp+noFnQ37bhNEZo4020
2wXccEeX2th9A/eLLaMVwL3XxN2dtok5u6vxZk2QZyMjDFGG3opfx+QdzYKMohZNCXf3n3p4HkKP
stDVJdjW710HBgAS0Q9WPxNie9rDe0Ze7AwS5zI2IJih9wT43m7UcrSq+Psvbm+jQNdWzP7f8067
JZxi6Ams5tJCK/sM6tjZo6DBUSIPiZY/oVSLNi6e9dL4QAYnf+GNYm//EOc/KEDoQb9IMplKkx/M
dXp6s6QzbZYxvDzqA8437KisBXfPkGfmkOSNqJHwh8CPqn+xCPPrVGJ9eUPMfeT+4Al+9y/VLuTy
4EjZVkNUfzqKLAPTamV7eTt0mHO1pU074g40ibQLbHk2Yip7vLgES+4/vLTiTvJldi9raEu7SCOO
JZFrBkYFnNxgAe8GlNhc928MPqAOhafNpL7tJ5W0GM2ymtgc/MuLnfIh1jm6hjvJYVVrd8lUsNju
6rGdEHDX+S38BJb0XqlRD9DTIPBG4WzoAlTJcOkXWoCXK4f+Jb6r0d3eDiGh+1t5RmLUvEtT+9TR
B4kbUImD5jAIkTVN2UW7Nl3+Iqae8NFeXrLjDRcGSNd2yRS/cSWa8QsLrgYVr2mbBoaKs4DPFRu9
zmefizxaDJo5n+CfVUGO0jktrJs9uLTmuU6Wi4HpoClUEy1flcgmnjBdmiIdM3F7cMuBVeFLIvf/
9TPLOeOAEdwXI1AKGpxCNKzxVm3V8+9QetFJ+dSdAeXmuS5DpX6X9q7XgWPabmhuOq8UFm1GOyVZ
lunY6oY09qJeBdn2msMhX4U4+o0VGmITWbPGNLHsnjW4n6oMWrGM3eVrbFFWjoLqMH00ZgKocy4Z
U6Ah6q8eqClUQerWZ7PRJmpFjw0JhyC3irSdLClMSii0HU69I+BYx+gzpfgmB/iS3Sirr6tLuQ8i
aRXnV/7ddN1rqqFAXWIR4ehTR3nILVgMhKNx80C00Pl4LzbVa661HL0uSB0rRvwlNVYn0/7BEW9j
9Z//UMtExv/KtNkA8Fozp736UumIsja1QQqdT3yS48YcHc2t0mdOJGmtmJvEkUREKFN2aydZzUwh
ZUsmVBoVWQw+UBOiQCDtnWyVPXB2D7Lr/rPxyqCZw64Gv2c/z1oqp7WjrGGeXl62Xandc7t7sXJd
TuCDFX3K2X8GUW9JHWFez0DMNMa4gIEzaN7b6Vy9vnMWu7aIDUBsq1ri8If9rkGhiN2C6AMcnO1l
trTEoQLVBZ7Q97nA2Urd/JOUmmf/XwURFtDZAfwhZJeBpqHWwXmBMXUJnZip8D09Y6glSUvWSruQ
h/295RwdmJb7TwH1G/DeAtY/6phs5rEtQD2nUE+NoWa409pkXAQa5Pw78RCklrP68e04ZWAFBNZH
vNSpGH++XN5Ceyo5metQkSNQUBkzSrJ0HmHQL/3F/Brp2gQVr+B2HI+1Jq3yebUMGK/MsSfZobJA
EgnCThfwgSwaarwj45yd7SD3V7EFjkUTuRVLReSPD10jLKKcokKo5XVOWbKewArfUm9Vfo5B50AB
vQq2t406aXS2Rmcup5JiIXy+JjLxx6aCcyxs86ety5yQHSNjcFk5aWpDsjtXYba/q9ulhXRT5YdF
BaJUAiW+yLBXv4nrZzTmL+bsPTEdzYrOI/IFX//wrxiemeCnf0wu5fIomgjsmhqNuhxj18T4NPcq
F6ugiESfDOPWYMO3p3QUxLHcktoa0KJeH4G86JmieVXHiAc4/p8s6hIddYO7vmZRT83L6EF9YStU
ur+BodeYqeiP78Zi49C1c6DobivTWmwWhklp6mr3wtaUF0yP1p0AvwkrxtGEDJC+xvByqX7FbFPB
A1Qf5Hr7VlTeYM7IkKxvKRhc9z3evo41EzV76oqJGCDDR5Gel1hS/IkQ+EHU6x1n7T01KhPpZ/bU
lwAuKpMJMI5oDSU7mawpyAz+riRDh7SnQHzOozbFWXMDwL9u42dmyOVgw70+j5y6aw6anCgOhINL
SI0jizcIoNVFmwW5qZ+u7NVI7b/gPNQnakyswP+GHhMMXiQyM020vkitp7CFeGm76evZl7NX31pa
4IQ6yFzubZxM8Qc0LacFCHSpsrnLFrf78hsKdJ5OAQvC8v55NufOItIYBqMnbFwcopCfMqR4EJvG
LH93B0shCHFZxIXnmSs5L5H/M1C4BR0iKl/Sb+d8ws13rqGp0b5pJnuwofriMFYNfdj63ojvZMs1
Go+/In40lhbGcZyYCGmrKqwmb4qjP7mfV9zoq1q/XlhSh3LQUl4UlsvTmjWR8elkYu2Vi/f+7ieh
qlgXHfroiN7xVAPKhK+aLcTt9ZFzCAO5OL3Havd8LrODVTVA7bxyjUMexV+gOWjidkhGC5H/o8nI
PwsW90vjgUSfJpFX5iKLrfyx40bx7IlMXPYrApBtWuoqnOJhbiRYZYC3LFd82S8dCKUVd6l6Ss6G
m/APvk48eHd945wZTfJRMLbANALc2amLAftWvt20+w2IfntXjzuob9MQ1pcYc2wrnebjQ4zVxJLm
IG3nVx7d0DY51My/EKAIKEhBIhuy3Aun+uBuoHaiLYox9rp7jLPw32siQ4EcH0hndTysBHPGv0lO
Hago8VrGlx8hVJskZa1DxsfSnBGtfHCe3owjubCcZhT4pmIcqMcZPjhMgVs6nRWbGgmzCnFUgYtK
M+IGuHxHhnkmpaVneumU8Kbea2wn41lDzl14My7fh+BcRUsvqwtlqYSJMr+2zSFdPGTTLjHQ9L4h
kB38BTDK9qJAdVxehXv1DVt8pKVnCzWrmkSE7QEr/u2EQMqccTH8zoUf9UbjZHa/JqRlC/QOoN4f
6tMpzG+v0bYaKcVfdcB/9zepyhOKeAFvci5vwmWJPH/Qsk9NRs8O9mi0zu9xSaJ97s6dXd+luI4R
1o2Q8zVJQYfS2LOnCGgNdlhGzbujmkTDG2gRO7IrCixWXiwXThnVH8gokBCEonFpBZMHDQ+PeZ4a
oXxrPBZij9lrSrtRcnc9YSPWOHsDmmnLLKfAjWoSOXxg1IetJWcpkF9afJFeECyQ0jR9g34BGRhG
6GNR4fdRfIOEHTDzfB/ny8aIol9iFNWVDZw4H3ZjSNtxkPhj4pDay0bJptgoon5tOfYMUqmli3gp
3GquQfmgnJWwsQoHObHP04SuKL8SZdkBpnzrcl0WmqPTV3jgjVC3dYJxp2VRxmklfJRJ+LqMiiHE
olmsFUCa+ldiKqNT/cWZGa/Tb3QljqDCSDpisTgdXgge+il2g/NXlEP04C6T6nhrOGehMC1IdRnL
a4WUpSc4DvLxTVsLiy5mZFz3FrzGCuwAPjZZpipdcFhGiF3mIVsApKlH0jVTbj/dxFxSO/em4I6J
l0VfR0Vdt6dZ0Ci7qTJqDqMyMmqY8q7/IJOgFIjO6dZxAo+n/9qzA9hnV7RFdj3mJ2tIFTASmvts
8cV2zHrh0YgSm/23HotU3IHNMXTYyBs70YWaNrJ/NiqLhv5CJWJuHu6J3owGBBrZZss6PsFxTLqs
nVvLrWT52bnwDadm675aBctcRBEALNwCMLBkTVoNaEf1NbDGr2lQKVBzimB8o2oTDh+3FbERgyS2
uiGAeuW8llfs9ZBWSnaIojL80/qvFwfjX6J9SV0ipkFqlVfIL5oilCKpgrIPBoILt3csV1RLlfg5
ELfElvO6isQo0mUDKzDh0puVgwn9ZcgZ4xf8Sm9rPdrW34EzGrx4FrkwXHwGWkDheuCmM3YfEBhF
e7ZVv7l8cA6SrBMO1EZkB9C4FqB8ALL8pqjWGVMaC3f/+T0AvDuu8zYCuabhsw9f452JdpoyRiyi
VZjuKO9lVW7oax/9lDOGT/ryktQDiQ/Vcp6V8ySaN5XMpP+uy6z4bLiJ9aHoHQbxty+vWGTeMBOv
pE64TBbM2o2v0N2ni5g5EqKHBbFHcVJtHqsGjwFpytQ5qFrzC3faQJqoHM1qSsj2H2frq0ixaKiw
pijP78Dtmu97xU9OyQ4yBmFnKGkkOW9d+hE3DdkQFqj0Ugkp+yErWPOgpyNX+O6Hxu+g0dKXaGNC
BbW1oqeBhhh5ZGyiRUK5+e5zoUJygFVdiblf//RV2dPfzzxYriY7FsNj6gXx7lf3YTGldKEaqOeH
vf7wPJsQP4YVzQRSC4XQ73hW7oMv7pd6czVVkVA8JHVRph1+r2xvnu8E38t7rYllNsdzsRHolp+3
K9anG76bvykd/r3jAgYIQhwngzscewu103Kl/tD+UAVEgJjT27agjIkSutph6RxeSVwFOWSba0PN
kj5/VQtuLThY9rq7PEtZHVWwMqK7z2hSljTYgygkkhNoc3kESIGdcKgRTmvf+izaFWgkghSM2sVF
oF3SFiToeW9FyzdWUyrCAZq2oSOj9w9XbZJxB3SiGmNrxGqdfMlHR+3eNMTuN22ARjpZg/WdNC2r
Tq8czp62SQStgroRFdEb/T0eZsifee35FqOd+BQ/UqvuN0ekhslQ2gqrzLtMcYDQd5Ay3vNwi4Im
1LaXZbvEG45HvKxY3kjSnzRSbPhoYCgYAa8wOX4q3JWb93pDlVVcX0EzBsG5RY3AMEgWH9vXXbhR
0ul/QfSRFjbgUSzmTlVQEnMYjpmKQMT8qZTmEQQNInLxxbmqD065qowmNo9H60/cOJGLkM4k7sWW
rsuRqmi003zwyGWuBeizJHVcYCER09AXdAHB2jTtN2vmHEOYQ4ujfkSD8xigdUD6bTYpZ8340ztB
rGSdk5RsYsXvywNN8x/5CXTQfLyESOYLHDxxc3CZMIAUVs/JAyE1mzdrRO/7csDlDdL6yjiYVMUD
sPsF73c6TgAeLMJ3XW3W1P20tAkw1jeGi7sB8Ng7q4LMsjrYZHyqtu0PXiK2mcvZbLotsEaZxOsJ
DxaO32I+11G64O9gnmxCOJkO1X3br4ySX/2PqT/iGZiL+ncU+VKtn9j/eC+E8ZYyDqqtqWcI6Me4
v3BUfZSEBRYqoHTMUIrql2rk6GAR6rZ1f09FQzg8yegv+o3hdj1Ne/xiLfhKHXl/H0VhiPkYQGVH
T/eAy/9WmQphQnON22JN0E/gn7weTk0h/owKJ8sh73fZECaiN0UA2cIhYdU5E4V3mXYjygeBaa8y
Y+LIl6+A/wKQawu3E/sv0JozMIvg88m9ehUxPniZq0Dpw+tRNJisbBQl7YPPwB92kD4UCcb+rz/0
IYyjAlxIRzk7mCtN771t1xSpuhXj0nRbF66+7niHQqpoPgMtHFzccdXInUOBvYCOy1qLdLc0NUJ2
J02tut4jOCblI2mGFvF3nrhDB5ih08FyQGjHQuCed4Znv/YsOGLEaFc/FPFFCek2g83VHr9nahH+
d9FFNNwxovpEi/BwSGXzHdlQnwHzu4oEhZ+rbWcsJdfFezRyimph0U6jg9NANCqVfA4RYw21meCn
FyK+VBp8rYce4n93PW0h3IzqRTesl9tMKGYYHErDxbONP3stmovS86gFhrpKd6gUlvNmaAYiocvJ
/tBYL5ijwQgOKl62yLRPAlaXQHZVdgtoI/7oQHLli/f+ZpLJ9HCmf4RePN8sJ7t4TDtN5tkBP91E
WB9EXoFE1yW0Z9b0AVq6/wIFuL6EiK2qsxXiz33pwDdQz6Zo5doH4rLsEwX0pqSldnBJOr+OFsfk
kR3tg76Il9VyaO/kGFR8wt4Yj2CP0kTnfDaogr5kqD8YLqjI5Q5ch8EqrcTfrNzDHdVuDlov4dMv
FJbfTHoddWgHNuzpyQrneBmVlCfBlKJCerl7YrZIedNj1UFXrqyBqsLrN3gKwyv1az6JnOgRcFo5
mwfxfHkgraWas56iukk7ebeJIe6tZRu0xaA5tLQE81dRBdtRm+HgBBuzsfkVfZVymZDNuQlH18Ju
WtCWC2aKCaeBqCMaz1dcgvOXAs/8REg6J+RHRVdps0at8hRiVSBUJfXn2Ot8NDvXukuujXAq7vIC
4yXgUjsFiimH+G32Zk2ZnCH1aPyRds1tv1hkq2CqID2aS6HaMJ5zK397YOOEebuEUel9rc/bS5MN
Yn2q5kdQaDO70QzPZ3uv39DHhpDBwICsdsaKsb7S8swBCSe9/mSpkL4ZIHS79vDzZyUSSBhK4SPu
ikgEqCkjaf1szcWnnMksy56/r3FNaTFlfDRcJJRqhT34Z9y8tMogPUQfn3+T7FmnLtG2e2WJM9Os
QH5OhGZ+j9Anrmn7uRs6UdLylzPUEPhvJT0rpB51IETqFD1eJEUMtTGyqvDNEOjaWWUHCvp4DCbr
kKE6OD3xvD0cfeOzZNCVaXidFvoThARP2AI3IdDFPdBI8uNcSOVMSEifIiVYxyWWplspgWimtdPq
EcIHZ95ZRxWjJuWOmoJsXGQO/XClEudCStS6PjMrLqc7nuaKQDGoiNUCeZSYUKdpVJ3WvZ6iXWWe
yhOg08Mk6CqPBzbtxm37Wjo8Mk3tn8AuAKdrJNBE1/iGWYmjiHhIRp4LOBWeagybbUDg+VUQM4YM
9GW2bTXg4MpO/OCo7ymLUv/G8Ypjdz1Q7YXRZ6qU6DXBXB8t/Mk82hl94qzoVKU7uD6uDTdMiSNT
hkqK2U8hZS9EPPFnhST+aR4m7y6u1JjMAg5CEpnV73yEfv/PvTSjTzeE93lmds4ijGZy4PfhvDsp
xW7l+ZHD9S/PmOPUfOOZGTdm/SjgzLqk+zygMnPTTaujD1emQLqozmsv8mzBeFvjRwYwozIepj+u
egvNSx23InSdyFA2ZB98DijrzWTcUpnqadEp36brqyJcmCnJ9qWRZOU71uCfwTpFurilcu3eG/un
OX6VEPBitseb9yPtoGU3KynpvcIfsbpg8hXVsNh4q44hs+8W0ILWv3sXkz+6YZIqwnO80b2vd7+9
BiO7V77SHp15+WFnrR1V6KlMTKdl2pZ7gp8OFNa+WaYc6kKgEMBMtrHmVq2D2tZhWeSp+1EUhmSE
lymm0bAWw5+2AdYgqV4v5Tlx6FKY2w6z2NlK/q2YctK/uIa89PdhYFSRP5VdnWUP4cTeRfKt/6Yf
+vW+4znZSQfgPPwhfWCQ5G/M7GBtcNqNrU+hZLjdRrW0eOM49HEfetu3LjlCakpTznBenmhBCnSJ
yunRd/pe0qWTfwjmIUkYgT1oCWF8bF6PxeWZBziQHw+NwTkIhl464xiN+lt7tc/8PoUBROOdfKTc
D0kWkS9B6jDd3dJE0qVN2aNgsXJnQ8kp9nhf9DFonaF2mg1GtAuhx2r28kX3jq/adXcwg8Ann+Tx
ZsIKptX6FTjR56nl79WRk9y8fVKYRkiwX3kdFFHe9yCKjviFDHRFrulOm4aZ5pWQcbn65P0hrm15
+iKeTOhH9ygh4z82nwHVnFcHoWrKI5gajHU+tqHPZrftI7XGAlix7l05kB0+aHMGCwI35efIwt9n
zxSH61Zz9X59mw8pE8rtWq7eOeASk0w+QpneqUKieLI9NWFTjDU5+000z0zd1RfkG8eLPwxyPwVI
nZxAgj6DbkFvkyehwIP6ER0M8rsm0Q9sRaQoXI8woHlaqZ+QEfutjjfgxXprJoUwOdZjzhvWAKbG
QSl6opjolOZJllTKIryR9XPD/0BOYktHQ0Y3/yRU9AlVBMVaHPWXMMukhH8k8wGB5qFJ7Vd5x4F+
h34fQRWAEU7iu3cRxdvMxF4N9n915ZGwFmSxFVd318woXYigxJ5Dbo54Y/7ENDbGuarjvAFJm7Wa
Oxa2JtiFIWiYRrhhqaRrFUm9Gosro72npaEf+9DWzJp9yoRFTlBjyxNjXkczpnJ5mx2ylts9v3w7
RBvxH8xf80OOC9CdnHKGG4jkod84PnO5MQ2VMkpEuM2tjPfGo/VQtrE/CcG5//QXECeHs+UBlFrr
l02mml9vyF1+AMtzo+gt31RwMNnq/8VpsUMEff1zgMHs8oyTfF/uNL1j/sYmsEngp7k/ZOAMM84u
hpNFXiK6P5UswQtY9sdYNiky5NoqvgKNdRXH8YV/aimJuhsKrJiMPDSPlMnsKWMklgl3TS3X0gIr
p9F0wLp/4yFhBc+Tw7uVePQvL/uBdMTY4cWX4t245ZAXyWgfNLbDFp3cGr+NH6rDCjMkUCdQ6PHt
Hj6LzpswOI9CqMKSJDccz6gPMkbYUm/1JG+Y3vDDH1ti7V3RGTUuBl0iOKp85Kmt1pZ0Mz2ntUJc
IwJtMcML/MThh2/MxAwZmOZqWPaS4e46s5b6UXbFvJtuL2DMQ5SHtIatPyPwnG3bBT/a0AUYY+V7
tKGkib+9JZBgsz7HJv7L0VAcEDAgA28l+pGfzsrkzEhiQcehqiMt+r1ZZAS1WzkNTv6J6KrrkRq6
EyeMmpYa/qsBspnh6lJQaAS3jp5t5UeazYGKYAEkuYbmZDLQaCU95tFUwDFLSHQteRcr3flhVAFQ
m/Uvh94IB9zMkzEfcFCSNSYJCD/sYwnnmgVIfwxpxONne0boLKurTErZvZOSPaZ7Ndk1gtfqmDoY
xuOvkRo5ZZS7h7h7jlYwI8hPxNW7+3SMqpZXo40taY96QWM48SMcNVY+4mRxVeADy3tK8Dr4J3Nj
IHhUEISE8QBcrEG00bTXb7g6KaO2oyWu+OAukGoZpP/fcsu5H8BxrfcQ+YgbfhyhMEBCZdBGn6Q0
6B80K2vI+6Qreu9EWKssQPGYCXAhVHUsYmv5kGXQ5pJ0EBC44FJj+Hyx7z5e1cyiibKrZCO8d2EV
Q9uF5aXXvXPxDxcOIjawXI5dYmH9XM7QWiLTLey4iIjnff0pdYGF/oiw/kVbxdlRW/xgW5QSf8uM
wo/8JU1+K74StKr2NIThR147nauUEEVn5Fovnl2KaSukfpfs/VYP5pUumJBfO0tkNh0DR34g/RmW
/c1iW+qnVm9OCGzQBf+82mFA9zFJaumQRjrtmV41gZCOa7ieGiUo1LiIZc6DoB+5hGu1zZcRKGML
hQDXH34NREqgxXoXC5yWSpriALjy2zgrts5wbmUjxw4ZRcdrvmK0fBLi+UYcPI8fJ9/h3ElIic5D
0VQoi0CvNF7j14RAdPZs4cwWh1p73ufAXkPbuQ+Jo7vpUiQmsaEGfaxBcolzfs0EOIPjIYRgUSoq
jLm2Y+DoP/flFNHAPkdWk4Bc/fPOHQTVzHCObBU8HnRLb9I0Js3Bjmlmg2N0k1AI7h7VsA/5hhMk
chV72Qu1RvvCAktdXzqLWw==
`protect end_protected
