`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R3v1gh7ror2cqCntjf8DZw/J709OYPyINsVCBl5HTTJnFQg08f6z2TMImi9zQHRN6E1c/u1qiQsjmKxG6zOPpA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MlPLW8UKMPwZtIzBHtLuPwMGL9CgAK1MRvO2r61WEV+KZhmGQmHpJlha8Zfu5RJp0k2FNi8XZ07GOxizZJQ2Q0Gg0mzhN/fv4dpPXJd+PDpRyBMdczQEeudMGehzsleV4rs57HeFv+Yix8SqJZppOjIHwu5r1c5r8F5czvccx/k=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ziik6buE9TJQ8xqqW/aAXzEBttT5AbaCBtbJbSMcr/G7LbJnimNRxtSOXWxrO7+cXYWhkpfzC3b218HlBabiYmBEyVfEie0ynlatL1GuvbZfDPwek7zHi2Be2LxWAHgS2yWeQMfINXeoWUfNDc9rLyag35O3YWhtoJ7rD3pxEWvAZH/UWgbBz2HYAX4yfjCWPG0/VSYfNR2jphi7YWyGIBxCMP7ccXTKYIySdRPgu5YDK2hFWkSFfMLYGoVmvbcQfr1/ax3ZnWumXHxVY08cERJ4i8V0nFFshgFyLYl8DQRjCUNsOHx5/iuSZVYVBG/3rbvYqLOpWVKUydbOXAWhEg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nCANAO7nuypyOhPQ3i6tirWPHk6ix7eUPGnoLrquGGLJw4m6f6jQABaHGsEQfjVZbcKQ3fhDB5rHKnjgnXoxhlj3we3YFkPTAWRHdF1sGA01Gs8kZA+D0PIyOwVKngS28ksQrnhW+OYnMxQHwP3wblwls7HRIsnwwi04o2Lh00Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qvbYmVg2NL3za0eI1wVfMP5Anvwmtdmi/G9lLQaadlRdYfvqIyvpnCn3kseyEe9m6MSoOvn+JAiG3eRqz5JfqEo6yok5/YsQWJqJgAPobfo3GcX6bx9m5cYuhiWed7yxrt5SiDGPA+mSMVSkIS/KSDwfCbuYhR/PLMpMcwu1Qy0osw00ZGi9TgjsPFl0Tolr6LYw/+M5rUDwYGRDp1/MntUEiqMD4HBP4L1vDf5Ll4Ayjmv10Fcj9LbN8Zw+C3pbOts/n9Rt0LQO7uumtLu5CBB1WnmxBSfs2HMiW9pnmIaSIQnI/WbWKyo97kW1FAxxq1yMn5thE8l1X77N5lTKjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4295)
`protect data_block
enmSH9SRchrCZWpvjwGEzbzEsoPZmk1P3EfnzGrxB+ijBm6RNSuy5vrpKDh/2y3PTXimt5Ibk2QX
glqeg4oIPsaV9n3NHsw84S77B6drlam/VTcT5dDmGERoo8AHDR+NAIVY1+aeWjQNFB/W5f2su6fD
MFnfuuhW3AZcfHfJSINGkjbfb1lBOC18XYuTjBPcGEKj14HZNFTrFYVlqXqhLPQNUm6QUL+qpOXJ
5Z4nBcE8Hpf0shwAzqBXgNvMPXd+yMz5+spzymX3idzjTtagMH0eg0uBCM+Ef+Qnml5A2xZRl8Z7
X99E+VB06XgQKyFRQdYGftXMMnFB1yCZabAXNP/OoILcl7xDvu41Te+ATB0sIsp2xwkMLtzBm5Zf
FtT4wsFK/9TlrqwgExOHRe6rkjJWhvR7IeUfnc1cJNoN1ieY5slmcL2akvuAcizeoJp+nDlTNrdd
NRRK1+tmM+mV2IG343Uq68KLM7lahFJ9v01VsYMuAFXq8AFnm5bVwm0Q0jVRCrbhaPk7tQZ92ysg
RqTugvF0oGRKg2SrO1fW2IRst5NDNmdu5KpcHK39jnVbBNoTUDU9LohJj5wpdS1agIoa1hkadH21
zA9+sg8I7iGuWpvN5a4lc0hQkVTD8alkHXoDwllqsmkqkycx20Y92kaBtvMLew95in9L3fFkwN0q
XbUvcA14WWoqjoJzuX6DJoMHe5ZdIp1wewOcoB+hzYhCwuixwfNo9DiBtd5lD1r9bP1rHy30e54v
v9SJBe98sjHzf904ZmrXNou7rBEc5g3P30rrrlFoHQ0BfQDbb1HMO+ItpzlTICjAzRBTCCf2xPxq
QWrqHaiI81PlZf/U6EdBTrmtHCCKNzV8zNCM6gH6k9vEjD08B/qZegSWlmPa7TrOn3YUu6YRrSJL
CAPhy6+kMEqiOmKH+9n3yyInyFcJylVqgRKvrsO+29WqKW4dudPcqlylJe9M6HoMPcTFEt1H3bgx
Xse5PAr1SD/h5/c8zIRnVnYuVAXCMBba9nYhGx7+vXTr225DMieSsJQGD5VLeDyPDujxjwwjsAN+
s0gjRGzMowRiS5x6kTsQnHwUVaGFbea2mmizRWABfxKB1knDkw5vlHcvcZBFBF5ICKs5i/NDzhTW
utjXoqDUzvjlS9RfUpYJ1X7XTyCRNZl7mR3sT/umH8Zib7Ye/0M0zxrENF0Jm4qxx2KX7/9EBOLw
9QrspvaecJKdcPx8wAedew8LVlTC9W9jwxLVaSbC/U8+ceMAokkyjQE4AyXDqLNd0bJLqWw/m8Mw
9pZaHgW9c7X98TQO/3fk1Y6HGOoYHK4ikfr9JLPYUZGWy8+/e3Ahbs06Fwl9/M9+c7hL77NjN6pl
/CzzJWqWDCpS6hrcNgwLkXySf29BSONDmmo5l51i1ccSwM3CJnZl/bRgSUklS4Kq4tTpkp6ILQ+R
bQ254KaHV/BLfDLaZd0zGL4N5NU97gR4fh5a2yRGDYGq+rPdbkjv+aaCgmYdmcGoQAGZEaJsWWmE
tXxVjrODP79Qux7iEF3yfoTe48+3ReQFimcPkqTnh+mBJOB8MSq5gKd7apml+Q6JCIkXGcdx+jfI
2THURTvOnEO/wLGi8G4mduJQdUZNv0++YOy+lXPnh8B7WQF2mTdCGe+cfA7thyL2SaX+qdQnyAu+
2O1Tzm6OkLamI4sxr7aBdoNo1ggPneHSv/x71rjR98WaaoZ93YNAnyacU6l5rFl2KTef//Gi6qn3
2quWeWfhMMSDKh1Vh2JbU1tzFX+7DFN9HIvgzujG18xy1OYY/NUlRxy06NBKXXap3lJu7Uo9+0yi
ZWE5II2pRC+mbZ/p7maWCn5FLm4qcRW1DYhsMOvGjacyI2jBaT7JIKK0m+cBqEnQSPfmuMyqHjiT
49fPQ/e+FOhK6puG0TZ2GwelXqg7gx0UtFtXX2/ob3kUyDbLXcD0ab29V7rIa61E/bhO9gRiRBlE
JmIhC9ct4cn3Pdhsml8jfKyj0PF+OjewmGYl9Un9wPHKyu5IuajAIG67xFG3j6pra/o8/m0uoT2F
C2y1SBLIQeafdtf+rXo1Z1FZH1Li9Kwx+O6tmJdQ+ZQ6oBdz1bnAicbEPJZ0jjRxRgZWlalDzmHq
OfIUs27IoYh+BtLYegpI7MQQZLhBg2ZBEla4TIHg7H2/z0GY6H4tkx2/4FRyThX9biVZcTkLqGvG
SA6Opqm69+jLYAfF76zvaVY6lM5rwaOn8v9svnk271cVPQoDG7B9w8v1JMY9Ih0Z7kTgpF3Fa3Ob
ob4jzDqzmaXD9VaLpCZDEHoC7sA4aurk1q24x3nBqFFB1YQhuu8ZmCW5BGaWOwDSNa4YtDxs2rXE
6ewHWvsM6wpTI2ABvn6BWhBkoygO/om5NNTPXIZ6nytQjJpjBVVVd9dKWjk9xrURgtgQjbeTFNDF
PR+94HZJIPye9184sYsO6bICZhgjYM5U9Qf7PCRvXzuSpVrXCVeuZrf594sYB/ifSNtpCqdtMd8T
F7NHGI+TqPkF1DMS1oLSOd5ZRfhQqheWCzlttl+MNIPFi4lhlMhE3hR+I/dbRyRAhLWeEjv1XHjn
9yC9yZr4yGP69T6hBsF6SNw/K5XpIYI9BanQG7GfyCRpCpJq2RuY0Eq0XVfT6C+2Z+zoVCHdBclb
M+FeDSNd2+/Bc1n2JctQgfJbeylfveVzds/q1ytNZUyvfgMW4Kffup3Tmpj5xEu3PZtYCT2IGweT
q8VLwGnOVdg6b8GZ+T0Gt8zCY2uPRx5VDScOHSc2mH10oDTCSa8u4mpwopeTEeniabJ7pybqd71S
ZU4ZN0T4WEpw0bYppWOgSuqNQ7DGpJ4DxH14wOY7BvZpc9dZfEO8H+JmDPka8klRDWcOilU1qA8e
XJa9/PhsSNSW/GTqfV5xzgKlnmBaamtTNQs/aga2goJEEU5TvIzMVk8N8RuHQNI7RB1tjsaW8oEP
G9XnAdfzCbDgVt2iPdbJ49uIsTVtFt3qUt8dyG+PC9F56NRaA3A9LTSdYDSz3DZJN/6S/QLuMlOr
55DvDYlZP6wPZAkWm1XZjquwSaiB9opT46CWI5Vu9+R/h5nLVPAHaSCFLTaWMnfiGivoH8Gwal2x
ysdBBqe7E75M5ikOinUX1MwJgiFbZMERbo+4VKR2T+RSbGGCDsZGrlfHJ98zJBAdn1yoPun0IwOT
0KH+F2s0N0ZrTqpNbOh1DseZ7Lrxdx1MnL78T+ZAd6tYu+RApG69tXH+cO5AJjv38VwoGT6Gj7OU
J5piRilpxXvD39S9XGDmAWYdQtpYBnZDoGnlKwaH2sbT9ALqb7OXkPxP1etuA3hLdvaJP5fOEFeN
auv00RQumWZOx3n0Zudyhjv0kN0zHG2jjbro+CyZ0VrHiL/IYBkuwaIPz9Om/9p0Dl5hEqvC0UHz
kMKVh/0t9ihAmblfk0wpCoQqxelWnn+ESz69tK0gA7kYcvGrggwpZOCytO7PRjB3m9fg99cNmv/O
j7ziqUGbfxpuzOb7j7Vv0ny3+rGLHY/N4jd+wuFTfucnzOW2iSScks5eeTI2dV/w5iIKgTMYcGmv
afZUerYanYB/hg25MhFqK1R/XTrvRetsxJJ39k1HUie3JOcX0uTjVJ4rLskCxF0qYi2c/ZZPQTqx
p3wRS+G86iaPfbaorkD6jdTvHTkgOvw7iB3P0buu7uyUXjY807WOAkcqBLs1EmBxPrl/fblhqvix
uikLYU8fSPeC1T3B9Nm+fMw7A+zDLYE0XOb1eKk30ep5YzUiwwjaAt2bTv06jc/nYrAqQb7URBVa
Oywj+MWQzvuOMfZ7C9ZUOf7QXTdMSXsp1h5AOWkwbSFvjieX9jG5rsifTfeg+10Zr80acCVs7j+w
yH+qiYczKxxMfm3YOQVTp7B9XPCG1IkYVgIh6/r/9lyQU4LsIm4s+Ac1lw5ou5ztMCFlJRyW3onO
lvBJN5dhr+oWHefZlZg3iN3JQfhqzFGlnbuF0OOh80fCA/nHLHVW73To2PeGHmN1wASlDADqp6t1
84GbIJGdzO2Qaxz4aKY58wk/20oAltNWKF4lCl5e8ltT7lq45jRrl9RB8qjMNuK/P9wS0Ob9KUZ4
x4wVI+BLNKr6Rm7SBLaYNNNKk0udBG5oXhZP3GnH0hq+2un91P5RJE7azW0tpytLrm2/ewwJqUZW
ElacxD2IXooMsjEdcnvu+6BkVHzFuDLni0VK2DRa/7eRJB3Aw4aOZTNOTra0NvlDHBkM+h6mY4T/
GQTKhRhKpuiRcj9B3yCp/UmRCMhcV17X23knzCXIdQDz7K5/wXODTdEPlwmIriZ853RapGNbeMSC
BzqefU4mTfySWgQlZyB6akf5d18Y1ZVHJNs11Nxnz3hiyoxH4qzNox+8iyRQzz59+Pi8c4ZxCWtF
RRWBjRv8RPGa59+FcpnNgg4M0v106/5uya+6ARV8nkfxMLtnDXCf423PWKKgSXnWapx6delSoFgx
CAieb3zZtyt3wKQW2oKhMlEtotbfMpItx6EYl8EqDzCJWcsVi3CHGqUtZq/zOIt0h1fC8gYr2fLC
YxVGtbzTKYkwA05MS3qI0nHPL68bu/KXNyx8ecNpvqtVF2frgTt3Yo8D/oasVPCPMeo3Pq54vD6N
FKM3zRY+sEOk9KUArNlwjX9gt55iuht0QghM9S9yU8T9NL89MgrVm4nLlAoVNhL2IQ2iryer4vWU
ALZ01v3/+vo19TXRSucpUHdPHv/lDDga4FkhWQYI0yH9dSAC+klNRKdZKY+xRSjYD6OKzJGzs6hp
ywpgc80Es22UOMemgNhLUJY861HDKq8mJCbUyLQikYM4SNrqQUGmYQWsTBYUxUlgynvKkfECCmS/
ngqJhQYK+BmOl9gFHuyhBNN+qqFhsfNQuF9YHeSyxPk8GR3JrPRo1FEv5j2c2+6zYybN77WPi4Ci
zkGP8nT4FZ3bXQT4VJ6bERPNBhoWRFVnNhlVCDvtBDCY15bNsOit7aImrj5CtrRZCKwA/D/RidhX
RQHvk026RAgQXz1bG+avlUP/CLaJwatlyINoJCJKltOIvcfsAoJdLJPq+7Q58d4MZMFkeqDNfi6s
HLARgWnx1caEKsZxiR4earp5HhLgjNVew+QsncFIo75s3/so4mj1TlqNTjflO0tNZBtyodTWTZhw
6UCU/+VjdCsyYVtk4v2PkaGasZGTScrW124BAGlPzdndQxbJpU7vsfnvnxMJ9gwLxvJdlo2EtKLX
/MoH/EGXawa/k3rHr4XfUszAQJ7HVIhq8aP2BijKqAbsGVaVJ+Zt7ctXR1fF8iLzkaD1e810dAOC
J7GHj4KikGD2l7rLcmGF8F10ZNXMJAwHEbkebFkp4eFeveqzArEB9aKIK+EKHfc+zO3BAgc4OlgB
808jVcO00xBuuaXiPJn8TnVgOySbRdC2ALanGByIOG5mk77BoUIDUVXFQVD43YUFaTtSqRC02Lh4
Kqx/sSkCy7kQcpnUzW5lCQNcI5tX53hceOgA6wJOcJbYe5EJmBBa1GnkKDSevPnhytBLfI5qJPEB
vslXBLDqzCRbGljVmXbI6gyOHDxXOQ4DyoftFs5IgysonIEreyTEIUQQNKwxMXm77c9xPJiifa8h
/fXwY0nITuMAfqN2qptUhNmlqHuHYL36kaD3zCS7dcQ2D18uTzX6vuc7JPcToIf6r8gtSP5968V6
nZQ+0v7P97z7McSo642jakOT3F1+qzWjJw2gOvHXnthPB4iuz+0ZfD8JoUGR
`protect end_protected
