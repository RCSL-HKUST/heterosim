`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZLYzgQPGbZI0TaG3HY/e7ClzbxGEOfk03Y9K5KPf5Yx+CnQnEtPztsf+0kSQiQa33D1YmK5H/B8lkgGvvE62aQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
llbqEMDnxKK/7308gj8aK7ccPBEEW5DV/lFIt7jywOUCdUlT+91da7sdBO2ezYb1Lb6YBcxWJwA+6cctU0EIk9SVAkWazKaoixGxoqVHD8gLpjvCq/qUN4S5/ai40An94059/d8UtE4m6e2qWVgchwWXeOVzaXHdviJlJJr+AXU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pivI0mFOS9gfe/kzYyQkh6HeUOh8Ab1O7cmYW4SY+/+FH8JukDKAFQ2w50mnGvnzEQ2N6KId+yfY0H7wNAIg3PR6Y69TbxM/VNGnDhjFVkK/+Zo3FyBCRlsRFDl0eV3MDlo+MiYxoJII6oaiqHfMcJIryaTKaWPdqhjnmApZKnIJTtpdLQmRIas8lq2LB31BmEbUh1ZxgtPYpdHBZYyaLlsu8fcmIaNrw0f9NniY4oas1K+LO8+7OxfakhtqUTu5vtSWKIGbIfCfSt0WaQiFY5xQLkZchexTQsW3jCeoCr2knZI/1utxjKaDf19Nq6WV0AicmYyxrPptkF50hjF6JQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4oWGYsbQiqw9Kgtt9bgBTvblxL4PSBkA3GX+dliwLuYaIPsgLQOylNsTw5xHgHUCgNCLSrKUB/0Q8frPBzdx9bGwopgDp3AVhflb4cx3loOjwczDb4qds/hCysyHJuNyja9YcckBIV0eFa1GTiL9rqcL/fO2V3aoRstD+4g8nPE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tm9IsR2i7xHU5/y2NOHyrqARq+U/CM7KkrDbAUlFV3hYkjMS5jedUmu2aX5PRSitFERp8P0oIjDUq4jFJPEj6Uec4ko4f6IW9vNSxjOmy1dD0C2HOPXbhYdbA4fWc3KqYfGsh7CdFgQku4oS9CgxLn02tkWtOek3V6aQZXBatKuF5mUYJBZ0sitrHO//XRNkPeaP2VjC/Gl+waGgIbIqDUjGNb/O4rCFqyV3xJtKTpx8rcYr+ThbgB2zZCNsRKAPhHub5P53LCphXrYOulJyQiyxdIU+iotOdEISWQ4tTTQlKEmsetRbA2rQmf6FBynr8iFwd2EE0nFrGydhBgJDVA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21321)
`protect data_block
p/CLK43x9AW1FCc4/xnBo8aM5O9Sl7zCl+Erd7PePxdTOWibcZj3WRk1wF/u0tRrGGf9nZICY7mY
zR944WCbw20llIm2+zL05R6DPXqJGcNS5gOibOc+B/JeeBvfmUnLDLNmqX2o+RVnMkd0+9xNe3ci
ThW6b64CwkgVrjgh1o6ZzMWYL064eyJS8JHiuF7KWWXbiYQvnkGLl6HcKprlHxQ/Ns9V/ej+LA3t
YwO4WdAx5kbzv0fURMFJf1EmJ+hooDUGN2mMl64WrUEOGXSFTnWusjoP6B7IAxTbNXoivRgU7k/h
k0hlW6JEBpLUmmE0SA8OYEpLPPGZpla8lJ+X7+/D4cVGO8ET7DKSpeMJNU593XHshujqsinttUzC
lGSC500bWS38nbaTkXQ37J5Cbqgsiu+zJoR9PnYnbzu7zofr3UqZNE5vYNlRAK8O4qwCNWqBx+1l
tsjCD3bgnhScmFMgkuGbitm9jJia1vz7SvsEgCNo12leRl4a3UyJsRLaV7YV36ggCY4DdrhZOJui
C3X255B+koCBk2/uFpHryuDWtw2orelfNTC3Ue0hbFlePFdkdxN0mtNThyq9elOsbajbjXRKkEmJ
iVRMb8UrZRdMFP3j7YfgaYZaDug0V2AMLUx7ObaAX+lJ3rabMo1YS6TxoaPJQ0BbBAOWsl09TYr8
NHmu+uBVY1EujrJELC6zujAdtdoAQ++Oz9NRC9uV+tHsdCSXtSrujJy8IwO7gqqtyqUEBzkegQUW
NKirZDLgbJXRHHk48tNJWt+TZj+Npj9RnG9GywHEjOocAn7A6BSG4/txQihqgTpMOUdu9nYC4mZq
YLOS4cKBu3hUCafc3Pc2yZfw/X0rk7h10eQ2VeNQBDEw4wW4OXzsxif7TRhpxrtDQ+i3kGU1xwIE
Lp5yxQ7kRsEiPOGMyyNH5FxSawe7oBsIs8KCIGuA+mv3RCa3wqFCPAQYvbBYS5t8OYDrpsdYbXAx
baSdPH3euOMeW4KwbFFa7m9F05pYzHAMiLhfNuWjSsikgZnns7FfNwWunXYZ+QPJvzVaEnK7VoP/
T88JnssoERVZB8NJM/T8l2kb6N3/4CT6f0hPIvYbP9k+LgZnOW4va4UU4CV8uclt75drBgctTLDk
WffULTJTEfnaMmaqQGD/zFM7/esJzbl/RtCV8OHVpdwbktFF7NtlxM39ahEEeE20rwAePEeTUQi0
Gcyorb9omWXTJs1h+VgaFRtavmMh+zVBhtDpXGDV+luxzpW/fzcdR0nBcoBC9/bK6tkrcD14QjGI
BHc6sTKyuclHPaVgc8T9RJRtqaLwZ67T7lvx+mB+RCpM/0AIAIVHMpxj+W4OzjGP2G9d2mCkD/J+
AKOMM88Kqzoqwhi+GA9iDbTNHwpibW51UclXAc+9WpnOVJil+ynGDRxK4xwR4pLU4NOBst2FEq1c
XN2+CHpDkeeTcNwujO6Ui+EZPx5lX5AnF0hRQK1PPojGuJnybw6FJ9MhaXqBhZg9GtEFPL+B4WhU
4eZ2CVi3NHkKuif+aH+7a0rkMzGfZdoPX5msbCrZf5zoM6vVqTMqN/JK4vldQFa7Tzc876jWEQw8
Dp6p1OcdpMLkrxzwqnCXotVuNzeyYFIXro4k4futjm4jA/a0ggj0PMpbfx6yw25DTVGHIqtOlm01
UJMx3DDx6OB6OrGvSEx5F30/Q7Kprw+j9LVfq/9Vw50R0TOML9wkcZ90sjkiKRbnVc0u2gjE+Vwl
96Zzvsnmyl4GErOzKnMYmAMchOvI75Y7kMBAtys3641r3q0qTnkyzcOODGADBcW0Zd3vs3yzdakP
I7ui0irP+g+SSw6NBvu4htM5012TnapQ6FEjKlDtPiSc0AD0AmSqGRfpRCd1VlBMj7IeM8VGuA94
WaWKcLrPZwKf+/XRzqpsfFFNfjszgY2jjmQMAmdFujWzbOnrbyXQ5DtuYOHc5l6i0Nac8TC2G7Bj
VY/F2WckwQBhZj55znhCbh18tFisauWNp2Cy7OUi9qdYT1uHwS7Cy6lclKrlBFJElb95Pzsc70CL
mw8Uu5b4fbMWxOtFtgb2kIctdQZmYa6OQZet+U6Zkw6zc+VBS50nt8YKAj/xrdR9xDDpA2hQOgxi
TZP4cj/Rxn4u++c0GPVKyLOxP7YgSwyFBAag+pEheXRbVon1XTGoMZ8PJgcoKtvsVFYFncu1o/xo
vhrao9NRKi85Ygv3o6eAiPVIm7H/vH0bLMW0M4wuZ/gSH6simymBia048sny4oY0CbNu8R+Milf2
pbOrC0GDVIxMVlQ9WfD5noznmor8HWDCvU/SfcmqAHI0yoEK2QtTvCenUSK1btqXWSLoFEHjTMFI
o4/RcCzaow9RqMoIaIWy3IxjhZAQN3ATs1V0AFini0VmeOk2Jj4CMqU2Qh+je1XsOfhSHsHtqOks
yhGvDKFbaT1ln8P1Gl6rQN6mp5oo4/mvpCxG+K7tOjEp62MbtWfbxYItpYrPXINyp8g6N4BCsEok
4ndN7qkrZ6pdDKoQZa9wYYOdo2yH5i5rpJSkD5rVlCe9epEnMctFSkFNaeZpGysjfv5pSqgs3Edn
TwCZfnbZpBvZkuqcDYkbNplBIN4f5tVkphTOkNKPiBaWZTprtq8Eg3UV7ZNOTpYcN0xWAbfBbPhs
RX9tNz5ia1dzVl1vK3MNMtbX6J/D50uMd9d8Vljfb/bU9mfwhVNuVyyFkMWKpHWSQfoMRAy2SEck
YV73qcHZweT4YB5e3FESecNZU0MD/k7vGgIAxmYtr9QiTMcPoBMCRP/zQhPnPejIxbjyStXk2/v1
WnVAFApYR3m+ckM1/0i4nnD1w7RLA9VePmtBZqVUgxnImFbsRo0NMK88mHNSdJaWre/jUJ5h+cGD
HtGuiFinZYf0zJUJWXsF7WH2JR9J7C+ROjFCEaOIZBVh0QWgsk5BksMsUMEdWtVMdDeSZVuNnia1
byfsizKLDmA7ekxslLyK9hT5d0yiHbWrU2g4/TepYBBU+WCT+mnYPD76mml6c1W/PHpp535Jo5jH
RQ1cEV/4cF8GrMt7Ith7K6IQBZ+oir4I7AOu4Ub1x63CmukDl2HvzWkPzmzxIl03zRWrPVoUPULn
mLcC3LS5LhgcS5crC2e3w4bWIzoyoyEBzjyXP9V7qne1vMCaTSL2h/LHM41B4ZFXWpU8pthXXbhu
+owT0EGrenapQyvdLemAg6RfEWca+jZIIDrYjCbNdazwq9FF5fpiT6FtFSjuQtuGaRALQUgZFPT4
sJEdvT4FNPg+vINCP3gZuYTtiH8bUkdOH1bip0Q3d+DjgDCEHemD2C9g+3R/gtqQqwcuJK3i2bZn
Y6zvtafhKTUVGBsbmoVZ+t4fFexGiRI6QdBAMLeD0zVSIUldNJNO8HlD6SLZ1Hr7prCbIybzq6kM
Np4ijVM14GS4rE3B31HVb3qBhczQY5bs4hFxMYIBiLB+ZXxmv1a2tFgM227Q/H8JyHaQXsUtq584
88/1OHtIRkaFs9b7nY/eDmC9sNqHpMmB4QOlxED9YQwf7gFsPq0xAG1l48DpMWlfedaFlOb2l6Or
p2Kz55UEmlDJxDZKVcKtNxeSXuSaZtOA4VZHXcrNRE81e8/e2HYfk4f2YD6xZS8LuEjXthTptKJX
lKTVm0jPiJzEg4N7c95fFvC0f/VtLSZCPCl6rWqqL2GDnhEAW9ndUE/RSKxTChhz9ndVvQZQMOa7
s2pp/NHrwu334T/0J9KxBwurv5xq/7SD4d5d1tJANIX3CKMEwAMdPGMsoh6yvOU11eK2jafFBRi8
RQ9Y4Jdnm1wQSXyYxmK+6y9d1sej7IirNB3HD5phUUScllnJ/H2pYEhKWzXk33DmrRnTHrMH2NjP
K+6YnavxLm+uH+WKe/hQEQkb3itA6oHJPmxRy3m5Oa3Y6PQYKkouiwQToZcCTJGzE/rhZnsYznpM
mAI1p4KD+tSgHSwpJE4la6eT2Re3zEk+e0p9c4n84CxBI6Ku/jI5aXEmbfKSBoKQ/TmBylUWGW6s
1Fq/zlhQThvM+m2xJc3h7Zsn+AR/THOudUoirG6sfbaX9lMzqx0EpDElp8rTexvSrmkGMplMhCYj
1vNKz3urB4zIbg/k3u/N5Glub+tDJjjrCS9+KZ/iqPg/B6gu740NR2LR4qNA2CHy+ZE9KMI4MTDt
8Vwb02tCZ/4vR307/dlEM6wEKVWzlOdTLhG3hQo3/0eytzkmN2O5Bwm/BFMpOvY2EI+KvFqLRa0m
LwQyn64z4qdoWx/Jyd1vbQNOe3ARY0uoF1AGxEhVtOxvl2jM3Bv24ybhxLfyHRwyTFlFiqo8ZiBO
IzRb30iqaqmVnUJXWSLk/CSfXMEPYBxXWF2BNDh9lWVk32Y1IPwVwEOHDALnaNyQmoaGKW2vwDex
QOXocZHYsIO1wBChtcgptMj2LW+39JOdBrvNGeRrgct6FpLXqj+DNHvGtWthXxBiQw8uoxTiuDRS
RoGSmsDDK+puAKT4/p2mV4q1/5Q/ceWGm/Tr8fMaWv2weozrJLVmLf1goR+0Zn8hToC9Qpka1IOU
c5tw39Vi0LnEAfM5/GDlGx5fKroL54RzOGq/eBvQ0aL6k55Df8slV1YBi3lWTvKENqWLD205uTT4
+fMpsk4efWPHSZQm8TDSoiA4CYEEqYg/5/FXFob4r+AQ6tq8zREUUudXxUZVs93dKyyZR1eQu2et
01Szz0Heo1MF0eMGTwiL8iDvn80vLKifLeva/Li6n9+yNYdfz0V7tmASQ4zDNOGhPUP4Dxz1aVwj
b4/fraUTVdnzcMoPtGHeDLAZESETmFukNaF22niWcOVy85DuHw05QRhZoABIfeEhUoSknGGT/d2/
G+Pjfw5t0m5vst1ZOJym0SRw3HZqaCw9hMGVH7X12ddFJ32kFxiy19b10k4sWwhY/lh9KvS92HBN
iEI+SkzLRc45K3dXSFuQgwc2cEU+Bsig0kLOH5i6xl88Od4nD2Qu/bViY+z8/J6GRBWezaTxL2kM
ifmKadzWgzSg1DI6P2NyoEoy2/JRnAaW90hXMluEL+uL1sA/GU+21Bzhu7dBeETllvky0+d3wy32
Cajw1SuLbwPpVKCj6Uoy3ZV4uQbJ61Z/6sIY0oOvG0OsoyTSwMV3M+xpcVQIT5aOr09zqjkxAw/C
EEvVf8aOckKmCahpE/jMpaN97120oZfq9qKKcn65IPmdmJkK2foyCowoW61cvz57KSG2rhridB0z
/LBr3hQrHo1ewYjmjqNE/1BQBG7bfgrqXVlhYZCINLZA5GAy3LqiAe3LjZzRrBkOQUtg5xKXBvE/
KsuapioV30+ABxDoLDNJZrmQommEO4MsHrxD86rClTkepmu2hMO+vsT6urbZ4Aez2FG2QfsmxEjO
Z8yNzHmLoNghh5Ts0pDDDx3xQjeQ5MI/v9PN11CFuJhOeCDLArHwRSvrpr6a//ajryoTjJP+wywY
C37vDknM6Ilzb/vDsDL4M8PsglbDrUS+WzPlDSxJjnntTqe3aFFbUzYyylfmWJG+a0V+ulL+4G9l
1siYZ6XuI4x8gugwkNsbmMTSIlovoccThozyQRosJL9DudwDQg1HOAiWk7bc99Oh/xWcW/YpTr/U
IOkd8hiuNfsTJxAi69mSG0EaRQbOxz+y0WcmuSxm6Jf8is5Jm9r8abM6qPa/lsJQ0iR45AzwM4fj
pGNnvdoMXPA1HaCKYi56xO6doa/yPFiCEkdpi7VkYjIht9m2fDXwMY8r13mhOTvp25htSraaT3de
+2xXu3VteaN9T9DORd1+HdjgFmD3OFfDzLG1iVgyrZ+rsH0Qslfiu0R7gWLlM4a3uaE5ayb1APrS
Admgm477k2/0C+c7bI96N4pIiFbYo/JgL1VelpQ5IKxxx/DL23BExTWGs0HJ0y08mP2j1/+MjBcU
gtZej1bts88wG3dPUuT5+Vw2BXaG28Cgk20dB2NhsvJ14wPD15K9e6A4/WDLqT7ebh43ghF/TBLy
QcFwq1LdOIVg3XOzqysiX8OBrO2xP7HtIKbtP1Jt/vkMXJiucMggXYgqNZjrTJIMTqL0k8XQxRl1
AEzxj1k7qge00od7n3k46jXD0+UniVUeCzRdOojtaW1CkzgZjFF9TGNeS6/po0Ezjc8zN2KxjORG
79WHn09ZM8Zs0wnYdtsOdx73PLqXeg1syfRkxnOyVWGGON47lIS+OWYmjffScsqeqe0NSuTiqxbh
q4xM+7m0yRAN60p362bqFjOgN9A1oDmjDVQMJZJUJrzp3EElDtKl0o/kIhVYVijTFigmR8O0iI4S
x4sIyYsfE7wCJBPaQ6saWZJ7PuKAoqA2NBuMj60bdmfvJyaWGKWpKBd6cNrDRLPPUcg7XvZb9HRX
dQRqBxPx4okbNbvtlAqo5maG/9Q9G3mjbWoYnGhXT17V4IFPfxP8CwmsEpPbTixoXhVd0iIFOG1R
/4ycTr/1gcKhk2wpgMVu4ftfBNKnUHOnvAtBrJiyhWODFs8Js0WdXB+C7qfpOWwLCksP0Qqu63RX
PyIy3rw07hJ4xI8ZCRcSRILCnXC/Tpq7Bko46pwpEnNMSBOKkWk2gC/jH9elachV++eSk6ykafrZ
DBfxczWzpNdxIOhIQXsuwM0SWclY75LyMxHRRr8rbl7RNrQi7Ob/JHL1DQzIcuLkXP7Q238RPiuE
BmL0EyZXEUDQ+WzVjcqwvRy2Wl0ny+VE2CIa1349sy/qcbfjd11vJ9gCGMUXzQlx2WdHJMijodYO
IZ4S0UMRbfO8jbOTcD5+qI4crHGbtdqnJetQZila1ZmVihmVv0WmthpPNjPQcswH7GuzQ3olhqfA
9mucDtJXLgVS/4zu4o67qYbuMgY7chTIhNsR2zDjsBKhxrsRKymBkJfC4H/VP+WaVWFkO4ac62J9
wmV6Ki0g0QsV/l2eQ+wwmugWo14E3krf86rPOA8ihIG8S2e5J1z3KlFMdI7i7yvOeIFhHYMdfiJY
mT7poKWzBShLRZU1t9F0Mj3LhzuzgiUjNkvvsMywCsICryTbQGBLnLA1ENTmR6OsvYhjQRZ4iA/U
rW/KIFiUj+JbQkvV4lPPH14JNfKblV6Uh5KhSrgnj8KAuRhVcyX+Iz/NKPvQFVV0nuj8VIQfShRm
5pan/i0VYyipXkK9Dr3Y2fqH/tpXM+0X2/X510XGWYZ4eeOM1npLXnsSK3br7gFuHAg8CpfZ1lH7
LtR26zQPu8GEnGce2PTkLiZJrWMiAeNB29myvMZ9dV5cwRYhKRB9Lgzo4iu2sCLFkHkDRrTXHimh
qjtmgwECXA/Y0x8jEVloKcteX3juOvBGfCeg4bd3S/XSdqrJWz632rKZyFBsWqiWzg9fJtGhmKix
DT02kbFgIAJ7nLz8C2EkMcnmammD2i6XEFlHWsPAIhgWMUs/9ADIMY4Rf4/85/gbG/vifdYsw7C5
v2LjUuEO+rAORRKwRz8swpZdfUqvig+RP1Lt5HpFYRQ1MIsfBGi51B5u99rzHb39bioWo6mzT+UG
WnAqZVv7jNc2iPOQaDHn6e9845EhntXxECLH8IfOqgE+D2HIjnd8x/q7+Pkiyf87WpvbDZBgF96o
JiBUGJQh42Rp2ojBEM0Jwip2DMc/a+o8PM5uPDQQyT7b8XGM7a9vGcqw20QQNoLYhgRVq0OY3mS4
mwABpMfGrRu7D0IW/mjDC722Pgm8vwx+V3whJLHOa0+JjTAG/ARvJDFny1jN8Dk9jn+iFwlZ5eOC
pKhQdU4ZdtPXlDKdybQAR+EybGW4C+7fnFj8vQjOI2bYlQHhyiTYMyZPcwfZxW98uDB/XJVXkdF0
rmtKNzSF4LjIOyc4nQH5zKyOft9ffwL+xAjazPHFJV8gQE/VA333877dsgWro0Ccn72h3wTkL5xB
j9qkF5qHXdkSINj8I8fnlFubhv16wnpGy0IcowWH1o/rNMgv8FMsqbh0d+Om8USo5+QGkXMgyHNm
4TzwJ9WDvmn2VG01He+vd137Oh3TTAcvWeAGjVgD3vz/UP5JUYLXhwFjp7+aqZHaEKPd9mJmmbBG
AupViyTEXa+PAyiOq1hyZWw4/JwaXp0ydgQWsz9jRzFlHlLeWVZS7PvxSDiPcZqmnrqEMey5KSai
MrKnubq6PUbS/B2S+fWaJbEZwF5aCCbUxzUnrwzGSDBmfMln9y3IV7ndeejiJM1bOQsP6i/sQogx
kCNfFxoTMbcW3/hjM33GH329RZvnR+zgrcoYqoq7SU5+jg3r9JrNX/LEXaK5BLUS9DVviYYHU9uR
p6mdIlkmX66gjKGcUpY/pjIX+bKdkBWxMdXOHTHB9eSxMipDmsXS1AyDCy5guBhHcpwn7CHnbZ7g
et5KOiOBOGO2/9Wdl001g3GCY7lZN0lqz20rD7aQpJXLBxmAafJlhamniQX8qvkv3JbATWWe82Vr
rE6u64l63g+j2SPXFsrMpv8jZQ36kljPJnE9kjdHg9nqNyFcwHL0i/XbE9lf8o6p/4+DqDD76vZe
vO+gCcgkd5Yl44WvASqFVK6ways78coFvi/s12G3aSTg8pt5lg7v/6o2CQTDB0NURjGX8e2vSLsP
D5+zw9T+AQ/vvcgZIpVQWE4hXeGQ7l5u+zxtszUw72pKoubJYWQmRJYr+NMUM5X5Sl+zZ7JbHWUE
OaPflC2bi+kbl9MflD38udAKgWZfVqMO9rl3esGlBdlWziZ0REwOI07nHS9VpuVPsyGVJ8Y3Ndiz
3OR/Iv7jmAPru07xfdrrFvXZm2uhICSS42kNAhxW+Dry2kWdQ7+uoF+Aa7IUza9x+HsstVchH2wf
nLfgkz3pWbXJoYnxTViP3aTNTF6zBRAxNtykbt4bkw2rGyp7t0ahRD+DHNyZ7O4J134rrJcnbPrU
m2HzAOun7Xad1rsWxHsvTM8/VvnNPFOTv1NuVqklLLpaoc9Kz029d6qOO4BDst2yTRkQcraBg0T/
OGuG6jbqoxvqLntEBdXOlRegnaUeF4K4f9qCMuin5hC005f4CHcAWLQgfYvGKO+6K+CSMgAJqRfS
tK6rjZhOi00ogt8+JGsk0a6uqn58umdlQ8bv1jtKU7DWLWIPmJ3dLJvzHFEgYpHqvmPvNv5RaGQ+
VUM6JDqo1CyxSAqwhAgaaRmbRa7lx6QWThJWAlaUwfSxia30tG7EHP8NTOP4emjOjAJH7tGAa2/Z
H5IE56teU8RNIKuQkwJMlowstxJR60QLV5nle4QOH47T31V+s8PMaokoiQkBlKMM2ley+Wd1OqKf
0opJGlsXw+XqSIssgea4YkUY2OtTNhUSJ3EvvtUzg19/w/x/mmrWRj+rt9kuxdFkRsL/e103nlbB
kUZhFsHkMvRLcxfZPi6JzmMioYbVH8QFiuKRTVxZZ2gqilbe8Aciq7VK8rml1PPCXA8esj/GxZnH
XllMkb3Tg4kbN5hRrZOCeIuut/h/JfT1VT7wDw/nZXbUnKwN5jKmYgL2TFS8oZUUS4ZGIVQfUgoe
Wmy0OPuwkrmbED+Gjgzvc5yvkEjb1rjuVsR9bGpQ1MkEZDxIDi0ezxfMlF6Wt3Z7fnRBJSFzkmEJ
ggUBsyjIwY0EyzjqMWQ37GIzuhC7spTMgT3irq8V72Ud8jrHfpNpWQFZPF1X61Q/fvEcxeoRjb+V
AAeVaZ6eNPICot7Rzrl9OMdLBAF7p6fpCrTmMuB0oEjGphXZoyTVfgRjbe5F9ueS/G4ExA1Q0FCk
twD7AHsdZjIogtu+m8S+X2SF1BnExys91ZqnlMDNdCErRGv4SDYrZ/XDKhyrfyWI7EY+RAJq+wiG
HEYSyKfUkxV+BnnxhauhHboLpye0kNQy1fTwjXZX8zoKnNo/DZlwqa0rBtSu6voI9wJB4Ow6aiBe
ganb8ZFr9WLALnvrArSdMUHiVqCJGmh5PeOdwaht8jNDbyMnEvDDHLL9vA6QhK1NdsLgFV+E1CaS
Vsq3S8C3wgvQ6XVUwN+FH38r+3/dhCzET004hHL+XdnEVn2tzQx5MU0WIDby4TtAlhG4xmOGCzvT
l+DeLaT3gq5WVhOHXWITjBT3yN6iVM4YFrTlV8kQ9vdTkDkYFknSABtsr9Y/zS3s7M3diqP9ylnA
7Z3ejohw/UUoeTUA9AyOIrSpn70xXuUJsny2ND799jwQ0SorwBh6du7DA92m2W2O9GISOguy15hx
nPnYtYWVjApRn9nj9Jfw/S7lTdXKR7I10L7a09NLa8I6LH6DrHGim4G3Czr7LCpSlwx7gbCjxzMt
3PfR8ZBxRF3h1/yeyvAlpjjpZseArCTn8dGVLZIQYwOYsr156kCuBw9t+ftSHwfqzJbdADKElM0X
SZONNKfOA6U/Myz1dFYmgfbsgSJCLkCTmvhT2jgwYgDgSBTBSZn8sxdHZQEhAtlMyEOkaewt9uOl
3AJi6XK3BfHqI968gVBi9S8T6G9RXb9O9snOH2PpkE84H1YB+Sp1hSFInzzF/7MaSkXs1ke3zi48
hiG06w6Nji9clAkX0cXJxypw0iyZPY7eQQ0DRkuaQfJSHaKikl49tJY8TYyP7I0VcqaQeoRkTJmI
2ospcp/YUvnJa6fBjK1Y8L7cC0eqjvlbfrcLO3JkqTolS/Qv5paUdp8Z+MKhN9/nxGCB23Zc7p2y
JVstYyaRchNsLSI3NG2i8wIEVtvND0AVXI0jFH1F/+db8aR6sNkYWEI3fVGeDV9/0ldKxbbdmVO5
2PmbghUVOTz53WoX+7P+rs0psPWr9AAH+rAy8C9Yz8whdCpZGRcoBfOhYsxkovA7TsseDzp9LRFY
TDhMF/4fj7/Q/fnpgzOQaFK7Bw8qWOY2ki3JMwkDDEFi4w9vN/M9ZCd/tO9H4BWEfpviFGV7PjtL
nExOM0VwXcC6wfkL/FBWzgOG6O6xeA25GRbCai2h7aA8pnZpHTrd9QKsMFNodqPvKIgwUJ9m4U1J
VlMGU6Yu+lM3wKpDwwiLPbdk5hggVbVp7DDONTnuAW3kz0aacSMcWjL83LVLG4BoIEhH78QZiRy5
YsKsyx/STFXx5ihJMz9Zjqd20ebR4yMRd/6oV2WHsqqwfuz9E5QIpGozBDhfVXbv1cJEF6VPb/To
+i+6vcEy+82jlL7l6IBtEVE9onTrqSPPFQEmYtLjKiQepfFao6ftv6caZGOVKgHne9OB8OrZLiWX
/GJis9Fx/NYoXpmbh6PT2ytbFBe4cT+J2V47eOffKAcGn6+Q4kD5/I6t3pdHOKxhJafZHYzrwzWK
ayfGuJhx6C5GSEbb5LT5PUtwJCliEg/SG+W02uL4czIZ1NqCdJ+WiAqrFgX36VQEAFoEavMGQgjV
9rh1359MNMerKMsxto6HN6XlmJXwKkoM2oIIi1lIkKKTzkIjLFmuka3+K+0ODTrBs9li/fPw/SDp
Sex0kswNSc8nhGoJ590hHSWJa3ZMZP7bXBazNI3u0IEgf5XQxprK6B+JViCh1Ab3yJ2BqbhvilLc
m9fyTEsAFK15MAu3NFH6+cXVxL3sZanBsaeM9SnbccDyqQpyJvW0YTf3Z3OxYP1xvlJR3jDNREGe
IrgYR/OH/t/D64zrH9r1W9SVwQB7zNOV0tIwljEyLf42Tq2JnM2sVeTP2hvb1Tw0binL7kEL6q91
DpyUHLDfuRB88JvcUF1pMrmz3gMbSosk+pcScV3/lMjT2kG8d3NnJyxsnh3bOUrWL7yRpuD8wQgN
WfVwr26zn+Ayttb2stVob7APG14D2zFFS6l6bx81KaeHUbSibO0p71PwP/i7hjCnUBauTrrJEkZN
RSxCwwSwQmveUJrjeLvfJNrZMI+ExaU+SuzQaw1fhY2UZyjvdZrfA1h2WcI4h2MSdinOg15QLNRm
FUigX35N4deKsXC7PYkJL6GgqIlaeofhYU2TwbVP59d/56RNSbuY76lf6aomigieNc2BeskkHB5D
Zf5Qp+xuLY10BKqIGhTTM/qSWuwLTol4GDpliZo3Fs888HE1B1kgJks2RnCd2ZjqHwft8oRPzQio
0leKI+/wqmnfxTEA47ryaMHMiS+7N54Z/F4+C0RRzqKO1oFSbHt1BzQ0uc5ZM5lxivM85TYwNOjn
S3OAMWVingjFiVirPDb7ID8+7NM7SMYqXhsJnuZTlHG9H7qF0ZEbFO5AmEGzVG7eMgpRSHJ+XEtv
F8DGfDu5bDunMt/J2eKcrM66jaICMxUgWIbR3WKcGTvna4U+m1LeS2Ik/43SwP/ITpFvOZRdPYsD
FammfvfxWpLN9lcyOFZOH+PBH5d6NPY7nkPRsb+MaElrbpfa/DD9+YyYN/0UC8Qftyi0DIbzNbAJ
/WtDk5kPF/Y3Crd/49v58m64cg1W/Sl//eTiXGuwgRdpnHWTvWx0//qop9XRmvF2Ddm2LIfJH3K/
oDwjxn7K4ELorMGbjjJNJhiYtGEgvGRy/0V6Q5oWEnERBLr+7nrO1VC3IUy9gC9O7Z3tUzqcqfKt
IxJOKn+brqL/G+btkMxN4p/SZ9nKdO4OSizqLehfBizTbExkmt41adfDTRU8Z/YHwKHjHeVl/AIk
8vYpPEeugH5HShImPf5SHtCoazT0HkQGzATZFsaY4RVuAEDKA9dkVfDozmuvpApN4H8AkrqiVM8C
HPUdu3XkIIO9iWwlOYJY5xgcSeOXzU7NsZeM6G/6EJ3Ont4hDf0Cd6b0ernm/jO1Q63dm6anbsAJ
bWKxw/wsz78d2Q6ab179yV1BGvv5ebGsXGxb67uOk0K4jA3Md26AkiZJ4ttLyqDdoNb8XYpfi0fZ
jCKbyGhTVTgsnZkjhBZz95BapcRhxoSUJuN1PAvs8Y5DLGUakajlChzakGKSlSXdQyD5N+1ZPkv3
2spu9TXoQBkQE1ZEzhm5wGnJE1f0eu8OeiHZf+UuCu1EolfQs/874B07jqExfPII4V1VGnmzUngX
4HmN8NSNuK2uxzimkO9SvBR/VA5gJQM5ltrcmylSPNmhDcsa3MeLjaJGoXkdoqyJ9NkKi1Ww4I9x
M+5BIos1WpUsDWgey+QORvnEcJOCM5gSkRynoP2Iqb9xPtycing5KCBq0c+OlzIeS25tDsDviRPX
kvQjz3iiCJrSpGM3zrSp8lQTQsLmnnX+yj1bKE/JTY0/WFjd939GHEnMxV3CGQ2fvDSML1urJvyn
X5m7SgHNYxfZdOHyOssjRKMnE2lBmzkpo/GYI3tuAD5lvpA5I2Pilt27YnbsJ0o1BHoAXHbW9bsV
BzIHVaLXXLCQXuIzLonCqjfZ0RfNpe00m+XmF6Yaqc6TycSm4Gi2nkIfKIOmKj/VkfJMys9UXZKg
Nx/0zLOohw2JQkmGsDEj2txZKCPY1d5eo7VzLfqCEPJm1sxwyju5CbMFrc6CNdFvRBIWDHKaFtVs
DvmiMHvgHHy1Pp9oAR8DOM4dnpqjw6SXOBtTkMgx05k+LXZTWBeX/woK+RnGfiIX2rWkSahk6dh6
AqoNFPttfz2w2J1Td2LhoB2tPKLP1shj0MJvV+4IR7yna7h8yojCmxEwvry6Kj86dcwC3XQZ7Uy5
5ccKNXtCIze3th9F856Lrwq1vgRyVazCWKvHOJHcGIF2pMoUmlCH5fnfengo7iu/t9V3a+ObatfL
UxDxxttxwkRasNHDKmPcb7jj1jDUZjYFRSgFt07pnwzOutPbO1Ios/10+A6QrUBuMbkHIn9ka6K3
9HyPdbM5ZYY61MlwaDGM3+ELgCy0xd81uCW/vrDcOxBz4cFSgyKC4IfxmNOCpJ12LjD3oQeBNPS3
AMFK9nW56tOmOu/Rm7mIZdudYAU4eZ2SWe9PtY9a6p8t0xTB/xhF55qxrCJWAw3vC8qMteud1Pkz
sgL5AYv8IyYSPh5oWEfWrmj1LhkkRRsK3zZUJhcX7wwImUF61JM2ocJYLY/cQrpaPqCi0gcz2SEx
f7YCcTg4zgK9qI2vhgYZkUf9UKscNNQwebYhJ4+Ui/J334kcX4Ud7b6JhU11XxlbL0QcWiI3QJek
FjKbXTwx+aqrO2ohCy1pS0tIl/ltfBOWCKb6Yy4BkU4uuy8exFj6t0tOYGYzhzTEUvHE2OFlaxNf
3YwFL1PfDOU0+FsYOioRXBm82CEzfLkG7dDQI3kG8nz7SQ8wlZ7zO3DGxmBV0LE3gfiWGiYO7++3
ZE01d0SlQ0Wu79E7501G6SNLdrX/QRNB19UMC4aYk17YD+uDteFyYTcJ4RJ7B0+WxfPU1BvHqW/E
cT5SoIwuWP3zP6X+3mJlqyWD/0ujFtPZd+xmYqssbBwpI8Zfkqn1hBNp4j3n28dP5ghRLSKW1dM2
K5D+yp/ITfZcVFP5AygjJScOJl64nrqfRC0y11sBLrOi5cyZGRNb4eaVuoQ+6pJGOfXLEfgmiHLr
lkpxjqZIEMNUMePwXS2nbFMiM7LdPUeVGRWz2ER1qqykvO1kR/vBBLgFpmXfow8yFcwiLGdptkgP
N6SmqI0sQ4sC1SKL7ank2JvJTZCf00b5mgLph+rDy5e+59h5nBoalsBnIWSnrFxxAbeLfGQptUGI
54NDAaW+pLwogGExkNH6Yy1SI/tSrJg2kKNgtHGUZfKqowS3pGMc4heoK5vhflr2LIqpZ7qA8Ebk
llxn9mVKLWvFvvVq1vXzJA33P84huKMhhcasq7iKtTTkB5L4b7fqqujPx27UsvSNe+auRI4rwgap
mvfHyjXb6PTWjKjq3eKPnIOp81W7JmzAqSgF/+GzEQqyhjOuIO5tCoQpLfXh7SPr0DSajNqGr1ZU
ajvz0kKdCYQdn/2aP5J/kHUV3KxAQw3Eo8k5aw8sK1YfQqKylE2Jkg/jhCB8df8HgG81Ljx6adUo
OIeedxvERzkvX+6ZxYpFbudSdrjmXdF632eGM+hj7rtITVp75eoOc4KjlPVSKnq49/kYxPJCSiq4
2qFYgWlkiAz1RqhRxSqW1aDoc5u9dT7zh3KqGzUzLCSmSW2cnUrO6Cf670igjJAPLjekuoMIip1P
3+OariaApjAttlRGGdLIhQwH4LefzQt1glTIkPCUUyegC2SJkOsKeEo3uea6yNcpNTGhBLUQXbQQ
wjsIICSJ41T1M5h1bNtg+PSQPQAOaM/whzqOWdk34M4hT7XWMH6vSuei867f98awdi/RsxdJyGDQ
G2t2Ryp6XD8Z9zTo/vX3uezs/L9WN/N53wD7GtiPicb/7ZvoGuxcQ48C6gmfWkYjGiQqCTskL58m
4cFwFZ0ZooYBfaln4RodtIa7cxpK6cU/WDFJr3FG1l6OC5nnVhH+yZ10lX24WHidkmAFAUqwMbud
Nhjx71dG3j3GetM37KNmhNCQleIK1rqBIFYBJbeyvETAylQTmibaB7zi1RmvKJidGgOp8w5M6asO
kCRjtbGxrXLcUkRDZyBl2TB3UDXne/SARwl2QmgJv3lPZL+XxqV9npe4a/4G1Eepn0L5vqTsa1iU
MGGjPuPe+vPA+o0p0rUN/DqRzq9OEvxr80h8dXti98F+iiy8+AN46Bjv8fqceNK8E1AIi+T1TzbL
RYZtUp8cYEEo22mkB8uyrzGG/x4UB9SSugDQ3OM5YcdGqdBUPTiSHYeqj35Tgvtq6MGaBUvby3Ip
YnNiN0qKguWnIWfjo38CaY9PPIxYgOzM8/6Qud4TkssMXeilQYWMJGmVZ+veuvMa2fnhgjouLtHw
aq9gHbwcU737WKJcnFNWLnNNyJ5b43RhqYvcEADyUFJyHo98kBAyI+6vj6Ksy+zt3NUE3hl0l8+Q
G/4UuqrVKanRuTpeTow6MVMKswergz28j6/SGOAGH8iRX6Pn6AedyypT7zI3fFor53x77iIHsgPj
cVYb1Y73akWEWznKX5puYIG1lyql67LaVyKZExM1S5jsxz2gFrCta5v/eSTIBC/pWqehvZ40Zm5p
EjtoKh9wfUPYHUVKDCfjcR9m/Z32YNlkall04Q/tU+I9C07ehFe2IVDDSj/S0e10i7TmAYXaAkba
fJEcNJ7OFeWjX8fzlonpYqg14Jj7y93E85ZwRCESL4D2aYJ2Jm0T/vZr7rGgQX9MqM4J37GfpIu0
3kHkqrmyiuoFR92E1mLZfhXVfM+06Lloq28vuV4c4pq7XygI2RUEGl+oAtHA7Tn/MOE8r9IarOcl
JYf28ZdzvJApvFCK3Wo8OtdrmatxCngnyxnn9taaFqNUrwhLSvjUYIeZp5VkOXoFdcnrv0hmkTxl
OOhwzp0Q8ysEppy2C3UfpN2UmUYtiN7P2TOdiLRBXYVfmRlRkzfsfppDYJLbjQWyJp+nqwYjdA1w
NxDOPYx5Is1/JBtpNREFsOrc0YLHV2bte0iS8yW698UIjJKyqPepg5LYaKNiqWxUexN/y3O36cbL
StFAnxW4QLhiimOUTv0xcFATUzn3n5Z0J0S2yoeemgvzGD7f88EfiWI9mnadxY2EXV3Mj88r42qv
8IkKG7m5o3F1fwoDZac4o+k1BMcmbPa2B1iHvmKG/ucCQMyELu4V1nMgTzMBj7Sb6nNQFpyy4Cun
MYIvYuJzJD6rdK8AjggROTqAazOopt6cYzeRRzH6DTPsKaIPHekmk3pozf5KVXwUnTbphx7c0nqz
0bCZGpm5/ZmBWPddB3yBZei+9Ygp+LAmJNOSI6lPoZM1npB4gPd0N0nMNq/hJLKOQClO5mLka8Id
kpITYSAg56hZeV64ddQebeRKFIMLBXmaRcK9cd3SNAZ6VsFnCxegtGa5L1f0FKMh9ogG8jpfvell
kEGgnTdGvkDuJJCagSReTszu3IBKzlvQFx3qZl47OaaTJUisoeMl0rhZNv5X0z8jg3ED4Y2K7ohi
UvM66KRiqBxS07VylypLpksGNuAFgZKhOcsQ5+XcjIk/nhch4l/mDxljK+YrLdwedxMODRcQx5Ey
wJRtOsMUIDtUQf/z8X7M/kY/CB1o2WL6TSFU8fHrd/cbT9QfNDxWUZAs787e8V5DgM1yYbaQfcBZ
F4uQU1moySZaOVRYH8pMr0YcoJNckvKs0CMT4mQqQHEHUwIVYbRQTNmZWpzTxBy7goXHrkTHd/g7
6F36vN2dn30oTzBurOEcTb+uhf0zqLuoZsZv9VuwvXlc4MX4udZuGeTNJ2HQjz6cQa7UFW7/BRN2
RruI6qPFTVUxLlCyMbIIUkY8b5+RmTOvWbmkyRQCsJXAsJDSUuSvNboXDXxGAl5CBN1Wgv6WiU8v
rWUd261+yLeENV3NEls6SXLTD/HqxR+fTJv3eLeLMVQ+vZPEH/VgsXDYf70LzTNFwMnsQ9PiSocw
TZKt8bOeqC882cjxV1xMC3XbivZkPYWGRFlqDP2I4yvuTnKL+6kESmb4cpN9FYHdS0pTT+Ob4H5m
oraNebrD7B+IUgs/2YxyQwCqR6mYnun4hoGR6uTguVK9qSVcD01QjPS98MN3sUIOr+way8SYP41u
YSGoslTbH20OVMzaPY4ZUdzQM3DrhnroCahDWQTgcidata1xdAHBHgzoce+FIDlt7EhOYN8DN2gy
1JhOMfwgaTMtiFzNWlX/yXfj4nymF00fBI9T9eU/3pIYASnMbabhIYyUAXkhFQ4Vt9YMYP8EnIoL
8Zd5xy4mVOnynJmvsTINo5+Urn5+87XZRLcv0OiMVbj7Oytr7C9cKcKuGp0FoqsO1qQC9ip19ILy
WZ/FIw73cd7hjOgG9lbUoF3kgGugJXZzhrj8AepuO4URSFOdwc0WKxze1ADXnU3xAIOfmmAgJyrl
MJJPlq/HQAPOteo+9beZwvSoFj8COqMLLY6uTF9yfz6NoSrCox5QSPfGR3bexIFLJYNN5VhAUp3N
bYf0h5+hQD9OSNqwjCckUKUXCok/XF1KPyp3yktFByFZzrL9oJz76oVAnPkDPyBCucn97b82tTpo
xukOc+RuCPD92RUvGb+GDU9NmYdKjam05kFZHgKIrK4jqTJyktSMeFFkDRfWMV77GNl/F3Tr8f/F
Hj1hyZmfhDlyqgtzfI5fA9TFniILUHsTS8jkepdOz47zrgOoS+LP7QP5QeQaGmBrHC3l28oZ8ElB
SPSvYzeB5pjTCJt18bsoYPyNFyxUyhF5msEcU2a+ok9wtE8pHy+yNWIFobAcIJCmenPVDRztcpyy
bkBEtc8ntTPQ3X79qrVluTOiKbE3yc4vrl6WZrJ8DyZsQbrY8tjNbJTaydjqSUB6RtUEFg1B6UJp
fE218i6G6Lv0J9iyz/NPgBeawyxwiL/mfWJMKM7VgLOYSXD9axmBnLf52lWg8uQMqqbJ9A48Blhz
yFmMN0noXOWgdFjQ4GQOHdtNSlshMXu/8gGJ4bmiBnzqDde4SIyaeFuZ+jqzTnA4XoMtEJEWiapq
F7yFluWa1nY94vxhdGV1Utu6KWpoNTkrneLT3vP+CW7YTa9ywtu5jeseGwPjsSJPiPnEotTZFGJY
67G8ZWmXN9y2trSyP4xDPx9Acj1b7NRNG7cy2rcDp5EFFp9fHjRAt58/GF04gY0ORQDt1VcCChjs
GKYJRi9wYTe38XZR6dVR1YSmJIialg+/uSNyW0+t2c4eVuiG6+IfLdv6BQl75YzA6nz4DxqXbTHg
4bUkJDPKlCkwZFpB6cPcE+YgqnYjqviarQkIaAeevZi0GUWRAW67ox49wc9nsuEZuqF5NHu4/NSx
cjA3Xobge00JmiWbwJgpTAb8i190xTqgJxQE0Rv+9OkahT7qPBhH7EtPONQf1Knkwtaq8EVgU2P0
nmkUuNG1uHwsvgmd8LAiVCZ/ljOv+jYt5gl4QI/BcDrKPaCVM2xOJahUGn7S3N3E17S7AIehDhIO
eOsDu1y09Ld97cAPILJVHknFF//xvjEoooP1ct/2X2LWazP0s2EO2VgL/w+xN0HGxDGIdQyAbk7e
70fqBT93lY7OOuVKN0U+cR0cNKvMYJoMQtB1HJ3qhl4ROjrkLSsESGVVnIa2oyOaQvKZ+pTmTjyM
0c55jund1Y8+k+Eq8Uj9ludmudrpUa8KJ0Ty8KrrQs5PPBImHMipBDlBMK/N45BFnSlP/gs+YrvM
TR/W7dfutxtRKIjjcWJlqK8MQhfYIlWyxrfsO4F3rMxXXiv2HHOSGKB4HD4tYBKz43hC6to5vXIA
6XTnHajamKLivPFJ0yc6/Xzwmp5K7HBCB0jeNwxoSx85CJ0Lw0izmiUfeQfl3VnlWBred0q7ANHB
76YNxabMF/6fNVDyAHTM/dWgspJRlUPQTDX5dz3rkTv5blMHrty4zp9vIXr8yiAlTZYpiRXPs9Dj
WNHhTtgzv9m0YZSgKwIoDwFxaaeByKZf+gHu5pY+gY4nKz9gqBgqXFfSGqYIsNCwsR7zwgQxmWzs
AJeWf6+8SxpIej0n7HWZMwT6j5f2d8RAo0311b0cVZ3avgV832a9W+zbQ3TD3RX6VFC3e96fSBIS
V/XICphqskrSDwvF+jczkQ/0tloy/XEKrqE/IpnSgYIVU85TNYqUZD6qy985SiRrCtFwmb5/jhfU
r4yB/YVoF5RiQxtTRZC231qTbfdffhImhxsMQQ6jHyJFVToN/AmCcoEw+T6qAQHIkRKM+6/Dh4ij
Apepxn8CYOFpdLR46UkjLp8sNdyb3+P/RtpUx9C+2tQS0AZ+xrB3k6qnsvtR8onIbzJGpzHS0b03
1bYZmJlEMZcMdARcfMgvJuHriqv0KCODZvIwvkLJ7FSgq3mptChq717VsAyBCOFNGohwuaEaTVIk
STcJMWFxKDKIGxLLhJQ7PK9GMw/njJ5+FPv+Lj42PyiNM3wi4w0I3nSWraHMxcHoHrvnS7ckJKN9
hilT5gwsT9hI0VfVrYRYpsjk/pZKQt32ofhgmRayKdKB9KfVmPuSJivkOUxbhYFfTKa8XmDh4I3F
Tt/XcvyTCzKH4bWrAbUHSlRSb/qoWK5rlqij1+mSXTwMHrhbE1tWk1r/XmA9s4p/2MzHqCbVIysa
oQTF7jFhUtRgIRsBfkzLQO+69xFJvkf1Dmi9JvpBPymbNAY7N2vbWfiaTKCNqJuj9jZhJEAuQjZF
gieygW3fN4lhpmxskW7k52wfUxTJ6UU+zZ5LNTQFnQ5B0Hmqj3gO0nutm1mrgg4TcJV0RodDIg4Y
GBZx4WM/zZmIJhPPSltF09mjWr/2YkatkgPXs9zMrPVMxQ52F68KzbyVgB4d0OrEIPSFE+KNJnzh
DIqg5tEjB/6WWDorYjx6khBdBCxWz+h9UIYaiR8t6M67gjwler4sQdUqx3UP0EReA+7uL/4Ji8Mq
1zlunBA3XJClnjGxtGjxvjY2Yd232kMu2yPAljmZXNpBcKAbjeS4C/VE/shQ08bA+E8UQ/6pdFxz
nhdEEVZyPwLa2z8oXiF1wzyS7nYVS8UUgY+zFqiL0amfJ24LHAQSD4lQq8+lHmzOl2/Ed3RLmFlM
6Fg3Ub1flGxuqtvB3Ffp75GXcbjw2R4g2wPw4xdq2+K7BaKC/TN2oMH9mIUIubVADTt1t/VOAp5k
4ts63gipuPRPfyWMVdDfI6hx21wAMjuc5S+xp5OYRMY71YbxBaYB29PpI2rt1dP+e+qfXyOk55ga
gVSy/7iCsF/kPNe+grRCMcIcBg9vQaIa9Z/xWtiTlyv3CIeJSpx5xFYVu5P75P0z4P5doZQdmjwb
rbcLRFAivh0egDKoNKTUjw1+Z/F4mwZtgvW7SRHzXPI9hjlv1Xrv33abvuOLMbFQlfUzLqN0FdCW
QPkjD7dyllL2LbgM6DcSaNRcblDvQJtxe6EMb11dzYkvxADAKW9AKBBXK5ikJBRc9ExliSPpQ1T6
gkuwq2/uLM9JYHE5uC8/mLwioDF3aKSbOcMc495nG4aBSpVVE1NxfLVaK9YUHY0KTsUUjqTJTv4Q
K9XdirxSOEUy/DvXv7D8FrUMLm4G1P3Uq1MmlN9xnq98naOBuO7FcdtmkD75DP7WAdAw4D0YRxe4
NRbYcs5s4g9MnuNOpqWa2xPxQcqYNzOUKVIYp4xYHf8BtzOLsbESlbMQoF7HDGoNI8IUKidAGXnR
g3M7nsEoavtfP209cEPCfcfkvC/tmBqZCh77hswAOhNu6fE9OR5gzrwoV7zCa3/SvbEVzbS83kTe
e6TwbZSBlJOiqAtaK/g5mh9Ysrf/i1BFOZo+gwZ6C1SEY3CNucqpXxXwxj6dRTAtF6WX8no6OQkS
F5fkJvhsmlDlwP/9gdDpDPGFK1lmD96dmrwOrq1bykVuPao9NWB5EuoTPcXlf1kFGF/utI1Lveq2
LbgmXu6hQptTDw5R0lEoOC7E+31kui8/yEmuW6I72wU6hR/4xKPT+J4I+5hZIP/C5k9Tjk2sxhwh
r0q568t/npTd2hMq/RH7bxNP3K+oIO9YPCVwWbhtZNtOoXotNvNusANYKDu7eWH9fBj163G+jE+4
JWpIlpG2tIvRWvX/Cu5EbndFZyyBl7JTkk/s7YkSp3L87MIn3hxzRt5rjA6oYty17Rzc4XVp3+u5
+hWewEIweYPg29P7zNwzShv3mTx9r24G8aw3O5QeZO2/PO/LL9kbhP5YW9M5p8EjJqCLVOaYUYkn
gifWNNWu80060NtbEeyA5PODT0jdM9z+g/CELk5/mqSSG8+lr04RTRqkRFCjeED+TrEFbC1vdNol
+f2Y0TGabIGeqncx7zjjuYVn6/Rm/7CPUOB/eSp7lGjEv1MkS3TY/lxy122Cc+LuyM8hzH4TTOOs
rl+N3lD+3RJmJM9m2H7uRCFchKR3FhUNYng1nsoREibMY3pvMd0kgvsDAPee+YPWAfpHJ3ZAVPWr
6Ytw8o1fhWJfHFLCrzgfxnGDHoTjuDcuF4YLROb/fC+b761JcgKHymdZ/GtpR7Y46kvN3hzmUWZI
DRx0U6G2xplSXB9O+CQwRxNw62A7anmW7pTzIt90NP7l1QOxv/UjoDbVow7gWx/4wDM9TcchPfOE
xedu0uWCY+Vs87gtIC7xHzoTykOM+7Q1H51C2CnTrEigf2hANShNcn2wD528l4Rxcny1xNm9J/pu
5gL+L9iHJzUelDo2bnco/NLqL9K4lrOWWFdapPuZtKJ/re2IaNJ+KvCxAXXWUC4UemP0XMlLiNtB
LXxGCKZm0TpwIfQD+AZX/8sQ9kQ8Ojz2sVkm06TGJZZ9ZNjWr4b1TP4Zh/+1v+ERO2hCS9qf/kZ+
DJxT8WGASkhAmHJiuTueBERh4o6RrdfraIjKxxzbHYe4MPIK5BrPKNXR0yUDiUf9se2PrkZIKkyf
uWIAoamSGkOvr6qXMbqFmWDmiuBfw9xUheId/JUNHopkAEWJW8cHSLwWzTmOSgJf8yOD7CIcbtiA
8kBwdAFSHWp67VGtxI6Hi44SYaoot+WU4+yepZDZHvhYAO4L0Va3xBEuvex7yZ1URe7f4jQwkDFC
relijkATYsejSTclDmgXTwg7lKSJD9rouOV6ZV1z/ikCpCa5zFfxQaDiMKLmec3VnkWLUSyk7YpV
+RdxYncSU4JpNqwwOsnbCBy+ZgMGLa2U0m0KrG3ikR02Nmm64bv0gU9BF9L5Th30saev3Z6Wt1PL
OaxuV1OJmTBd3LD2A2q26ku8FDT6u+imcM5KTQZmZFzHTHQPrKHaitgZrmZsS4p+xnbaD3EVtzVe
i3s9T4UtCqgKd5yFMAMmz2xtkgUMNPiKe2Njos+dAEMDYkze6gT0NE0lc5+ci6LUEU9uhPNtdYtf
RsqPeX1+CFOEr0n6oCd5mIT5tA7K5lKGlLhQEL9dUhhVOE4YXGjg5Cm66StLuNzi2Gn8zotmpiYJ
FQwjU9Mc7m/sTq7IffaRMG/Q2pRcCg/wfUd7NtEoBrFjI+x+cl15zA8+6xb8qW2u6ctte74hzkcn
KeHK/43O6rMsGBwjyRjyGDOY1Co7e8m3ceASTA7W97fjRWoMC2YCPeAAUX85x8SSD7UbWliFZI1t
olaUo3uU5fk8RmnSqDJHwAZ1ij5j6zHouavPyTXS0VN1ApNjXyLAjv2jN2tbLzZT0av3Xl4dnpld
e3yaBukIANj2kGvIDppjpu+BBkUnslNuTEHJquZAlftQHm4MuPunL/M8+iuGt0ZuX0jBzjvzLyUl
j+1T3+7QGhYugwZ/o5A1xFaLr6LB1aYG/2CEOpT0/lXV+61xa/sWKx4PYEb179FYJH9vfmCl6GYP
lWqwlhqUn3UvEobc8AEKJCtYDGti3IgIWgftxXaBRcRI07w0w6OpfTfOhauwNXBaduNAUH6/oi08
768Yq4RVVv948XmP9vM9MPLL3oSsj9xTBqerJnhRJBuX4HEf90kJh/oSaDWw2opr0+xP3/Odm+z3
NxsXGBTPcdXLkgdQezuZCvrp+jrdAdBzroqPXEEENSfhEctdoyJ2hBSo8NWEwB8aDgPSwO0DFsEZ
AU5lO0ANsj3QjZHCsZCYI1MY8KP38tECWn6x4OBXyAvyRMbkk7svVOIqp27DYpGS9NUFBUy//WdZ
ihZCAZk3l3y1hTL63oAhReKlZAUzoBqliJ0PPKlYYNGPnIv3FXP6O1pmVOdYyS41dnA9rYSQFbjf
SAt9Ux3rY887X9eLNnpIT4g4Cmmei4tyfXWXiA/qEppJt8+eJuX/Ag07PGXh1E4NVcbF0pFXhhXg
hzMnEN/ScSq8tuLLMs0TqPslLZUGMGegzRMQh1UD2dF1SHecDbpREM6fns3TimdB7qx8OjJKsOOr
u+bqvnygcHWHyd8kZ5miQEDgeFvvL/qCLoQVLIFjIZKhwdG/nsb65QIXLkU/51YHIczBeF8EsYxo
x2I3dyktYwztGLPsq1UMyPHlovxb04atz1JdmIBZYBz6RJEe0YJL4i4PLQzBzn0mD/VAmgxMsWcV
NdUpMLYI7/2wpMrXnsgvQIG4d6KPZTTLKMNTPrjnP/wTFuZFfD+im7gl/KSgPko3LP1fsM2530vg
dMOmePgGRUQkDlXkPqqWE2xiTRXQLF2Lm3xEWazEgROd5huu9jmJfAeamMk0NbUy4o8ruQsvZunP
TIYKxyEm521OdRW0/9JwcHwJhjPT2qRp85wlgLd0mmOZXQ+T46MyqPsRNzkHJwuMzJL7paEK/aCO
urse4lZkZUMI4Jzm2eozEJACXcDaGGdupPT9L+9N2jnamrjtba7Pm3UZo61MDT50e1c883kP7c3/
vBR9Iz+ovULdDEA5hbVO09AHeJeenw7Gy50ldDwmjswD/DhXciC+6D9uy93B6V3l61+KJy0YO21a
6EgkljKzqTSNV2yET7G+aXniqjkz9P0J+fIjG62WDc+q6Zf6Kqs89diLzYYAS3W8/tZGKiE969uK
ImXns9F/I2VYMxIFP1koyVT+8aD73urRBmNm9HoM7gAuyLAGC3xDyhhAQyizftx2L0s9bipCMuHz
/gyfTtr1CUlJ6CeTI3eVVHxPNQOAmuf9VpTcL9bTGsx8FXgLAQHbUBg39KVz4gjiPRcP6slW0rMj
uF0TFXLSo4yFOyYq/ZFAtua4PN8rjp9L/wgJmVU9v5zzEpuUkY6vm3HNSaI1NYWapE1TUhIQ9bIR
48lu0haruM+RKTSZ68CkhYbyhrYMgM1KOoa/abEIT8T4lttx2ptLsbrKrnlr6S8xZ+uooGmHv+sY
tv3s+DcqHMwPwxBp+p8fwmyHzbZuEBwu0XVsrH0ztuDZrpOXcKRmGCQAPU3ls7kPc/2IpAzQ0C40
z1MZFcvB7pL4eyi61hY7GP91nqPTsrTsieK8MkQ4SQeBK3Ig20JGfu3GRk9k+mOaSIY9dwXkxewE
5Hiq5q8oV+423aMmQpnWKw29uZhonPmosmVD+VuPHhtdsHIofdxzJyJ6jbBeGafxb22XbOrG9Gm9
giOPnqG64S24VQGNhzMRwc/FweSqieUSWVLSWuXxKwea80KxKQDEPuz6pmz/kkJh9Eq2NrJDtSyc
KAYoobMyygJbV9MeX/d2E9J/YuDxdmkKXtFbFTZIEIngFPsSyEPEcyKkDqpdNBfMbRcd9eRxyPyW
/+gfZpO2mfGCndwj21K922LvSawZeIlTZ66gyQDuU4VgDNH7ymOC2b40ukjNYrsykbwyFyiBi9k0
FJQ0jsOB/3AdHtxhNDyPTd63LwMDhEeSFkNlIlE4HxYPjWUaq27TUEIxfksm6uh/hug1hfhY2md3
NZEXorKkdX6VtdyKqvbnJGThscZznK85IWSmaPW++wpxnyVf9Pf558Mcgn1JK+XUqYjisFq6PiiY
QmGx9PxaSgAHYz+HK6usZI4tbrFcOO78zyDseM1KBvBaj5rfEHcDDQ5kFoizds3AHwg0K+0FlBbH
JhgFd0PPQWZA2RTlQz7zIqRdMrk0r/65mA4H89mUjE5aovD1axpyPlvrHnr0ztJ6/vGX9lA4EK1l
a5qX3oMZIkXMGSoBla++VaT1ctPtUxF1QufGEdLrSaMU2VQEPLqWm/OvvqGiAkG0X5PyjnMSJ41X
qRIJu0Ci22bJmf17TSqiSgo5r5l+pqMY86egiawecUDdDquYJw1qlc7Qe/wZT9uYEpr5NLZL3Uol
gdAQ4OpytJm5vZ/S00zoeakEZcgu++9Ss4AqA36w6OdU9rYSvJ/7s9Eow9oC3OoEwdwc1taM6lQu
mi6J+bVA2aMKBy2JHvbQLD0qjJqWtFK47u5XqlA27nYCT6ibTNwHDXb4+x23AkD/k22+FyvGyoxL
g9gN8kfCBgYcb0LkPU1P0ZY9TEkce/kf2vnEoZhby9LaH+f2F2LHRvxr9y3d+7Npapbq/BA4Ja8Y
qVoXhAaHDoSLYq/5qYlTRfg8J+oSgw8hesaF9yYlS+ki86qQjbKAwYYZwMelnJPjUrYshV2enxEv
caz6mRTDBp0Qr02/44L1XkBLNIG7D4r/7wJiCu/tkZrmABMX+q2KSTg8Fp7rPkN8prExZUKjcR66
0p5ib4yOp/+yZhDEL5o1GI3JeiYfxmj6FuqSBmO6jsxHkn/INjXxL2MqkbNACCcSg2KpmB7khyX0
2COOYz9vvL0+pgQl2Y78fz1JQuMsScp4kFDVw5ZMCs+CF8b7ed1fST3Dgu7ZEq2ySoWqONchJIXj
15TVqq1rYZ58Ox5Ez4BS1FaB5eXDTeqHP08/7BXX+Nj9ND9TL7imaxiwsaJCXYE416qhscVy5tCE
ZnZn/X+PVsuUhjOASVVv5IKg4oFbjX0f1nHmlrZOL9ofTFbs0IDXJu1oucaajvRuhPRY7G/BvfRy
P9By9Esa2B7p5xFM94lGXf6n6fUvE9XwK+di0aBR0+HHUnC/k+t/VmRuCFiL5vMZWHqkH4aQlHmt
OYaZa+keBLLswfBI1SbN34b/VdCQv3xdKwWAbX5RCglAwVzVSWR3LmTqxIpXVNgYQYelNUenvyQX
StXOPwZyQJtSuDr3zl6NCk4b4uUAbglOvfnndNSfNS2hp5p3cwlGF3+JJTab4bMXkeXX8BdsoUCr
592uewPgAWs4JklDhrqpjN3C+bO7zyGpxw+t5EoSVt34oPKuCo5PS4z2m9Out7A6wS9dtOs/ClAW
jSUSrnNVCFlvu4WTP40n3yAxS2Yjmz/imPnCI0XK10AIzJQMZMrYdjuyecgb1Wd9fY4zahwf4Tc+
UWQBWgTM81rETaToNuIKvh45CYZYhluj+YbWr5KmKFZbqhIcM5dwyq/hoGXvM8LpL4dyZMS6LQSr
uGJ292xVYDC/j0TYUHm0+g6Jkb34I93S5E8frZughF23rUSKloLExsvURAwIwwhp+p86VhbDbghn
jo9sSqHMEhOhO8/I3lz1AxFlEzlNxZWWFZwJaKNUuLK9qibfLjY87bS8eKsz6o6iWyQCmZMWIZYg
ivmExlOdUFcAsQWymhLxYgpE4haBTuAH1a8NNvUAG6ghSLsxcFTFGm38lAO+CoJe2EZZeC9IZ8P0
vA1Xpx1ykgus/cZr95mxvx5Ym9AKp7bfHySnY744j/71b06+wMFUw6gQbWaebJ7hpAg35oLvnMyu
cWJBbDcd5Cj5EqPftC/4Hb4cIU6f3yRRk/cwUlae9DNWmXp6LAPOlNERF7JkWJyJaEjlmQAHNjEI
ETUAVmK7ayIBI0ROUW77wtqEu+ecpgmTSMpQqUs60+EwqTqO3l2iTD4joEuc1VH7FXcCzR6wFTtR
sN9fuATnUP7jW3YLN3tFuU38lg38h7lCFHY4AD3Taf3C+7/NyEd4ycirbL/FxFhItGxq9zG1GUA5
Auqa8FIRjthCVgwIAiG1sTIfwQfLn44ZBPxa0n5bowC52v9MDE+iEZb/LVGyQlegMk/me6aM5wJc
B3+JUuSMudKW6hO08Svfu7dCsh759f+L+tuZqkK3aaZDZkg64W9CYpF4AMMas64GcYauZYgH2tOy
KVlmQCP2MifNdXf9KBlKkL/IbMNLJBEFusq+GK9Faqyp0PPkZIeusZvyHulZiV4qkl5M6p9Lkzzd
MN+MAuTz/Q0LDjyqS5YbyMIiyJ6h3Qkf1LbKEPixYmWBqBCTwS7HZ0MlgDHyXA6uGL5tP0vBGsZ/
7FJjlLjuiVvrqtn5FzQnz98r75TsFo9Qs0cymbJrMB7vpOwAhwIs7T5sct/GuSzG4kE+o172PJnI
73bZkkbKVn6YJ0wBeEMC+fhl/B8nu/us7jrr9zzFw2QyDtF1RIOA6TbOWgYMH9S6x9dSiqOSrKZS
NtoJ9mi955EFOMZGfoxAAkTEgMWGmuQVVnv+hREL+IOtwdbS7yAnu9VAXsbAlppE6ZzQLv/qfLXX
WTYrXkqz/M9I37OhF05q1mfgydJYdmKEAHeGAqN2oDAiWZbNV3H/ajiNjA6PHupgn6dN7NQsqit+
L6yIJS5S8ZVvYtgj5OA6SgmKnove5CAg3gA/1lS20alMcekI2eoL6MU1+IeBk1aZk/3YAoJjhcKB
i9rAr8f2QpysIWflJKOu2JcKCt3nsfCXK7pgyCuOud0hupuGW8tmUmcx5UOi8lSGmr4d4sAWP6nP
VEnIPVZrE4O76I6ezdAL/ZF7SmsGVQrlbNEv5WFeos+d+3+qK0cwedaS1amMuqmS7WPsrX/+Y6Jy
9TbOC5bwhRJ590zvW/gXvaEeoOunzQPMa52kfZBzpsdsEuCfJqRrZc9O3FPtZiHWEuc3DOw66a3c
UjRwWUHWKgiP8sLoOO7WkecGOSFjeWfr532r1eEvY70suuAW4O2lJ+hJqwZijs6ThtwaADxZZh1r
Z01HrCQJNwbid5LYVH97UQiMYSsui3wrVAsKX8lVyJFYrltYYYhmRUYhnNns2HV+4U8al9DHyHow
uMh2rIGOdChjyoD+3gqK2qq8Qzb3wXX4tolI2s2R7vPboromQN6pGDC4Tc8dXiES5e5S9UCZYEDR
RpivrTQ0kdEbVnyxq0qQcpnO7yhPWYx2DRd6IapP1Nb1wOl8RP8SQsYQmn0kBXtubGB/B1VDSyeJ
u0S7gkiAh5yma/8+xp8B3FaejXXIRGO1Rfjq+IZBy4NXQ6k5cglh9DMnJ2ZAAp/c8UA/dYhtQOLa
tTEou6RwGShKAg6cojOn6xOyOuaeVpfmAGU=
`protect end_protected
