`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xzu3iNMxcYwWeGE7zBBSQYEQ/PVQp0Qc1wcsI6um0warEjZWkI/USQQ92OzWQVkESiLoJTTmvxIi6SnxATpK1A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jRjdEgkXYK8VYoAf8QP+gWpohLZwa4QF3Z+xEhWa7JtJHPPyitr63XbI4BA2S1gieeBT+7Xj2YKw/QIeDWh0/9IAAKtXGp8MhxDiJLiNO+Dq55TPPj3xBbD1zcnaiGxMA6uO8rRtCpUAhhEoCCAZc5XoEMYzBE0dtfexZkGdKrI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
2K3cKS2CdGXXm2Zwv3MYZ7DGVg8qiSxXPh6oU41wWj1xHznLr6N7fuu0kvOF5Ydeyl36zQQpTQRyPXtTkq0LtOGwq2SfF8qseW+YLJx/rlcGy+w5jUMtCqNSBT8egyYNkIY1Yo60k908QyMwyCl2zxsZQgD5dbZwU5fbC/ZPyBwcGLWQNThT1J9BL455hs/UTqXrEyvB10EY9FaeS91b7IJItT+0B+r+bF+zUpu5UzMve+c4HlWMEXY73EdFdhc3R2v+2t+mZ5J2/DkRJ7TbcWLV9jw7fIRg6yLDtoHq8SV3EhWrlR2DWzr1sirlz3MGmEu1QIZSk0g0aNWFannj7Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DEq5F2evb7FcxAdhPW3tkZ6yQcQkvnkHnqUzthAlI1spohk3yB/bKt0RCLhRRi+Et2XfTv06PprGov524IvGZvJNL+NjinUBHSPr9bx5IyjSSrm6Oc6P2rhPzXgoMUh+siW3jRcEd4RQgAiFxMo5PH69LFH+SsqjQmK99j2UBV4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I9FSPm0HNafdO7snEEvGRdh10jbv+IA3Afl3FQLgxK9fFdfn3OnpMiK0ykaeF0OtRk3bzfpYDmO+cqjYtTaIbVAczAtgCuMdjLuprDl8+tGw0hMX9jqS88ndb5XYEV0gv6Ev1d4nOUOzbJAngBiVa8ums3xiqeVV42yeMlzojh1eNTuOVg94JRh3oOjpxqn07eT9Ywknc/xq6C3ah2qf1EmnJuOdnIuATjPcChLLTnKO+JG48N0PWqyJB0qwkfj8p2O2GsiQpMs7XET2hXrwDOXAO7bM+UKz/9fyr/vzNOa5pF4uDLoledBL8R495/PcK6nT2nCmS9FsiISM80ITag==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20298)
`protect data_block
AVHscbdBBvSEXtrttH2dXZIm2phkn+6bPxTp4wqpG2nRQJqOaz5IVSJrlxQh1NwTO5u3+qBaaHu1
2oJxMNjedEVwJOchVieJa11e6pQ2zruubf2Ra6YXHr7h/X+q6/3UmjBC81cskROJ8k8svHnlFNnr
W/leeaSANjZHob7ox9VI8d+a6GFAIrOv25lBN1AlKiIn9J90OSoqPiFoxQd5Cil33gAge6P8xCam
56e0KjtPnNAl+BgPclVwkML+7+ybDosq1fHfbhsOULigid6hzHLlswTrksSYKPmgBCXU2uIOM6Hv
f8Gm8UHlaEDANZVnm1GPvpfXn5WsgoRIUBOSJ+5dfsP2sCwGh6rNTGidVuUPkCqcbWEZl6srkEU6
gadJmM2Un3puU6C6WDNItWM7/1V1wKDQ4AU5CCO2QQ4ANmIdY/JXf6K8dqebepNziebMdEztEpAP
Uh6G+4XNROSwakJH9aX5R7YKsfFulfHk5my9aszl0JaZIgJps8rTmNW8esjhYi6ovwzvOQLhprx/
vbXKwtbyK22IuRHtq1Atib38aonB0Aij0QTAsskNJEAEgOPG/5bHf8BEAbLFEW3sdpmaTTqnNTaY
QOVLGoGP7SotFQWDQsxKV9xL6EEYqCg7eS9cS68FmknWBhWKXDTnHFvp4aanoJFmw7VLWmFts8H7
tLUofgXo6/nIPHYIfF/8j+ZHfDMMpPQFdRXgGXhG9IGYpCoGR86jH0JrPXIK49X7Z2uEIoMg14cq
2unIDk3GG+OXFIJWDgWxN4qWM6TLi3NPoL/xABjnmneKpT9Bb5bezakD3z1rchTb1IlzlrCcJcX+
C7KVMonoxHsDo2mKYFbvqguObBLtiJnUNqcntfYVbw5svvJNZ2EvDiOqKC91W12bMgTY+nqR1DsN
ZF7dCoJBMpLn6xl85RCu5kdWnvujfbLT8kAkF/X2QL7ejrEIWEbxwG0qQn57Q0Li9NehrQ6VyJjJ
guYeCNoF2blFe0VwIaVNQTUR4lsbPFtuu+N1mCIt64TPY4PUFlDQICyEQdweOIZ9yHT2paarOU7V
qMwQB8gG0ucnEUDHjNjMEqU1/zx6rYXNg68CHyKBAtMMKsrakM61Dzw6DoBOcw1Eg3ghJ7/KWKQ3
ceIjXcEqYc9DpKmlE6tTpw32c1y1LOW8CLX30Zg7WfIKjq6t+SEk8O9qHE/VDcG2z8s7S/NmJz5K
nH1ey85+MojX6AZ/BZrZXD+NkfWyKLYXRCvlv15DNK7ov2i83pGGjIE95d1yu9zmwqST4vafXuVF
meMsyYiqCiHfr087bEpzTdibDZ08lfeCXguefWOx1ZKAoV120GLwkYDrTAnRkar6szHR7c44rUhJ
69bhhozxkvD/hVS3nvRKnNM+EM8mDj4rGhphFClletswMLvj939xQxRiStXatd/XV/iOZZ8TqpZD
TsQ1J1Gu50XcO4YBAvdoiEQqfaqoHB124qUT9jcw6FURyuh03JgPBBDoMrOQF6LzooFoV6igsgUn
MJJ7XOtbUig0sSOfUCN5tT4ASnGxeXKasKwkBXgQaiGKnZbeSIr2RX1CNTKqIKMUQmZsGF2dG+BO
44HA26ANZmqnQxxnkIJo2FXtJgNk5RDi7GaiYQj83B+zyZTqi6uP2SG/oxOugpFIIs8rGsc23cRW
QrVluBgNnSnhuRp+5rLTb5N5mNP7ri7Fvv6jAHrmIMlQMQ3JLpGgOQtjcHpcJnrHnUupZ2OENUcK
eSAd0HK1A6dB+GGmy3YdIn/JBKCQgiep4EbohHZALR17QWqXDuDydPfWuUxx5gwPZxfgn1WoHNmJ
RjOXHLNvM0iLUd7XA7OIG5gHycw2TfOSuCV+k2RQjDIM6zJLaTBsbWOVNj4x+uRnRkjcfffKGskg
I8Na7j9/ruqUIel/5rY0nt2NXpjfXmCOhbLs0uazVXnKAWkBkjk84U/UgUKO68kvqRCTe9A4DP0p
OKHgrnNdX8ulLGQX+/BusRC2AelgpO4305B0iygd6YZBasRvPI61idDl2VoH1AkGZkJSXbQvQAke
rbm++JNZ4lkvUptLF2ydeUYRz24DsWgtzj9AZ161WSvG0yFMVXQuXd6tDUkT9viQpC0RHTUMe9e0
/GTZ12mKEIdnUFujy+A0UtXT5Y4U+a3BbGoK+Z/RyW6aCoPEp2QHGSc+emQoNdyZxLORcDHvD0W8
06L9ug0vgNpWIT3PA0SL4gUot6aVoRcta4OfgBtza/v1OhjAxdgdamy/02OXmSfHm8pLmm91t7aq
2shRux/AvEBaJmlQFsGouAZJA4nQIo0M/J7Tpb9x9qJHgEDAElkTBQh3UFVmFTnR2jyxY4wAO9eC
BdqnTC/dIPEHUA9dzWouHwVKZszmrJVpliJwnm6Shvn6v6qP698ov9KuP13WUL0Z6mt95J6A0W7r
C8MBkpi8WkIJOPpIzK3ayRCXmphqpiOI514qYOt7aZ8YrcUWH7hNxKOjC1p9hT3wm4svMnRbvqyx
ZiGe9kGPn3OtLrUlhFU0gZAFtI6VCEv19LCvyaG4/DuBu96/Hknu2+vcGiLBtQGpmGjuTcSxE0iJ
a1or1PLYDu2hNRYnnU4JfQELbI68PbsUeCcCo9RuDsEispRfpfVlb4THNDCpsmRt3FPO4Az98HBZ
G17Nzw9kKNQpesVDugELVMNRnsVV9K7IA3Lu5lWrg6DNO3bhOkIsdD99rQskXxsSd7aRKer1oR/m
YvPr0uUAp8anctMbEOBhH+iyQufjNtGaDcCG7eLLS1wMjxx+NeaKTDjuKKabSqu2Pj0g/g4GAmLc
ykGMjiEJ8DcwtrQvLe1cpA14i+6190BobF1n0MTx8Seebe6KGzqmInpH3wxAk6DHpI3C85n2X1B3
REbNN1hgWu2XeJEZpYOOo9IuuVTWtwp7fn5Vle46Vd6EVYojicqo0kY4bIvwzYSuF25tpVD/sznd
qDW+0J5B1BtetiF6Kt1Ek8CNIiflTJ9e5Hs64nx2AcN58iD3n+FcXSeOJHoyZn94Rt+uvNdwKcqf
ag4MgaXZzWYUZI/I0NtQZjFjIGsyWDsT+ds5Y2IV3qFn/HjEGTL0YBtB9kLTIw9K5KVPPVSnn13T
vRv1d7T4FqttR6tDNZOx/fPOOMwH6kXxD03M+rtkhNwFbaljY7maSFsHYAvFX+IoDTJgi5N/SrCn
SkMDfm3adYrhadpSJmUNGb6jHzWB0Z2pZn8f1e/E/pYHqdAFCkEAgEdHCS1fUaYWFJ9syUgxNQ+g
/lSFNBsRg2ay8BqbiZVv2NaLyFFekDwJJZUoFfRLYG0gWTWkiCePDIdCgZUqwW8J36BAXfTEu0dZ
L4e8sDRT1oR+LLoRUhwGxEvTFwxjApJlOVhfttcwytSiWYZlxcGWGvMkjlN7ktyGy3VLFyGtkiAX
J2N4xWAGzLEMrclUGLB9R9CLaddUsNFdaUQtiK2/VYZTwNkH+GJ2qphiHtUVEwlowES/nwMolxaL
pddsabPYj4JRBr6ukiTnbY1/HrTM+QHXw6lI3ShFVgdXmB6ISMGJeqyEIvZDrNCdywc0/U19dQOS
z4Ph3jMekii+i9JcLqPJ+BIdT5BNF/4WpYpL1GfzhI+WEcBR7DiL6eM3LAa7oXoZPHRZdDYHuDLY
Fa7r0Y7pAwObSafYMhopFXzEGOozDoPL4TDZfYYG79lN/7nZn481eBSG97CgyguoJYxJQtvTUTcY
mogi3tobn2C0a6slQScHUVzxV7rYClAlO9E8vanCl0P1mpb7cqey73+Hx9euvCQsgWZYsk3COWb2
sCl0FfpqXvfv3jTpIzOYOOOQtxLX1PZobTl5uXhln2C88ktTo8Exbj4w6c9+ydB3+CNWZWq4GzSJ
SgnQJuhXlPp/iOSHV59HzhZlKdvnjKSbLhBaubur4Qeymwb3ZKbmKXXKras2YQXwj5S2BRR3w294
1REurL8kmUdO/f5WfcF5SCnSuwPODps8iCW/5rZHEGO/lBuCR9Vls6hVQ9NqXZMaubh/bYNhDKfg
44HdfKl/uRTnZqJdO4HVA2Qp/5up3iM6fwwRnZrc2SwCW6v3V/ZOzCW0qbpIK+prGUWp6n4X9s56
/233UiSOd4zv0sW97SNBPKYbqjGsWzqb+FWsdSzFw/wvyX5c4d/k3hcSi66Pg0e2Igj7yKVh7g+m
EjUEiW5jTAiFf/TBoSDjIqNZ8w5M7qTg6eX7/NOff/W7+XA+QAlxn28NsTBUkClrirIzQ9CScXtZ
i9zLYhPBjfrtpd/xapEz0Y+lgrNCRTtucL8C2c7h0l68mYBbZ7+MVkU6VZsoTFVvL8OqshxYx+qn
ahWbjEPFHWSukE29zaKa33gRH+WGEkNygQgKndk1w1yxgInnvmougDQVCv6RjvaqfucLs/n39+VU
m1tvjhgV3Cc9nHegFlXQ0EqIgfWeL3aeBfcB0Hq0yaMQ2iTY5Zuv/+NAwWfA+NOVf89PFrXOb46n
yZr3LL3c2iVNYHcp+CvEOm930qs8nDjGWFDSfqDCzTFafha06FZumDUFUFQwtA6vlLBJZ0Vz6xIv
ubum3waGmEOU0vXXtT9HGRamSRCo/PhjF8KrobbkZT3SUZgaHB+TjKBKwn9oKMnaft4mppzwXMGA
cfL7Ss/l04cNwUaVC4NKDF4PsNWk8KELemH683ZRkLSSPT6Jih0Od4n8d4dlJHCSoxyOn52TLfDy
z5+bpJaixe1BNtq9spJluASzWfPClw4gcr8ZrRPx+bdJ72+pyH9G/QDYyiGOtUYkKI3Izx6M470S
Zgi/plTr0gb62hluKdrXkyCvmQ2tCr1c6XQ78+Npjl6f1J0Zr1LJtqWSClUC3yZ8Jlzn3S7+cLZh
BIgKDJ/NvhLqLw99kjjwa+XThpvJ4yvr689b4bvJUOId580Owvsg78dvpwUAUGKc899Ux/EBGraK
mgmQV/DW6OoOGGdpe1yg4ae0mrRJ4I4KeYSxpfu7sTu/rSkZVNk7n4O/AzvkjizTUhGYjFSDCbqd
mcw3k7vNKBXNQaIeHw8GIxzotZayA7+v895ERHEdJnpVveuAArSwrOO05dpBG2O/iJyBMscsBAmA
vO/1NZwy+n3pCTyzqhUncZ9VvWunCKlzuvXKhHVNHg8Xn6FsTkMDqxgis5LGycqaUquaQtv++PNr
/bTSABBmxg8QmYotLQK2wH3NKhvnQoIclCBa9wqL8QBIflqAKB4pM4r/t+Cna/qEWo03jT8ykQ6w
vWnH17kWeYJKBt8/fHf2qQW5d4+bvSKg9VF5F+Wrj4otLecLlLhFp9q0oia58o0XcsoATMwFJ8uw
JSCkTz4vxmP9ncBLH3LDO3YLREv7Ci0/RtH594g3M3tMuNTGbfzdI3gEqve56vQTDZZUpdK6cPYx
FOqSSsFJOC7izfpCiAVySyVGbKqzISe+0SG/p+D294N0lrkxLDxLifuHouOLkQA5V9+nvM8FSIrL
5r5z7EqYaR0CsKwn4h2qSj9ICQWH6aUQlkqDXeDJSHsP8BMlG40kKc3ivr6C30HfQyo8gulwUnvJ
P/6M42DCJvyRfQ9soVlwyRtj90uuPjRTezQe1cGFdnVmdQ7MdHFylED4RUHiKYB6JNmQ/Ddj0o7b
/SywdT52ssPtv10vGz4SmBvNX6smwbUnb+tirnXGIOEU/oFcMfZLyuUHo5csieAryrPe8+NtaleB
HZf/jsKduODzSudodT5+wH601SWmSHAy4z6BVDseir33fyfkBuCitr45tBlIHIvVB0oBkaoY8kSb
+yQ6nMre29NNRrS+qVHcob4Ls0ueFZIiK5Qtl4yXcELMYLA85caaayXuwOai+zOjZew4RmxZzCCQ
pIx2ao/+PFgUOH8LftBcf2q/j6slsYWRuZl30IWBg1W2PxTnTVH0XTZ9FdueDtkOheH1kaTRyKOx
hsb9cQ2mjnqhGYBJPFLvUpEGyN4SRUuugynkJkFeXQz08zUwU+WGuCpKtm+jJ/q42byyYc50zo+G
LIf1E6g1PVeubEvDsQHYSJimpzD0GM+QE02gbT490WUnYqmRac8F8xLx8qKmBEpECXH8Pr3UkVtc
6iN2P/kseRbrjmOu0RkTt3VWgYucQRs2t8UYGBggaFJhij6cE8ccjaKLLkfnzbgLRU//1xTgrEtr
M02/enU1uSR3TjJjGAE8IxaJfrN1dW7gzdpEg2evW69HOmwrhnXjLolUmxaq4K/ZBUuNkj/RszDy
ety2Zr9Vz2ODNfRsh8OdU6mWZUR41zb/GdyELxmfgCc1QUPZB0NMYSDO01EKyDI7KE0OsCOF97Ba
X5n5P91xX7Fgj9qNjmzpcUziH9XRcL6bSVDngyErpxXe3zb9bpX8CypgtkrNk4+qdo2mne0P2Hr7
IVdvEibPtbvlDbRXQUu2+XGsjWB1w8iFuXTZ4eBcBH9NGjnpGlEQ790wEQX+0xHl2LDw3RwpcAhW
k0M1+rfXPgty/vKXRzBjc81TywYzDvGR0J0oEZXcvwaG3/TFrNsZA2j+/Fa/G1T33AEvYGiqNSR0
9ofzWSW+mu+7629kJIWo5qJTDtZoXpOCbgDlBWSEEB3M6m0qbXGM87SoKAm5zGbLW2wHejZT/Sa7
Vl6nvDLlnYmJn5v9cOeEh0ZrIoLROnu+GCMiO4XqG/eWmEKOtOdb2hwOQwozRTbURbJngZnmPdGb
ywSJZPxunQfSDLumkSoNBlL6HaoBkLeP2SUC+1nZ29e5hkk1qoidDs3wESJfnH1bgEnN3PuOyxde
9DcrmlROUt0OtayQQ0yUpKM8q5TloFDGwVS3oz3PyJLFUihYPnvGkWDlyA40whADG1TY4PC5l7fh
2M6TOHhJ77UCT77JcS3pH2wktY1aUu7Pz18etyXLR3FFDJd9DfqCCpdKqUgtcYFLcMsjsaNkDpEc
7jaQflmjQM+hDayXGtA6rVotUliED/3H/KNKOpXE2h2ZPDleCoqlW+ElXLIWoZdbfPxUDFTCkX9P
UVy1kkF/gWEsllXLYrr9uCAwHjpASi6f9aIIuWfcB8UYmsV8fXVYdIm09QJb7YMGZ7AOCLObyMZU
E1XQWNB4f9KJ16QE7/D6b2K7AaaP9O0KmMPvEFXJUTezEzV5zoBcTrza7TIvP3pae7Rl/p1Eu/xA
bJdAGOrc5EQanJdZKZ5FXI3kBxXE23LO+sE66sAlqZ90apxzNU9Ou71KmFN6bDo92So3WCI1gdaL
zluG15mdHTd9K8Izl2erLq5A6cGbRY1flvweK2zg+n+woSWWu1jtwehJ0crt6N4FsKYcPdlfhs61
noGRL6NsSSmWWWBVuZ0ELH+7eywY3Vr0yEHf/RVod2ANva4a6MlYJ7RzqzOfChXdihU31/qRZixk
QUHNBRtInuuXftkn+FQXamkR3Zjr9bKYx0tnkPTrW15rKjwmWR17agrMD09LKPaiAnWjCFm72thy
LPM8OJNbkLXs27AJzv2zT7l4fx4ugLifEHJaToRxOJLmcdU1QxND0MIY6eTU3yudGalrXZo0CrQ3
YgJM4fGYsIfrKimFPzNT0ZdLe7QcLJCbPEY5nuTeEvsI8SulZdQvsBcBrXU5YiUDJ/YUdohQ2BFh
BdgGhLUUyzP2qwnruofm8ieMroEis0d71KqPproqB40evyqSHabbmYbJaXc9Sx8omVXRpqhRHb0x
XRhdmhgsL6AbUIDmMq87MTWfBkf+tU21z6K4VWTPWyw3VQYi21JG+EiRZqbrDunh+3fIgiA+zq5A
mhpV7ntOeLyDWoSRj7Ha8ebSS+6jjyhrqhQFms2M19xXqf+47cQQXCH6zhnVzTxLXLhgBR2Z+yxn
fUZdcBydeGL75yQ4guLCLG3LO5wBrZ+DgiEaCfJt/8Xc8j6G5JGbXnvCzBPjUaqUxWlFrsxP9I67
OIedQZv3ZeFUFUg8dbkHCLJKl+P5I2yoOsgzb64Nu1crvLTKhrD3dDVkusskPrqopj0gJk4Bzmr5
S9gzRE2kcA9WOknsX4Tib7v3CaHGYszdqXxtxPHA3eVwHWeSdko+oeH67t27mfALhfEc/j9ryW8O
PzPrAoS5lZZ+wPzh1ZpoOon+H1brs2Lr4Ms966l9f0kuqdBVhcNKHAIa3dOBiNyodFssbIfDNHbq
alaQ6DEtpdmLUTzpNpMNTWhV96OoIAwau3u93f/23lwIYiyYEXZ610LfxN4dIRdKYnHaVhcI93Vs
XYXz+0ZFbe97SsZChdPN6o0s+TUVKG0zIOrhWxImG2A3W8pRbY3C1QuawoAwYKkrma8ToCoC0Vyf
RBE0pGrhr8XCk87dxIoWsE56bbJIij6XTsQaR8pp3oC5fs6o4XESseMfv25oAt2XvMrMuGqlGLOO
BHkxJBC/lpTo5JEuQekIhkMiZ6xZUKsNmHilB9N0TCVylne1iHjjuvtFuJDeJfIqxmxUOM24oE8x
u95U9BlET2TIlmvzRrrorYh1+9yrDjj5sU5a1a/ZAKeaOzFP4/kdGpF/CToJZjhRzbaMSaZYFuXH
t+fuq5lI1KM6n5n0ZU/qNUBJHnwPamhhy4dnlN2sKLoGxidBqtUrCFAgYECCpRwVIeN9ZjPZ6x8I
eLlpE9Ma9OzAnjkrMeoxkwS1Wia2RVSMapGwe4Uk7cml22e0/z6W2TLjOYvDxHMFLL0vHxzBN7rG
LNmUTDAbtIxSTy+IxUgko0PUENA150dWGcZWb2YksiytVJ3QbR6uRSqzOe/CM0bfoT/TXYylSZsb
YchYYZLdm2wti6NrXeBOEFVClpB8bM2Dl5StFVZ/s7UFiLB3YNjW2JgMpFZWbICak4OX77c8r3q4
yRSiOFbnocLY5mLHADTcBJAXIDa9+FoOCLM3xMT2Wb+4LfH0JE/UmurFuwFwNRxtpOHNeVcWRHM4
JE3kGgetTFgeOPfRvorhPP1F0yyQIsxrPVIVxTFhDYIij3KXxeFRomzMzoTSyDN38P+80SiZo4CZ
8gYzQDZkmQckKOwBgVs8RYoPWuKVuo7uB07X/3oy+cpScqtgGqDq8ZlSAE5PulFGk9YTOYryLEQl
avL4JzEvqOmetDjlxXi0nkWYsmEyJQYBMY29AqTp4jXy7DPms5Fx7WI0O0KHIXozZLN0GSgWOIUM
nZHwmb3DAeItrjWF3pZGovchVzbAXBtQ/GLgJ0Vu/OFsuuRbBNGIzRmFTMIOQECJ+ZEqJlUiTfMT
/wsSjEmkA/d3D5/h/3eqfpLeTiAL8+9uZSGLptNSRNOcXhQ+6rL1E+/TtOkUseLn/MOyZpx+qc6G
As8PH+koRm3P3iGRvQAAptdGgy2NawKomPp1YWDatrozOMb6ZC5Di4DxcvU+QHWw7PqnUDFc3Z+2
byRqWwYyMBvo3UDs+6Bks83tHbn2kkKi5443K/Nxy6E2cts8focklBIJ1F/pvaxtA8iscVxcy4hh
ZBjZipiir19U3qecabsGwyShwd/iZwkJWpwV2vlGOESpVmU4FgLkpPY9acQCFDPe7vRyGqS0/SU9
U98W0w/Nu4wF17cRMfzE2XARustBPyapDQ7lgDNHVLW39LHCp3YyUxz4eQqTaogKaM3CS5yc2W+u
tR7laqk8fKVtlopNq+Pi5tT222agm5D2Dwf41LHADcskvELyXlflcmRt4AxmR4EbiLcN/LbFwqQo
3LeoDPZx5ci1ADu0SX7VYpva+euHvsxk/ucly2q8pMkpPclf0aAuYgEGzaf6RmS8PPTLobDFhuKT
8ZlelIcHVUAxU0hrcnRb4q/IBNk9SLdRRjhKstlltok8o6ON/E2Fx+Pd7Uw6CHXrubV6K/f72f8d
SduWfLzGM3TL95zxWmmmEPk/zCSufHQgMyJE0jIZ/nqzHMJuN8Uzr3RyosFiwhgWpfWyxNJZN6ed
4Axue+2p+QUfChvwmB7MDtcfGwCp3wyIJhCVU3XKRrvTK1UStv3bTm/kZiizdtrMPdt6S5N9zExZ
KX94BaHGYS7VRCDRa6v2VhMRuZ98MkScHj6QW0FDgAONCr217cyDu3ovstAfPpO6MrLh2ASPuedr
7GE7pX9LspXWRzyJ2fpkGuxAwmFY4gCyO1vOFZtysIMUCdCs3mHajfnUgzW1wRX7N+gF1NyEW+N+
7WZ8RdUU/80t8ocHO3i36P2fKYQx6IAitxaY4VTYlcGxV12cEJW8/ZGeVr7AEI0MSmHUBgRb0Enb
nh3xHEuYnC2Pe0VFN5VAGFz+BCLecAW3dWdVEPEpS1mwFWK1qneU69HJMQPBAwBhpMf7K5EcpU6q
XltYAY0OezbKe4ZA5KQwHzOYQN32h9hOCNzPxwzajZ6mxb5sUTtV+V26sy1dJdXMOqulStBv+H5a
jCMLh9rxsb6vaIek1tK3qkybD43oRFTNFHmevTYm37vp9rBZO6PaOFwRcEZWjsKDBOtG9CdrIXwT
AHLEhJk33h0Be1XLEKp2F69Yt95Qj7lcwsm/CMkgDyQq2vNxieOc3Zrq3qI1qSus2V0yjQhSjTP8
f362Mns5NZAYO4khMpQoqUCfi9nZhhXtn1zYZfCW7DOujvt5NWWUsOnrw5h7FhvQUJGt88IsU+DV
t7OJ0XDxVjDgLMinxB6DereV9b4TteSGBP+okevmlX7bJAM8huwsW6I/gHH0tFb3jnSx0TULszva
nJHiY/9v5pXXLn/iQJUyhYIv/IApyjEdy9bE42NPIA133rriw4k1L8/Ju3wLV/7ZuzJ3dXSpNQOV
sNZg3kiYI3gSqFP8v6vEVKLXxbSpPNHWefhVqG00KYOhc1Tdk//Wu/dpLktTltacWVWK1jre4BVI
1J9wBzYKNBLIpFXQkNvDyafYKOHtLoLjhcuHe6lL8u6F3/dlTe+KrE3vynvIQnyScRrL+ssc65wF
z1g651vSmfcvweEQA3xvHTW07AZSQ6FA2g5R1X1HTZuiCcNl8fBsI9gf9BvFTQ3cWkp02IEsN3js
cVKGHSTBEwKJSYB6/hl/VnRObELb+TEaHzfGbSRe/GKJwLpcwXGFHu0K4SjcwzP5C+EBNskAf/BK
pk6n9MxOGYRpf1nBeg9aPsSi5y06Qcqs1rBJ8OoUwTo5O55QCZHIg+bNV5sZ5wh3OiRJZAp6ao6U
5OjMQAQpBZmZQsQjREE2YUhL18voWNYDJ1gZyBK3G1d3PMaTAX91ExfSAtY1+jlQ3pAW7v+bnfzz
DcYKb2Ag0jvm79UlFs8KPUL/tJLPdE1vtIiDBz/y5jtv0KQIE2pXJUjvmMNv+DUuoZvupYQ0frLi
+yrA1m/GxDWvqg+DbELKULrNzAaLy+UwV3Lf0djBLZiuW6z+5z9iZmfXP8vhrGxvXIVl9B9rU+Df
CtHPP9jq9tscPX6jFy1HAHBlbuqyfvSRgk7JOoOGH8W3A9nDmrQ8/ChbonzhbFHpE2Xpai8hFo73
8hD9fi7brX8Vqw4BYI+EsoFCnY3kkmURJy6lH4ZxmtqFNfPkkvx1T33/RABgmwPuiCZ3b7XjRa4G
jTyH2uLumcTuv/0MhoZuwZ9Va7k5BJwNNnAVfuxWui1VIpukrqiF8dUKMncPZ4paZWRsKbd0C7aH
UGzqwlfgyHyfxuARHu07vgze58XR/fZeNuKPSZKIQv+QKDDx/dBXRcEHs6IY//i/jxdFSYHf5Jt+
qmUEqUaK2fxpjyGInMfc7jAwz0RbX0mkqbbJoodJv4emMt8ctzKSjqhU5tbhK3IhhmVmrngmrMiM
8RwW2KdX4DJ3iVPDGAeHstR8p1ddQufZOGkiqOIUNUlMuqVIvleGnUwUVRDMzbk10KuFD+fsi9Rq
nG9QVVnZ2nSKzOM/nXVFbxlEgykR8BED5fpYQv3lIB+GT6tT5nog5Z+ebn/twILiwLS+c6KrqCf2
uFL2LrSUVNFXQqPw4CmO6RW6yqPU28k6UwWGZ8/zWtpVGLnpcNgAznxBONwtdyWqcAbLy9Ly4sgo
db7w1D/YFrlEjvMvQgkc0x1rOEPYCpu17pnGeULrTEMhkwmZHkZwl2bcfnYpezohZpvzDa/bV096
zoSGR4+PYC0Fe3DQMskJWNFlPSuWzk0jgbcXh92zGOz2/wkqH7zpdn3m3BNHPdyxnNYJ+ywZe1iP
B8Fcvu6KcDHwFuoYcwnk1ZGGct9pTIjiFnKaUYMkvcxXVk6KS/p43QUdB3HXb6JdF5hNxklNuUod
zbdcvHOZmY2RwaNxsr1gt4oHXKThIBbGITK23pp3GEO/gOFHjijCiZaasu02Cyp09YYJpl6rqMoJ
P1gFr03QquLaJZ4zFjdbdAyAplO5CthxTvn4X34MNl2Ov14e6Vde4LM00t6Cs+BGNzxM3lAju16U
ECdUkSl6KomFgfOPoX2Y5N78LxLVN+YoXeZ5DnGcffqx4K8AExe0W5xdzSKVZNO6k/In4ldDOIFy
Ktf2yYP1BIC9jQtO0yioy/hre0dwRBoAx2KXeReYKqVkYDXsp4KCnhpPhAphFHL8dcH76yDp511Y
TB6F1C9zdRhVgCsm90UPqJde6V8po+7YqoTfkJD6m2jaOJYiOp5/cginsJCDfUQaPm/HJQ+6WU37
N0zGjc8deVEywE03yYO8mCT5KunTOOnISNI5jH3+j+nEFtdt7ocBZc02NfbhBgpx937XkSN68ZG2
B+s8oMfvr4CJ1qBAqJWOJRdSLSI/ECG8OzgcSqN2Las/V3EavAfOIiPVMpIecyPzxLkssBbGFmoh
dMWccyjwLGb5aVZgbjqt9TG5tRVghj8G/Hj35Rn3EE87z6syShQm2m7N2bpmiEIW7gE9jAfx/KeQ
FZIZkS7sMC3Aav9SiGRRWtAgl4RPT2kdzA1+ArNggeT3mUwRCH5OJuWRJcvsqnv8OrKg14Ce9oLa
fsS68pTI8QQp0+yy/BO1t8lvd/uhoosNFz76Cpz7Oat39JgjK6hI1Vjh/KL+hfD6fU9i/kypAJwn
iUwMUdIp87+9cFJ8pjmF+bOoJbPs9+bFGpS4oklJw4J9d3oUNAOWFAkVlmfPjRl4qrONP8OuMH+K
5B5Cyn1phjlUcBh2/32DpVVyQduHWTNZMjqyL0ipeiC8z5b2PBKpb+vBIVJlYGAJLoJKjqI/jiXc
DbHz2PI5tu3Gyl3fCgNWrK+XiUSN0cta4HoLMOgza1qm50VoyljDcQaSGn3sGjDrkKQI2g/jNBk3
fhnMAhNBidB++Ng3/Eq7hYjvCjEd2Ev8xM9M7+2zjftRQ8MQtFdR3N4OurHJBuMrO/qTc+i4xk+5
LPhe3a/wlJ1Ddl5yoZgDRKlns81mphSGjcHO8opepuyF1s5c3SnhsqkfzqpFUtobnrzAXBLpVVW7
MeDCuBtXj24TYO0ftFfONpvAxzp3O2tecxinytyUMJrXbxafM7Wb1Qhpwci7UcIXi1fJ5merjKpK
p9zd/Lu7HivUd5ZZui7wQVKF8pZiWmSaRjZTrQcj8wmdc5n01KUCH4Ce7EbJfossJrIEYYeB8d4T
fBoygBn/r2iln951MkBJy4gJgqbekruBNMi+jsMLRyXtmoMgge/pj5hqhfaKad7uhX+nk0rajUzF
F9gfAyD4xAyuPhMWa6A8LgbGfI96HWBc6Hpb2FT3RqhGii023C0RDl6iIvXFUxCmZG91/E90eiAU
/HKob3N+7VyvZSMsyoNL+49aDa49/CfY/Vc3y6CSli3qc0RcVDbN3lMrb5fpXLKCmCP0HJb387UU
wH4STbgXKjhLihafab4LeyzPTy/CpaotX/j+XF35hQaXamr3bel0WMPyhIoYMkWbhnwOFqHuQleM
EucBtLVYwTRlatgEREV++LIqFvr/59UeVeiY3711WGibS/7xklltfzY5ph+S9Ck5lu34yKKIwRZI
ON9guguZka8tnrjYNVVAH5Hfp6lAWfvTo1KcldpC+gCknE57pulqz2V/jde43HfZttf1b8iQorrf
UNMnLfMrB9AK8IxE9BOrwmLadFjaxiPIxVLXr0wjTfswB2f4K7QFfN3l9QqEfunToYhf/NRx9OIo
AUES35sA7dgK3Lzzz5YaBJ8qlz3TnVi9ro5ojaf2Q40nHW3hQmU4Gu9rTCKIntq8jvXldc3Tfr+J
/yZjO80r0rRBi9BT94As6GU1LuPzccnwFxkdPJXQiW/lMthIZ4QbyrNX+oqmtYhsKxDHaTbJRefM
Fpqkn12o9CMbFWS/Drwa4fQ1TV8T58gPwDTiiwGCZmh43M8e7ynYZLySkCP8KzaYBK0LNl1V26an
kTu69I/M26c5Dh5SqoSxzevxVm/GC1Mr26TMtDPexf14eXufAXndOd3FnWYsBZ+jodks4jqKtfqs
FI/RPrLH+0FXNokLFxoEtyndHxj1KEXKoQnMoj0NRjlUR6b8shKN9kWc0j6Se2czTlmVmUKUIA0c
hEPMXQfxg6DzAFWgyLNF1plA7kFd7MHNhxlbm4P5Jqe5VuPe6b6mLlR8obFKcRfMOTd4w3RzY9p3
Mpvcayg52gVwVtt++4qpeZgI/R2sOvPVDrgdLxDOfRzG2R06QYAWJ08B8i37JtKJGa/UnPrAX28R
Ngv61v/IHGm7Fx5/raGdChqNBl2Q4f9yoIzeTaWrq5ebqJYX5pQ4SM5rWff3eBtKliYejuQA25e6
ULZULAYXkQrnUN1sI4JkEDQ1Xf6yE+w0hfS2aVDXT0OJjdJMBwYA/s+TUTB2QJGG+oCJTq6AlE7q
Pfu3Ih2DeAc8nlMgN2ZvDSVGnDhA3WGQeVImGKmwH4+vI5AZIb/RSZASTyln1qYd8t497mxjfcUo
+aT8aF+zbqj/CEeY9T27x6UVOijws0LyC5ovmjL/3qfJONf21vaMUMZ3xTUsuJQrQHEBq3gj4/8S
Lqi/iTrdemhkA6I8PD8ygKRE9Gw3I+k1F0acm2WVz5Og2rjpQnZNE3VizR1eae/On6l9tAspUhhf
QOYF8or6tOWeEeUwkQ6Aoz3hlgKsqoZGeIbqd2MJuqEnmORiZAqFugWdMRufyGaCw2ISexPt5RL1
EzI0vnZzNCRYVfAcRTb3IRHOnbdxNmj1DQrRWMiMQc/e9plJ86Rw3UVnCPKzkIeZ8Z4JH/4bcXt4
3Vvr26FWk3YzRDbPcDBmVt9fs+4zNtgvw8/+sHsPr4E6eJVVCDZv6ui1W6r4jnYxdC3DaP7q9i99
jU5w78w0KGVs1DVcZGp8fyiRkKMeDrnCpCQtgFEqZLNMk2g5wO7rMIqfqfPYJahazYroiVh9k4ip
WBlKS71lgYNs0a0CPtqqtQ6Uyi+Ql/x5DxBeIAzjWMb88ka7bmnmvAepGVvfcHTOAAdV17ZyvI6N
kgr7jwijoKveK4zUj2nLd9kt0HldODpr1BwpmxLKonBSR3+2ikmueAGNOxie/kRgx1kY+fOg+rxb
18tWJc+sIVJ71tVpj65peWT6XqXgHDabuBmGLFUypIlgIxWbiy4yrLNZ7dd+1SvoiFbsk4YbMtil
wx+aN52p27inWK8pKp4/mCN7UeRi1ezbVHrIrGETwNV3pbU67VgYC+7qVsMxrt2ID+WhxdCGO2rE
0T+FDNnv/7Th9i+6SjUoXTgbezoyI5PM+yG74dt/z2DJ+sxPdL5AfSAz9yyEcMhE3uPGO7bpF3/V
pdrZ5cd4A3ZiKzoUW5rAHnzbxzitM1p4qYG/hTxTA1fz9QA2DA2sMYwn3oATbOa8jZH0lQqMNTEx
OtoQQUXi56S3eXe/4Gz6Sr6HzmEEUAwI3wPkJue2hUf5d7UbZ5g1mjkjM46nCNqhfBESahLTDNh9
qmNRlNp7eSdI+mQULo20RvvC9Gpv1rskkNtjXL8jnQl+pq0NoCFZRt0RqyFH7rCmT0AgwwPB1eFX
/IBi+2rWU015jDbGkSwrd3dk4yti/L5jkFM2jehQAhwdNzYSygQWbwGQdHF26EBKzpg0f+Pu5lkS
M5VIfNTBNdlwqE0flCL7AZNJSkaQkbfEvM5vYk3v8CgkjNqixNODNuIZNwMY+QMrIp58hNyJVsbX
PcjlBJHP2pQtpJWnB/MVagmBWMt7gR1f2IF7xE5ZAObw8C4AITg0+WWA2WffDaOHkBl1KmO17yIa
LhIR4o45jjrmwqtZPI8H0MhH5I7mbo9PrWBjJnxlwBVlJ5uonm6XAuZF+ER4bogjO5Mk4rXyuLZG
UW3VnsKAlBTgdjSzml1vTYjmivSfMfTx3BsFhF4eFrgNhk1T9doCcM+OAiJqdpF/pu6GV7FDUoMb
LM9fArHCCxtwOqXvS52b49KJg37+wRor/NOt18HUFv8ZhuXLIWDXByFJuplNQO5KPzikxnAlLanI
FKztUOpKoLYzd99W6Zlo08bpKajIAfPKu9trzkWA+U8IVzeXgwV2stEdq1fOeCpi2ou1YqV8kVIb
DSlF9y77F+Ec31JM+GbJ6sVbH77SoqoUprA9Eb8sqc15/AHPZHZ1D3Sk1eDhiMBZ9th9h2dFZK6G
JcYjvnsC9vEk1UGpCWx6j/zXDRJ5vtRnvfJMqsCAlI58cU0EuD+RZri54f0bsq/S3cxzOmRFbOJO
Lgzh1F+EmenKkTsUfkXQ7bgXhLVlQh6WcN5g41Wr9DZd9Z8cxosfPxQW8HB0erWXfMQK5hfg2ieV
DNW44Q3bqMRo7V0grsNhpUOzZap3Oddj85Wj+3mWSiskh186imeFgQqgbBQCXrrxpeXbg3bceB0l
YTVKRbEcjkXgaAaZczb8yQvlYe0lZxdL2NmKtol2h3owv3LcHP3TTPmMiCrR7D7TYfiH49kfJNNT
8Bkj41UUO/+1mTNcBMf7csllNPTcHY23jsIbpqdevgpXNCT4kv3w41wykJwTpkV3cLeR94lMIs5d
PJS7rKaEKdTOcR09bGUp6Upq/5da1pDvp6yAs1HPCvuHr8Qe6VAG3HcgyDrLcmGkA51CcrgF/Pcd
dMrlCwDQ3E9USgGTuuRhpcxN4pprWQwOTbxPa5cvevLHVmtpC2XSzK/tGsQs3UxHgLCZf1kYLml1
3wmVrH+LcAwNUduTbOwmhbJdYEzBdbRLfpAHQfMWlmFbmaQqnPIGlwQ4Krq9haITlzou0U328OOd
B6mqdZeA3y9+FJIS3w+mn3Lt7dR9wK+3Jit7U4b0pug8HX4TzYWa3twoE01VT6zOnO162cYF2Swj
UtEvhL0/xI2HMdpxo3e6u1UL1ahz5TQgBuUE7Oxmpdvzrjsf5VZqKmgFHs+VIxGwjw+sJk5+8hCZ
qrXVdj98I9sX+muPB6PYKuKP++qva9MS9owMK1qbSSdem493lsSrkfPozD3CxNjACdEKLOcO6CcR
Z8SZ9jxeI33FOSN1Fbt3pS+OQ1Ae6vaFR2VIJOKLpvc2AmSB6Xx9gRjzzYhGkPRtB6kcWls/MCNH
csRwuY6fLJeLmAmHEIvp1MsCOj7EemY4bk/rjS0J6fJGOVWDO7JLpI/5YsG5Fmx42WfQDauI9HZf
NzSVRGhS6dsr9+MElv0csMBN6Ijw67viHUuUHT/jD9yiC6I24gYxfkZffOtRMTn1+S/2EEp0B8aB
ChwovahKUsCx4tlUgGZvlhqDfIfvycQrtwTaHRADEtnk/V7D7vd+QM+jmTfa2DhP6b+sYLwRVEj1
o0Wm0S9gx5ehd3aR37oMUFmciKxDRXEG4euj7JWd6mq7IASx0cdA0LMDmrmM4t3pLxPKasrt5wZ6
V52SMuS4W/0OBJx/u2/SAdqYqdH6u5TIOMayhpEnMq9k1ofQKzIl0yu4APxorOKlKKapQDI6uyWB
pQ5fHdVoZADnpPnhFaY6Np4SjqF8eyc9sPo18dYF8NKksWCL6QPSxQ1BM79NIoM9IFvhpZ7jSTY7
RWWVPWiVMUr3wbbtAVnMTUCjEoBE62pYWU048OQtVA2U74N4M3n9oUT07Lw/XH3ztY1h9YqyAUsZ
vlTGdmcmdhrsFAXUxLxC/hDx1+onhZwRRTUJwFfne9iPhuR/qwU7jB4gzjhoAxNL0Kz25J9EMWPC
h3HeAvAbxdCNbLOEg/S3j/Sf7Aa8/HQKgLOWz89eoAeOjQJNOwqd35K89oy72exY7fUyNwNb/ZQn
m87FhS8zpjL+Ka4y60jpyAjYzFdYwjzYIfpBtwUy3kMF43BVmh/ZUZlENe+GIruyj89/bKPdQUpT
kTd6NVELMZ9bASkRfrGvrWIVFDMYgPi3yLpf5ezDZUnIbwYDrj1U2nm56O4cC7ibJkU87Z/MbXAU
LvyRYjumz9AWHMd/iqquHPEuM+WqJCVt/ESeKPLo1LX4maDpWq45tyQEThldIFqwXFAKL3iXoMUq
enG3lthSj1qwEQ3vzWoblV5ozuN/kVB+rnJqJh+VmiLHJtYxZAGoSB2bCQlRnm0muwJW21st5EDT
rOLtnci4HWd1hiwyIFOSIYMPC62xXceSIjjinVjybIlIJtdF3QvW7Gi9i5HJA8cXjN7fpEI1cMYk
cnG3dwtDDpCopPIHTfjs+TdvrklWg7o7TENpAh5wVy4AT0PCmKI4+FWjwYB700/L5gO3q6yfAW3T
ZKhiBKLM4A2tY/z8DGmpwXowbXzuui4tVV3vKCRt0eqe1RtjWeJlYQdcBfORxtOn+wChbmleHtRJ
MCKh8HbEUE7ZMCZ9WOaR2pioDL7vq4c3AUsHS5Lq+/kr40uKoYnaEp1/Cia2AeYrUkHUYn9VKMNP
i6/h7R8OktRy1JEOnmj2qfQxYQZSQTuOh0mOkvYn7alFLM3euaDDmfld4BHOdNwLmykXPpXwHaqH
Ya573BFOse7qELcbnHChWVQtJS94rCkZJQkhCHDPfznQQocOqTvzRF71SokfkfRuySB18JRSmfsI
/tHRhIXluhqTRiPQGEzrcs+epfOwoCEvUZfbZkOgdpO8ufoID4btaeNt3atlJlzafvYF5pPMtUrg
nqwlY8CH9sC/nngtoBj4Fw/Rcbm9zahHmazQFl5FB9KzEz4lIfY8zvWItDl4m3GNa2QVTAOeawuF
lDvgvLvDqmXQS8C+tk8sbT6v4K8mAXBOk4/eC8ef0EfbzOy6L1ApO68rdFFAKG6xgTI9qnCnioHU
CEuJ2ix4laT/WS0YUNP3KlKyf31nvlS9kDScrcCbn479vq9nD5/XwljfXsGlx+5Nlf4QwP/ixLmw
9AqAJGFyZ1+8vuqRf+DAdL2aygOc860J0W0U2ZzZXyewjHFMiFBS8T1XTGw4tM0IoB72qGxKsUoY
hSeRHmjwbdn6kRV+dLmBrcZ71YOc/L+1rhBNoSqF3BezortBJaLCcaB6+2DVnaMaRpvPATYIUR5K
WUvM/v2y3YzKUg1Wm2P/6Pe7AsNJ5323MX9frOceee4qnpKq9gwwyE3X312Ywdwh/AwMKk/nnG6d
NkeVE5PABxTkwOX5P4JURuae0fLFeIQMa/FGXjx4WofpAEBaSWH5S5ebhpTrPQMbUNrlYdZ2MT7t
SKMmoVNwPYCK+ohSz9UMhUGljItqOpsA2JOyTEk8ksq5jipzrUM1bRUC+cAP2oHlV6wr6quwVE4g
7p4w5Rs/MhKZ8vPZy0M+i4t1TrxAliZ6stvfsL6f0OfAixKDdzqDWJYSfYFJq+dvuS/TF3fAlBBy
Q4SkBZxH/4PYQMlwJsLKW4fijzvdOvet8gB7hGjJNEYSZ+w7UpI57J5f+kCZNe0mtNPgPuq2Tzki
NTM41AK67gJP4izQBTawJVg5QTipg7Ben/w7i4bdwwq5isyvN1r2ONPX53OeTGmQ1pGxOGV3C3B9
/P9yduImJuIodZVpUsHsBrpKhz3ct0p+bqw83PnmRanaeYWsq7JNIYeyP25zEouRasAZX1y34BV7
cBbMVj6Ptcponhwmvz/NNUR5TAKm2RFklxEf71G9EDDYW3hGD/gDrpmbNYRgMmmW0UoqR1tjDie3
OnEx0hN4MizRxARoqnos+gxxKJdBRhwFofuAdxKj2wGg/75tzIwIEwsE6wOi2UI1T9G929lws/pW
RIMjnfV6DMChMNDFQPgfOfy7A9dgz3Dg5mcyQ4CTgB4g22kBk8WIjk3+JugGbyo0GEvytKt5NKl9
93xtc8RWX6EvdMvmkrsrNC72OFokkqWvHHvgMBmXWMfU/kcnyd/k4i7pHgzSUFNUXl1m6EHi6tao
Vvzep/BgTD0PkRpz1soEbgaZwQ20LDVSqQK9Q6G/fKDr0rI/sSSXUwJWsopmCiBbYPvf53t4K31+
qufIj4+bAELnIlACCiFOTrnNGHhPiyrjg0OT2/WCutW20YNf5PfwhvK2qqPDvtA5wJGPwSwXqA/g
J9IXSkLiVSL8plwy3gX27HAokyvB7PH1e6D0yJ9E6SkvHqwLdUrt/u8B2+p8qaEgbbEyYz3ccoRw
rkdJ5KWEEDMgEUFBpar37u1IVs2iYwfLiITd5etXB75vm6NyXr4hvyvWr/toq4duB2ZJRCdP+D4y
3M6YfUHBdTjLMWtTHhC2KlE8nEobW0PPcVwdZ5/BkbUZNP3//egsxTjfrI4DDw5IWwaRkaYLu75J
3ZZuvKRx3Y91lR9S1bZS9/42XwmuBPKsosXRr1tIojIP3m+GVC9uhTuz4fWsdxen1xjdG8WNrV0m
spUcxckOil8aGLB2F5yJ03PAR2me7UTJC798cELuG6LZAavXqHcPw59F4XIUcmFfHecd09x6aC9L
oxUM6sxn0Fkz0DBres2hqJHRHwmbB6eKlG/R+FLBHT5HQoh40OJxVGqml2uxbCI2jVTSo/6YDHk0
qRcgDLYHYWxW3cBZhZ46Udk3urGJ1m8q23DyIkl0KofROdzrNNycNnZonM6o3YStuhDZ+bOS6MAx
3FkxuM7tOWhuAWMGpPZz+5YHqjrZuk3CE689jA/8JAPI12MHGQdznlF+H6vDTAQ0s/kXPiQBGeG3
auNJ5aODNrdwwa0HCFiEa5+YfE04fNcMVaU5nXEhcmuX1dxtb6PDazAr7P+MevUiGl0e8v1lsQWb
HX0S0dNNQKAfoBZ1KQSzhRfftLmHzjvoEaxf7uWu4RFNBRfN84fsm5DuM5oWZjSDG+mQT092QLHp
g1OQ38OEq5JgTwitvTl+Cn6hLrfeKovi0R4WNLTxJscqlC50zigTchksGGGzhtKRxi1ypUG0fzjo
jGujUCGpgJmQ2pxO13dcb0lgnOOKNd9ANatpoZPb1Rw3WNpMQ98Nnj0cySGsdilrLftDCGNlL1yt
+PHilUjnh+XeO6s+JNLeT8L0DkL+ctB549pQjs04K2hqz5S/tA0QnayMZ8D5pyYvwicFOI58Uivk
Nt33nnCLDADbmo7x20KOAhb5gEhZB1vBwhqyjrORrUu0NNfqE2q5JTweWUVOJBRhoAvkxiX8iOz4
94vNLm69wRHC0vsQMEvStshr7rFHI+9Z/cU6N9duZPlKNPRUQw5KLC0APkkCuFvd5LBTfvQ6WwTO
1J8xP89FpP7lAWy/41UOBd8mtxFcUWqFrVp9UsUku1vqU0NeXfcumNWj2fcxKIWmtsEGrVhPkyxd
WsbXD71GmyY63mgv7R4HEhNn+dRTtJ/rxSPuR42Bq5r6VYOwEQY4W7hQdzpgIq5t4aHBMlVR++5j
Gn2MwO78B5HVQFRRnAT2sOyThPz/5XkjBFhSdVH65PEfLbLsxdKXXMM1U9I3Hl8d3W1PWwx0bssP
n1j6g0BYe4szYITgOaRX3vD4ty9srJzdJulVRfPurVxxSMgh2mnxlcAfphSPAQw6izzyg9BxSaiu
7xenaD5mSqipwxd8NlBe+YrEpbpf5foakh28FgWYNP53D7p1nP0CFTEvdC2Z9p7fydvTsXypyHt9
nNeN7xB0xt3blsGi6BM77kzPs9BDbAe4ta3GL24pc8bdTqV5fABj0RUCqO/l7U0fn4wvhem7dkAP
pVxfSdfs/ban4sJE5ZxNYEVpAXLvMfiUCjTLvfW/+ZZfLwZ36J5O/NcyBgY7X4AoEhxokW+hJmJ7
7ynWqTC4pRiqnEfw7aX6tuDalpC1RUsD7tIrU3LxN9u5nWyd8aXTza0VZwA4UpAw+I1caeiLI0kK
2M/B4yqpak9adVznhuPd4VkROw+xmyiuJ7jIP9G+bYh31JEhQ8W/8hO5X9y05ppLOmY0HOmd6j+1
9/1UwkpIQVfJ1wLiHJJgMi8laDK6Hc9A5yESk+X5FVt7k3nGU+BsNwpJioBzHBFimi3kOG6sTvs+
rHYsY0O4Do3PQ99D8XPR6nL1jjEsTnby49FJC11PuVQZ9fLXPTBf6vPMgJF5otsbpDHqoAr+1VqM
wA61ksW82DnUSqFrZ8r5I6nas0ciDOUtflU5PqEWYY5xZS3DH+JqkSvcwiZx8p94H5Ntw7WUFFZG
OCQf5qjrz5sz+XQxIiFt/TryuARu/jxSLQBoF1RAtXk+MT39tg5LJSguRFFnVlCYRxL+144BzY6p
EHboLOO2uTHtPzn5up1BX9TcUg/Rusxl1iIsripmKoadP78k9Zunp1VdmB1Ggj+AzbbEICEAtmIm
U7+YScuEG4V6PBihbqRktWQuc6/xa4esu0JtH+V/uJaIs21mbicg3ahRcZyVmMFadSzubGLqD1TQ
JkPW3KDtY7xD3ofhyjvXIMM9MDWIEXf049k9qfpUjY+qMlqOSM/CsF7vu3i2tj3hGogmRZ96PU5n
WXfIU9Y8AN6yfHepJwR52LIkFsx2j3f3/Pj9gSxkIhPw3hDlsgdXFNJm2UhyeA8wZjFQg4kRQBl+
k8Zyt53BLfEnhLrAyWjOGhyyd/1lvBd70QmafNFdLCxwGjxLluUlCk5Vj62bRk3q5T6q2xfJkiF9
9nwD739BpUCXiRXaHHxRG7puvPDUIDplX9c0o1Vcr8uWpN0bVKbDzWPU3pT6LY+i1KYKXEuwj5c+
KN6IWzRQd/RKzUJlYMV6R6DM+CT2Lkkj+cHVKt5WhSrBJoZzi/TZfNuVTjCpn7pHqkGdWGXdwGGl
KN2aBTytTezh9fBaPqAMtKt5ma3rYgfRDhXbCQYCu2+obQrWEEh6fJFUEvnCsIP2ETXS4Kh02fWM
rTv32koN9cF5CCfs0xmHO9n7SEOmzDWiBknWFtXSPTX9gYADmE9IKdV3a1an8xBdGp8gOqQV9e3m
MOjNDkjNaMZeYj+NY4EPoWwEXFE5JY7jT6dIF3oZR9pfMfX6LYfSYy7OShUrHT1QanVfzzVPMorr
FjdqhvnkAsF29ORQ/c/NTANq8NcH/X6RR+mtFJJQNc3Dh/G8nTVLfz5wbsC6yv9ChFN7T+mcJJr2
CK30PCFd2Z9VwjM1av7ihexzsaHdDj4fj0o13vw4H4tPopcVOn23/DS2am9XbMoRL0yJDYNflpDo
Svd1NBZj3nDEslkldFn4nzNu5/mZekCpTgcbG2zwNnx2XxBx/QzmYkutjYF/jqUTRPZhKKn0Nm4W
oCIduTTQduZBr2F/HdxnoOr63fhQfI8/r7yfXP+b0oPSn+VQSofb3IryCzGHL8Dmm7G5TEUuzUkL
mxZ6lkDTrTdtOLOM54EElBqVwZ3mWeEc56Hhy390iRD7a6BEwvtga0OvOiDP2/BwiNNK/PHOPsbN
aXOWhGP+Lb1PPI+0FendWbF6T+sjRS61DRPGi4QI3PE8RevxyDaWiEjY93jeUDIJT0e6w5CPveq3
9o3Cxe4MrNTVHWW/E53MxSStodle8MDJkW+R40647oE4YVBl3RuTuIREGDkowH1mfRIKaA8Sj0q2
bv/mpHhjXtFKn4TbXrjdzZ0jKXyJPKGEt8G2zEBAp4WW0Ys+bvq24o/Yd12e0w0DfNqY+Phbf2Rc
ss0bF5VzWcLdxZlM8h+gmyOBEC90EjOPOHZEWyykhOQ8gH66uuahxoHWpSzPy9uv2VxeasehH+Fl
/cCPmmWraOC0EbGfmCn79B61J9ppV2aXSgNNpeaHcArwgvFIfMbBYdif62Xde1HEoEP3CQ/U6YcN
lyjE45PrR7GVShGNiZfog8kXcdKw3E6dIZAsU58BdggcNE3JoQa3YQ9GyzVVEuk/hauUSmUx707B
iufY9TG6EVS4AjihW3cDtBxQBgVjsk9Dm04E7GeNtpl0Y6GDDPYi/+1cck+LCGNJf52I7njmk2vo
dxkNf8Sgg+H+aU8GGROiALvJ5Xlmy9rTIfRbN/Bd8qXopy5itoMNn36mGNaK6/gq5tBcLfDWLU/E
4Tx4GHdhwA4pDIKiPNamJvPwMznCueUX9f+LE/lnMoTpIQ1bBXKTfcGLzI9aZR4K/US48d67UWkh
UlOiID5RsLi6vbmdNJvzp0ebaYcA/lAEVkL/wxxxHq+A0CePdbBje4XmiH89EGpjq1ujBlFoWkgp
FKFZiWFhjI2g8HabitDn5xZyBUZOGjPYotZBvaSN4TVmiFRG5jsRNI7zyC9xMQw5kZOBMWLw+Jfh
c9e37gXABwt0iLBLJ9FNvK+6A/GGBAncecYouH3jLt2OzP9LBetT7QonFpImS/2cwBf3qpjs8v9V
euZx9i6rw5Yf53Bf2HA2hdSqLQz4vtY3WRNP92OyTBR47t0o7q+wraNPYf2nfwb30d6ZuyL5Onxh
JAvknKZvREOpKLETv5NN8LVkV6TpYVVDbw3AO/UX+1ud1hFtE/XpY8AuFgFRt3eLxWmWPhIEclAb
1WT8szKnG9WOZqDHiLeoKXddr4L78CsXH4U1ZkweaGOtdr29l8wvEyefQjwaT0cNMFQVc58FDYWJ
Yhe06jGNxcvjxBirkCrvHoVYCHK7eRzg+zzbuiO83RjRLC5I5GnCj8zITwvCj39rErkBQu62VjqS
TfSGDKjHLLYHlvBZQje++Mo3k5RotHglx0H+6UOBi+GnbpMmpdz7qRgThL300kGYCHXshn38rANy
N/Kdkpf/343x++p20VaJM0qe2ypjXckmldBdcx2YV3ZPIBxK4Gu0G0znMdSeIKRxj5ljPhhHbXV3
iGD+3mlFiu06WsE297aHzcIRu/yQf6i2mLif+xdBaPIxm/hSpMwiHPZlBu1O4mJgnkRG9jIraHgd
2j0xI0XwE1lzvWzez2Hfv4/Y5TOmx4E+QNs29gT6X9ZcOs6QzVCMKRYLIJBzSwVyefsSN/v4kUiJ
LvLCiGa1QrMKvtJGP8nDgwRzSFYpeCkts+7aWX8mXBZBy542FtptcGqsg0MCkHfG2LEQVDaiYG0C
J3FrxQF3heQfTHV5DkQPQXLK2WQIGLNzeT0gQ8mMoLF9B/BcHVFm0XC71ph3hN3esg3ucXnUOGw1
KHs6iGXQWjwxCYBO2Hs1J9/wqrau3Mk1L5aR8MaqAGsi4FyoTiFfIruDJ4XT2aA3RzmYQ5xSU8mk
CpTsoU6uKu6nVxiDwUtwnOb3EgJkkHGCWloktEz9EbcnvF70XEdS2Em35y31jvUFm/781AkF8HS4
Y7UAwG2A8QdBbAsG7im2amsKZ+jOAliRJeRrlZudw0f0+Jyl0wx/3NB2rJsImLHhz7qlOFC6bYbq
Ptjl7t+OEO8qCET1dFg0LvZn9rvwaqO7iyUwQRxDeUyy0RvdM0MUch4s5tdYzTTevDMl++YpKsyQ
oRceVzCaY89IpN4cvmYjpQPiNqP/1TJsMP/oDbH505B/3yACU3ZvHob+h9WdxCyoTiIjsbicQQ7P
uGtweoVHEAD6OavVAzmnS0XviEcVhUFLVXwnBSxklHilfsVZ1qWI8G9PI9R1R/3P3/m6KHISTfY/
aw2x4gnwY9J4nsDLhWQ3Dk4/zVDhCV/lvAt1JNvfc/0+ccAwoOCXgA6DT9LFX4tlfSYHQXoaeQVE
icyOt1+bbi9oe+SlOcv4UnP3+LtbgQ06or7iOjHSa7X5mBT2fBRUvG1Mr1ewlQBwH0R7sA5r8IpK
/2Il17qvHUZ7pivYOPO2PNtww7OKH59gEEHPNRelH3+xV9/q7Dl7+Dr1BB4ArYWavQiu+JUHBGh7
6ta4V/SYBt2COvlZJo7dnDPbTWIiy7Jj/tE0Xy86zlExFNS+D+Ry3Bpi6H1qG26LDTkjPODHmS3R
v9TmOO0CpBpTxb53OtV7+XXrIy3zgK6AeaxD2jkZUalwFf4eGmdLIfL1+mw3x03hBxlZGLjoZFvG
YLLMrlikftGsZH6Tor3VJge3hXNpMHigck+KpT9S2LJdrdtbAXKCxH2nzdsR7Sx8xyoK0NT9PbrX
l1DOP0Q6leE0P0LfWbzjEAd4N0XPOL9y6C/AYNUWwFXvfRsElmZdhkyGUSAucLbVt+KIC43YBPtQ
vP0u8ebVMG4Qo3LXtbJ2Hp5lIkFCFdyd1M0QEruvcpcnh7tsSlIyESyt7A5PKVJ+RjAl/C+pWC37
VDC0+J08dUFh1DUsZ7yeFIsnOSq6+zOSqSD4ZjHfro8gTFAXrJT79c3oMGn3H/LMSNy3X0Z8i8TG
mnfp2TAjfL+FUhgYjtPXbl0/40ONYft86A462QKSfGS1s6io8rJs12EYaKJ0Rupm3E+IuxV0Xd9z
wFFkZZ0DX4BfTjreZe3yXyVEU+VLvW1evgK4mgjmUEHC+bqhonqE6SJ5QnALZ7uVe38wTBMp3gig
s2u+ERZ7tk/H3d974wDnr5RCr2jvqmUue4yC0RRc4gvCfnKBGPQ85YktnNX4A/c4Gmqq3VmBg95p
1jECxisTMXXnUHbZ+Qh+KgwQ8M8M0tHFGgqzgyQu3WVT7yu83rKhACdZ6ToPC0/mZE2b8PPctMn5
GKgEDip+WbHWroYXrPoKbeTm42i/w1Zh5tAYZ7dtnBmoJ+0C5B+GbGZKu4TMBf8V7Pqq8ov26Bup
/i83RjuR8MmrzEyxwIr+WvRha85/6gjYWVLNoTX/rH0jj5O8D1lHeD0EuKQeKMR+GoSeIdM3gswC
fMNJ2gIdxRZUyoaxEqtlESaWLPlXiE5OZwDbgnzvDs1qX/KBZaJ6Xy1ZAe1qyu9PCWKxG4WzCG7F
78Y0u50gsJag1sSmh+CFLKqBfxjwX7uxpclhjtwGvTN1xaBs5xYRytBVwA/xDns3UIcI+73DmPWn
13m5T0TAn3s0XxwGc4nSCNiU5mAKzMvzETrosYr0wCpwPuPoMeTtMWTZPIk0IsqCQdxyPULUylSL
nHYsSHHq0/htC5tURQHcgb1XrxVexXSd9JAqvNTbGEVmh6M/wbtp3KMwrhjxsATWuz6l23zCRujJ
W4LnfkgLl763TMh/CxzEmUnV2jNB4pE5iKA5nw==
`protect end_protected
