`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
I0GfVFo0NMQ4T8uYkL1/c8v6w0Q/PG4vxH17LTfjFM2X/w0oeXaigJahAtI9AKt/JTvQx4hOIF1tSiaiMyjeWg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HOsZXrr465l1Gp7XUKG9S/JT60eHgoYJ4wy3sb/wAu3W9UIrns6QSz6yGgLYTJnrp0Y40EOk4ADfjyWB3gcf3hQ2MX1ljr6NLXR7ck6zfmK/XzUxWQTK1CF6W8uSt5FrO4aqHUB+Btv+WgJLWyj1JH/WhXP30Wh4VPqqKwybO1E=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xR9glEbPcZLd/TS8LbgBz5+z0XSt0RF+j5oRn5yTm6k8unRlqQFo1Oaclg1ZJknJtDmPp+3Hsexq2bcvj0NQ5bjim1HMFbNBhi1tBH7Av7r2iOHLL2TGVch5SYuMx2F0MkwM3rPmkkgECpIInV+OKFnUB4tSnS4m5ornGDFHxfrz8KIy23/OddE2dx9A766bR+RdF0QDRzafUHvIwBfcX1ijObgDZkQ3LVJaSJmW1BUykr07kqPnFuJTdWLkUQeDL+VtGJ1hCDRjxwZw2/NArDRUB9IYt4E0P4BDS9aF5z1ER9iDiq3k0X4mFgeMmjWy/QWFLh9bHg7/WWwN2e/lHA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XcsLgQxMvWow63pTVRB6R/GOIlrXaCKlDqcZGJq7jl8FOmp7GK4cwpeYQHoM5doLjnyRXw8AOtE957RZrGecxyqu0XH1GmBihHbMcSO3/Uy8q7NxXU9vt8gO5GIrPmSCfMRjCoy6GCYWz+Uxp8lHP4CwzWGTNPmzDAaRiSb/P0w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M5K+u5nt1gTyZy1ZD/VUg3iXAKmLBr6wtQ/rG3jT9diVtmuMfdqsmkbjmCAzXLsR59U9NkcqebqUq93VCM1m4OUyfjAIAhc3jVx28oTAjb14nah8EUMsJ34dcHgEsWfQl4I3kl6+b4RkNDnPPRyaJIC/W5s9Zp98hBAsFbgJLXmsTLix0Z4qH0aqsMbuCVcK4sjo+nE1l1PcuH551VeT218NOZ0B5baa+IgGyZ2oZS5phfQH5h4z4nFqIioW2Gm+44GFB3CjKHHM7lQJM1+9Lo0H6Olw1TmZHzyLIp1J2pTwKOk0qKhmmNFV7bmxt/onBWyWZeCQA7zm29SrHDct9w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3614)
`protect data_block
oOb7qdh+CLzPFMi2H1shSKbadYw8pcOBCw4WWHDGR3uEXs5Xz5VOx88T+LsI2Rrw8+gEJoa0lbc5
Ssex1j0gG5HtfyvBBJemJK96zGbSusa/95eo9KMdPsqK2QmxCWZ0zqa6h6GDCiSjCML25veah+DB
f1fr8++qllBQkR/Wk7tYK729fRIzQRgyR0PEWeVTmHyxIx3U5wgTnqmBfZCiimzPtZGCSCaRYn+2
cVvxnasGaefrThflHi4Jh36d2XrjXHghfsfklSJI7x10LuXV3efyfBuq/94ouXhZ7OYp4Jf7C5de
BHwkIyLNH9bAZvLLMfiHG1ax45c7yHAHY9ht46x1fGAX6zbCm26+C/Th6VgnU+MEFeKEAsVNEgtl
uJjQB2w/g8/43r1QYrqways1QATX47XIo8zuMrW3Lx46gjhsiCswcBG6r20oT7e0IJXJZu+4jIsl
GrC5pxmMJ16uzigL+I8t+3Yl3ALSpJF2sma5NrAkdCyE+dxi9GWhdOfAubi7CcIBMcwBUm5Tcje5
NJdllzNVwoExAgjBrWmHop0IwdIXvM0pPRf7KwD+ubwlQHrXU9S/uqNV0QpvuVvozJIEqKor1M45
/I4iyDi9lBmyMZ+82DCckc7w0F/jR5tyNKxUZ9+ERx7IUweFPGdatMgs1o7nnfRNQOz/SRMQNhco
blBzawxKFEg2/ceYrzxucU0hdNR4+/3bazc2KJADKx7CH8erSfXQzeoo0M2NkQzQJanShyvN0Q3A
wITIaJhcnWwUKSWvk8Q3SPjbCoIoaaDNGv1vZl/FjJ6Jsl/iixqdGUx8uX5SaAvFiqR0FyC0qCwi
ZKPk9PkIpllkEHWnZSKYvkbeV2ctkzPV4rp02XBG4/yOYo2+X2jRCQhB5bgKDR3sPVI7jT5dwjWg
A9b1sqV5qSeLqGIAS2yI6cWz3BgxkDxNvn9G03Oa4Ie4sbbKQaWjEvZplgzDe4MMEonPfe6sVFyJ
JcudiEDHWVDPJ6UqHFAd9YOkyRuOe/nJsWpO7qPR3Pl237uKr7KpXSKm0tySyb6ZZ5ltHF3YhEXa
1py9kqUgq5PWgMdJx/WGZ9cBLtSLuf1v9XuBA963ApB9jxLqWgaaF9cLgLJ3RYIL5qeNsDYXlQQF
dWo0k1NDylpAXnhnfpxlwbi2p6C6P4QMFTRlSV7eGyAiZfb2zkOTi0oyTk2ijFeBvBYEtND6SPgd
PNPegT2K6GdwyZZe9Ofn9mLahN9X8JBvyF1JY+lGWXGBmxfiRY7i4+gjoaUzOroBpe40XSx2clEc
pTD9UGISmduUM3wz5pfnwth382OecyY90HcEQDDbKHpmKHl7mY5ff+0N2yieoR/diKKipQvbFmLa
L+IdkZmotzVpHoriapGBO9xSkBm8VtSHIJhQ0am/0ci/fazdfL9w3HCmZirVuJ2Oi5PbXbif4jg5
Syj4M/ytuAnEl5+FT89zAwbqPbMVb1EK+XfyHN881QHYjp/RDKdooxEEGFOcy5LBPPofFIAil+K/
GfJ183plMrxJ/GOMkzFOaJRke8D3KMZ8N87+AGR843gPOcM3gfc2DpJPMy0Dg6ozNDPVY6Jc4Za7
9DrIZgoR1k60McN1BXUpr2c9U/4s2TfDzcf+xK5azkTiH2edxy1DYi6oGMpXhRV580MxCgmhBh6X
3EcpXqsNHzUoB25GOeXdR5VPcwDm1DunYlORxCzddnV6WdQFpUHh4ia8Lw6XTZvPZ+1v4PAb3uQz
ehLE2HTdZXK/DRssRzEEpE2EyqMSwUk3xQqnHfrUMuRMnxFw8CuB1Bk9LSjWQWUyusEZljnYmkZO
TEBhrAyFLe3tDm/JIqdSqX5odFgc++f/8RGsBxNmcJOfM/C15jzoBoxKMWkAS6HXvHp93xcV96A9
ANRi8SOEVGGbGBsEAKssy6Y4fPS6mgLHF43jD4YV1e2yWVtJtPOplk+nEsVFfQXsX8K36DQ5uOou
GjjNIl4AhA/nMoXtM4DKoWLme9nC36M+n6meaoeYWzQmkvDfjcVDOoztAWJ12pTapHFss5bo98Fp
Ss3v1L3QLfw1KgIcFfgZCF8F1S7PzvBVh6dgE5MeoOVyvveEezn6lFdsNlxhOAPZk8VvhSTWbvhF
zaAr/AjU5Ct+6QyLkF5QY9E0GbgBW2A9Dx4AwxE3FlJbfzEu5MQrDC6C9bWSbaTCRZWItn7Bb720
b4YgmtNCyDV+cRJhNI+IhH1PWCJQIw7I4Vr78gnT4JMYGq0o7YD6fmybR4u+FTridUSReRlC9pqv
cAsI4gk3I5GImQOWiXnmA00WOa/0VeL8ms7fdrjLcFc3hHdc7L5ddYTNsFBZzj2dLjz6udbgcPug
3tx2kQFrkucM+nw/a9dK2Zk7yfCe4SLeIV/KDBCFpOIStkiM2aJW48JOPCtoRCDZuUaW5X4m6wDJ
1zjDWOYCDrvHJNz3KqVF3PJHrT9+CQJW81ssXQoD5iU/dwqgVR5Y/S5m3lC4oZPmdkidHVVfwkys
a4dBQVbkMjz91pWgYOg4wZgBNkPcmBU2QyBCqCADNt/PMW01Z3SISIWPQh5W+POoGMVtZR+aN7Zi
jKpFr9svxYiUuEQiLEFLd+4ftCmEwlkc4aJ0hssqe0rLdvoppOWw3eWbO/WaFDolhlVQR04tH23E
74svfCTgEhWEQg0szwfvJmeeQ3/C5/Os8L1EYCW6OUm0NlR5cNjytNbkco3RBOPbaCwBSWN4NhVH
+I8IXR64e4MdDBWAPSTaOaShXfuLettjYHTpGHIE5gwavoZvqwRowqB/86QcvCGFPilTBhChMTZN
gCTrrvDEep8DW0gjiIjFuOXQQZfpiigmxD35pP/zVlGc/KCMP0Nyi1M47MzQdWjuES2KPPh9vwnc
zUEflwrX29GZT4NkYkOlQBPn9zhAAaRzWJBDmQtskcWTpkY4Km05MPlMmkcyIcjNN8nPM7ekEZrT
/YDB13Ul7iImJMjHHBfOdhTmkHT4Civ4G/Mf6BtG/oTmOjUAWJIXv4sC1kohAbUeZJLeMu0NU4l7
y9xAp38N425GgAsuK3LI7ldcj9Xmqeyh5fLwP/7uUZD/YqsFmGbv4McmZtwNSnBfk/tvXHSWo30M
J5biVpUcqj9a3y5GgdaLMq7oHE7ivxJWLC8jHf/P74DPtUwLfkDFf8Ls5ULoajaljqNnrPSwdTiV
2t9y44NdjNUMCNxmgxAgbEAnQR1viVuFdYvZafc57EjtocrvXbTdjoPjufCUIyZcKneU475b7hh4
i6yNnCgpoSPqjykLqzdW9UWuCWPwAlChc3xBziUAn0r5jpg9o2caiE8v0KMw14cW+G9Y36tF+tE8
h6+N++OWiVpSdaf68t/WfY1nBJKPBtEelqupNwZeF5fQdxfKRSEl0jya9d0kb8tuW82WUPnc0TmZ
+FoR1U/hC8kZLd6VtybUJDkERDr6ZEg16/BXsHeueCEol87xxvhdLCTwdgdbn2XKsAINVxDilz4q
dTGUCWCghZV/XFs+mLMLwM0LHIC8pr7GXmp1+UnaeK6CwY9wHWN6uMrKEhAirFKAiarsLle0tZ4s
OnqF6H8biu2165zt4a/4Oi7I0gp5yhjem83EMSrudetv19GIFhsuAkleP0Z0cNsOuNZ8xkEKFPG2
VvyV0tkpkgLbf+v/m099ba2w2WkasQ5hmdqr6TuFAsJ++KcEC2r295cwdJe5gUT5QDGvcFkgE2t6
VJx33BZQmdyYmcmHMn+9yrLSEw3RfiSN/HD+F7f+flrASCZUMZx8aliUA/VIeKb49TrSGnmkqGA4
GqGqyr52ompBSnjPqrDw+e76WfiHZKK+22/X41GM+qtHX5hTDPVRHWH/a1mSVvYrgJyGgH2RrSz2
olTKYuWqGUgpfPkXvov0lKR8ZY1at6ExVgrN7S5BzIx0dqLWGWEy5IZbud1OoaIjHTjOuVwAdr21
uCZ6tsnlge3NKEoEofCX+cvmf7C3NwiV//JcH6AX0AC+8NlEdmM6V7NIvl+bUo8o5AFWbL+Y05mW
zmhVfocQvBcWdA9uDz6vKnH37TstagYvNV8zZ5fzaqybRXU9KQghb6zvhER6BHglNJqW7DbTTQQ0
wlTp4jE+00ZmYw/86DjuEww0BDjFhlwvGUBu5I40EQszg0kKX4hQhTTuBEH7+8cssAeeeSGm7X+U
vHfkuxAzJLX0yMLNdcGabS70S0MgRYelburIP9NE7caul92INj3O2o0QxdG1QnHDp8NAmQ3LbDIH
P0121f6VYgSI+g+rreci5LietrQCvjODelnWTDyOFoZUMZqzLWTxLT11GW91T+SCfM/czPswJCRR
CrXs6k069K0bdHQ0qh6NfVMHE3oPmUe9nEqYl0asYEgHUlk3OinK7fOgZl0xaL6IbMuuSUO+FAzp
YAOrSBjsqGUaoZ1R92RizS9nNmQC7Z1L7oNT54sEyZXp+penBsIIStOmKxLZdmjXASbMkhLuvUKa
ODaFSfJF0rcqy+qtEQqnIG4BHmcdNr25Xo99UGmpAr2Vx6/GqZSCrAi7/w97T5WEK4k0udFAlb4h
Ig7UqdwK0tfcPeSRNsGmkzcqryMT1BAyLGfpSToNQItfhWBczKalPA6CyNgDkUXDhCXkuH0fP1o+
lLipHT999waKi0vowehTpI/AakITqo4B3OjhANQRBu6x0kusfrd7YbYCc3R0bq0pqZn3594g3c3z
UdS0C8RsWN992e3USpIxvStWqG5Pz8QPmlZx56SccbwOH/JBInmuvpQtXwGQap4iRhcss/huA9ug
l22XutzGIUS/LsDhqF9onozU/uAzAKZNEzELo/B9twoZ+P41CR5ri3E=
`protect end_protected
