`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WZvujqDb5ENENvmww8S/ED6I3ZUXXxl2CFhATrysOELUHtxeLAmc372sospv4rrhlZ2hlBFVOEsVe07iNnbVSw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
POFzSez0h6HOaIEABoa7cw0rayatD3ZqG+SU6F+HXqYBgfPtKV6y5nHNMcfUwksZjWhTQbDyRMkrhoJkU8NlbA4ps7NvOPBL+T6XLgU3BKK7k3STYfk3GvlyTANHpyYUV07pP9FxEqDw6fFqzDRSFlmQuesnVpI6pFlv1bKyzB8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KeX/ahlrJclflHPZljdKMBl+2PIZFHlgGCGlXOwLHvaSunTOwU9hWhhEmFYr6QsdNtarPDj5TzU1qenUMzWNsI36w2okCaCbnU1HSoWdUnA8kW5Tr3CwqC46aW428xqxbogYo9xXGG66ZWqNHXAb0E2H/crP5Afm9+jnE3wZA8DypwuFCOTPt1uxBtDbv1t9dBoUafVz6aqBAcNnlgRv+aAU0EzqB4Nl1Wa/NvHZ7S9ZBdusVeiQl14f6P3JFyGVepsTM9qdf/fYHt172X2TreW3e/fgB/e/6H4p0og75e/hbQgKWOwc4uyKhhrPrrFFyG2seD9Uv08fXF7LKJs3Uw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gtn3utiIwTlsz7uZ7uW2GdmFrmtWwiFeEfFq3H8pJ6QqSIVY0AmLa9wB6VFNomq4C0gor46eAFDrPjE80rIQHeYrLV6o6S+jbJaHWFjqkdJVaB2EY5LxZJJmpBUA9bWByWn5Xpq+SPaep4iI9CoW7Pr8BhqE2E9CNXfyoHlw/Ig=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gJdpWQOUPCoenG8q8BbLRlFbLQvv6yW+En2OYg+dPEmIZwx3E29vCxOce18lGG/pwxObquE0583i9ZRHqCMfLo3KItcgZpk+Yvfa9OkGUZSb+3ZV57b5aF9Ne0/aE2Ii4XwDddwv+svxJv2EACJgby7tY5dvp3ub5h9qKB0P1UgvE+1n9yXA7HHFrL09Ki5+gN0VVoNdJm8OmDRPuFcfFMZlTFlGPpMOLRyomK9G8HNwS/Ol4PF7cGsd0Z9r8IDCY41MMYl1sE0C+NpL2ucmiaLrYqj7zbsoQ5lA92TbACIv2GQBmKp7b8scsIJncFjfqcrtP1o48JOfVZ/3u7liYg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 414026)
`protect data_block
kHzu8BShSQ7o2RBlA196Iwm5yIXTesuG6NxFh2mxWRbPVGUS96MbyVqYApnPYlGWMYssM2pR59Nb
M/HxuzelczBDfkMtJnUzP0sF0kAl/wPbQVUa0tk22wJdb/utYTINBBi6ZJ9loXbXsyeY4aeS7Hun
fgjawQ/148+ovAz1kGor9wdtkCGPsZQ3ufUqt+KrtGIPmdUWOyb3aa4kRnJsiZE5mO8LAirDYOe4
rbCkoc7rdDN2rTmyoGexO6BYVUyS3EzmCw25ZONwvptSrXXtOjcrPtefJr8WQwN0Ij03qatJujGc
t6XF65q5imaJyQ3lhcL4NStNYtfThz8XmR1SKgtubPgGZLcafkpKs566sPH+RQ1Rt75AdrTx34S8
EGI/BI4MHQfkL2RQMYrtuAPFGdR4608dC7xl0ouNR00Bf9TypvXNIBeD7fefEzfVwpLS9ryJT9pW
iqJicc0QTtD0lcA4WhTcj1Jf4ewenWJtDSSYS5jWNo5qt0lupSneBi0+KKbDvqK7EqHqOvaP5NH4
dGUF572WxM4Z7rqn8VfyoWEzFCdW9Yq5Um0tzcUmxAoi+Grh/e+Nd6VxOlasGXbk3m6qsmf79ymS
jyPg1A/Vqc3KwMKDYqsJ9301T+UuCVtcqeu2QL9aEjWnESeX9wZmDRbFJjCOiHj/9Rv8aJ00XqK0
M85l6/T3leH6qA5cZ3cwC51H0yokGqUJEzaGhUERd6gsvE//Yy7rxQH2IPuCMyiypscAhdlu51Ge
Owt8sGX6NctCSGsKfw5JfgGWHvZpVQMBXeg7B9xPwrdZ271w/pg4Rymqic//re2d617vr28iwEnv
Fcu0g1rQElqG1zm7F758J64DgRWa3D6CuXmgJLGTtLu/qgNHIgHAED/h/9XxddFHZNUKmhaOXB9v
rOqWAZ7fH35K6v5Ri+P7wnT+A8QtLgmShwj73H8av5OfL6XRZ+dLouDhqVYognulaqTX8ViCNWVs
J4U4PkGjAAKGBM7TinThOM6dHH33UQcl9LUGSfywsRsgSFOxc5fwC5LFg1HNUNeErh0DPBzMNQbG
JeZZfhANdlOSQXeuJESeGCVWBTdZfViTPHhNukTXfDNfG8eHaSOs00r40KP5ADs7mqBUa0TrCokv
ppvTMT7qKe0JwLwVGZFF+oN3rxToi+0cM9MhPd9ysX51OWHsVshIKguFFcsq2yfEAUr0kkFm+5tO
OKbfyx2eGCxUG602udqo2ZcM6DluHlovNT+wh1ackyU7IpHNM78Q9/ZQuckD+2C6/snn/nyYCmVD
PyweFyC4U3zJjt/C/PeI4h5OqhQTNAAyEaHM6/cRqcT9WfHozBN3rT7RDwvgqtbyk4+DHwdGsiwl
M6wH8p91M2FqpNj1GKGbtv5T2TQE9t6G0F1MeplXP8DpebFbQ/A3rADXlBnX9eSJhtZe8XXUrDOh
GqE5iAV3zghzlAWF7UzgZyqcnpIOUSH3dTYft8dsN2aCb4O2eybv0e47l7Lz4KIPY2/EFmDZvAUV
77YhFQOT/NncOEKy/KqVrFTFA4zJiGRvMpTmceXG2FO9jbE9zhqHRqH/Hm3zcvk+dLlTd0FEGR7Z
XU7aTjeeuw4pbMlci4kk3zfID1Z5xzIxXZmaePV0ejBKLuk6Y/+OkjNaKSbLGekn5ShmqwAemEdr
FYT5tPosR7iJKnOvmWkSMz6DMh9sWs76bA5b6VG+gFsqlMxsJRc2dHeHrOssGlM+UYh1/z9sfXBT
cC2mIh2j5UVwqtBvh+odMZ48igN87feZDVqZNCRnlt9rc8bsTqgig1+E6PHE+R2GTAECp9vKpfJ5
BmULWHx3KGBzFDsObssO4cgGUB2me+O5UfsSUHanZ2eJ7ekrXPFqRVkv6tlJqOTtqOnAeaIntjPu
7a7vhkrCikBlpoYzo7kZIRkPuAmNqHvlNdJiKtDpCjXAv6fYPoNkl8sElz7Bep6glruy+b/CALWG
IM+yMgqm6lIaZaeMRpSjjYKPJyWLJwKlnAiArlxyMO1yrlxmP2GV2mLBGTTVrkznot0UfD5ZZ7A0
d+hiaYdBUjBIuhHU/pGfd1RW4DW+iJBGmbMuxotzjvFXzKWk880KFwQrC+wHcaTZpqctAnJUEaHF
Pcwsw4Vsswyj1TsJyvKRjKu9KZyOI5eihGHZxNPBDtMaM1v4kcz1WUYKIfWvGBM7IdR5xP4x5ura
IJmrv4KAleBCeDzqc/hBY/1XJL77SFl8FL28jva4Avf51Ym/W/nluKt0uw3wUujO4BmwwyS88g8V
Uz9MfI4YP82wUxhuZhzmHl20tPzb7s9WnO4rxjoiA1DUwnI4WC/AWVlAVE/fS/Y+Tw36xUafQ3IM
ERYG81Km+N+Y0c1q1zyoHlz+bXWTxPXv+AAx2UsFSs7JwrIPmhGofOsklnTlIpRcJBbz6yUYINQ/
cIvWRUl5Y60pRlvKpxHUW1UllF25nwhIPUXIaEoQVc9kBhgJQGLAwOtz4kPbqAvILmQ8LFL3sgtf
q3deGmodehd+3E5dDGJbO2hP4PpwkHu0QYGqlzRBkHnAP2QnhlSDFRp4rphmqj8uVvKAN3FE+LxS
Tr9h9uozFYDJ3sCR4tobxNzUcxbPJVeG3uKglqHahCBtQgREtOiv4zb1F9Sbqvo6jSO2Y10WSykP
2ONlmf6MU4aUWQoSQrvISIEZWXCHRc+vADdhKSAOi7KMpNbpn3bD9mMnXiPoWEdhP698LkiFPKnE
/Ttwa/vAqJHT9QLqKcrKguaDgU4SbqJu3p/pfiJ7xIviYkaW1od7O9LkEInGZYVkkjtfnKDbaqQ6
GzxoLB+xlaUJy9J1ik7iQvt6OiKP88dP7chFgED14LAbbbUyEiJY0WZddVKZ5r8KLAzZSlPiRKk2
Ome8jEwuX3E/Rg3+wvSwitcU4w/m4198NiF46mYajxUJIXJ2cagl6MQCzgNxOUe7qwRqR1qQl5KY
ayRpRORFEF6dKBksCKnR02xjRqrjZxIEkXGlb51nS/fjQwmu4Q0dQh54rYgdpkeW6iU1qxEE9Yfs
QcHU6Nd1FGJLaSCKb+iIvl2ziRPvuTjQ2w39PCOGp0ZZTyVEOqjgzhTLYkjhvadsKotluDGblJTT
9Dz2YW82dZd70KXcYdhipk97qbpCNsVrwUf31RqDXiUt+fmwber2SOmBT+LsL6hnZDMtFRfajLCt
WHzSGjDsrYsP5hyJycxMAUeMSwlhcEYtCFdrCU/qHbVFl0qm9iZecySlxQ0SedsSE5xNg/zOVObF
iRgJ8OCWnHHHX6q+Made+cGncpJjR5XNKnIGNqcY4A/fQmh7u1saDZPMVQ2tPD8hORFzu4+W4WMp
cVqeaHqviMVR01E0fZEihD3/t5zLYlt1pc8nsTnYLzMeiEaa1CS25n0XFG4JxBJhqakT+40fXwyz
FC+at27xqPh9ZnBpf+T3GqkKkabMuRQjTbtk5reOMeovSbTjdOpy6ipKhehN4+tIEIzIXraCef3O
ngW2Xkirq4hqpiXltosfQTGK3syshoXEYpsb68HZTa6+pnya4Tggxw3AvuKJF+3UcHPUHsUVGEda
j0T2IrdXcsli6LC/JW+dvwNoloH5SnEwSbni/VrkRJcD9rog+uKuZIZ73elPelWElqc4IpWdDjv+
siNbsvMVDIkXn/3wz/E1wTWG0lZCfPKaxtGklr/iHpcZrCjQNiw2SrXPNviXjzV6TNFCdr+xzX1f
Xs36K8ECzpzcWR0ItIVE6ZhrxfudUJGtxzdg2tMnxPJAVM5V1GBNl2+jsu80vJHeM577CMWS1NDo
GBX/1Hwj2URx2nRCUX3sF+/SCEllMS6Yg0DsCd/ehRJDKUdtTAbjGGcan2T7pIeG9aIsbWGI0d2V
Qd5TI9nsarYXU9TwiryebF6++/TuPaFxepbfBS7yP7cWAsbrHYR2fqQUgxYnx9koXAkza60eshuh
8RAL/hs8vicM1wQFZMmQQW0SQPAZMACcFOi60l8eeKiZq+zABq+JAjlgMWEYQvZesU7PzKrB+SOz
0nF3RKSta/3hnPmiIlKJfgYxOe1gGwk04busKVxDBTVq9A4MnEJG9EpaRXxYPTo7ABcfYbRmf3kG
Nkk+NiWhCLsuoHAYw/9Oea1zl9z3OGYP500iAChlW59Iwytnvdg+oL99RRvZabAIrb2Nv6ved6a9
VjTcr1s9ZCfRUSgmXQn4XEC+QODiLsyWi6sdSvvZNUjqAsymk8VG3B8qQ4LZfZ8V/V6dn4PoSy0c
AHt1Jz8OMGO+ns3n08U8HMj7SgMoZ136EmweiY6NZB+6spq1uXggqWx+AlcEVKfTA5cGiSRE0Vop
T2BTamETlGHsRKWDK4szIGEsW29KRc7h8WbouGu540tfsFcQlpYj5TenjACLvskz3Ejx1p2CIFvu
kEjBajvtPUkEHM572oiw1gV1W8+xvi5qJ3yXFZBZ8rJRAZTiCOVplrOcN34ft1+tGaq8NOKF7HjL
+uuMnJWHMRKayNgjQLF1V35a0yoAWo5oQ193IyKPdtE+WcD2ovEFWe6YQGZtSx+1rIZWUkcT4qcg
r5QKnwC6yz3EFgv965CGY7M5bmUfVHV1ScDKn1kuzDrsXKThuGJX11UDAsXWQeNDn7ImjpSJ7pvY
nKitdaXs1iWIQE03WXU/8kE+mxjzJaoI54k1i6VKNu2DFIZEiqS7bVWHPT7DOZh0gf+lmI4mgIE6
urDZEdkRAF5LtoDDa91ttiywjyo718dGM5ccSyJOzpcZ+QcA8Zge/D7gA/Q5D8gRVlAxEw5CbOZD
eZSvPeT5zpXSRRobqqS0Nz1nnm2t8oUAmst8JBm1nLBI3VajgGs1x4Rw7VxYOS4MNNyksZdOkv3v
Ls6vzURqdmKgfGvZrOLsOrnUZW1Ay82ZauvMgJS5HY98HfxbQ4AGxmBoSCz4gn9StHuyw8xUgDuH
SPIxLbuOlpK+p0ved2/nKLYQ2NP0c3kiIUOKgSpUgJ3LlI1t6+OrtVyM3DPdGu2CsRZHdlsfZcOU
yOcM8CHJS8QqfFrBdkPeYa65OPufgDY+0ONlxV7Q7A+Rtiggue3uBzIzhS3J7bW3nEGWYxU8vQzX
GOPLzeCUWHK8ez+I1nF23IrAShGIhWP3Rw9uieLYxf3vJF+QYIB5np9S5Q3zseLPb+YCyU51sfyO
APNxl84kx8qi8X45K0rP1JwXvPSyng0MjW6KQeGfx+xJu0EDBx1zutgGLLdjkQsZQzpADfyLBBQW
9i75Pljw64MVhxEyW3lFxSpAInGKrIGdNIhqaNYfbYFnJOCXwcLJL09FB1FLNadfSt3PrGQEpStX
NT5IFJUMZeLxGPFdB+3UppJr5xhihJk7UR1KkmB0110AgCpxEcuv1e8tYogAeikx0rkAEF3NIC4m
2Ty5joMGp0AuULUacT033YHYB0WbSvCqb4dA8QKSkBuKh/jJLY2Nvk9lAQqRljBGLJznDVCZ5XEM
mmT4Kv+CzD9y07txn/FPyN6hptsRfZBnwbpyU41B0I9S7oELRiHQGWdcMU8MkfcbDw/+zdhsd/Vu
9bySClKLZZv5B2UvoMzHwm3GXd02QFKoCoFCSQszdRd9XO4tVA1QkfJbkdahTC9ZGK1IqU1ZTExC
e1EPSzoZP13IL/TPm4tJxhX0a8Jbv6kcmRajXEqT6GfP3msvjKkUI+pduUQk2iqOGHh9Z1n6aDe0
EIhaO4Gp/k5KjlgJ+NT12uDIaBGVTKwmpb7uU9oC5ZDgn9sjJ5imJ7e5Dw4nlZSvJ/l5FOT1k81M
eJ0eqY812ZY+DUkGpGQKzVwut6iOMER8/+iqM/5m8tZKxP3RSS64RT+iTqbOntvn+cyaRuGjp0qd
By4FR2EswCNBEMITgN5qS3GTHotj1x/v9Z5ssEhEVs62lD7Y7NRTUUheeyFv5RDvDFd59zFKOoJP
KT6GIfMA5xwrbXDgs69E6XAuTapErHWyFH1bukHJIUPC4CQ64dC53k/pFNMYs0qzEKX+Ma3iAz1E
wa3zaIUm9zPwEkXtWrgsE58UQhKjMCVdfos83rLF/Fk1K1qk72oNNXzJOAbIy3Ta6DFvtlhcdlBX
syNzLVhQ4CQA6XTgpDclB8d+2Q+dCOI4H/ChtcEphOMc1ovCZuRYkbCv/uSsqr8QR04XC7Lx0Svh
4RrC/5qykvnqIxmCol9GMW8AD809sdkgzLTammsQ2suNzst4DmgvM0AdXnvVZyUyhoGStlTptI4g
B70F+xC3fSWndt/z0x/QPkOdYulx061iNTIxuyEiCrWxzNYQZw0gpmXGmVkFYYoe3j5frW8e9Ppq
KebHvp6y8x6ZMPvwhma+gBcmihwNdvUQbbQuRWOvdo4SlC2QNnIKAtMLer2U4HuxEhQvuNSxjL0+
82VPZ1P4sFDd+aAl5VDIGjlkCuEErW2QqemSA9oA0BcLnGoqTdUkEgY7O2Z39Zt9nq84JA3x2Ao7
8Tj4nr3pROcs5ZPXEJUffSXdJyyhgEMDalc2fRb0K3Tz9Np1ZpaQ8hiHy0M/+l5DaicOgrv0I5Dp
93dGkFQR79buyLHvH5fQpdVZrq5W7vlOAtcAFAImX+N4MN1gKAUpIn2cEWd2brF8f+2wokq7E8Ci
ayYkuUbQ+cPdqExTfkxwgxY528g5BS1mflocnj1NoWb4Laf5nlouAvojecdjWW++kwcG5+DHFpo7
KJJIPJ5WOXMcJcgakbcKSCkLs3QFzP75UwDV+g224pdGVrEhVZHIkulooa5CbnzbwooBdT9Elp85
QZzyol2Ff6qy3+5lBPKANPqLjXmKiM9/RWVLxPeC2eKKB1QGKjvgo90p70Taaa5rBFEY6GR1sLP/
wQU6ZbmvPYGZmF1wy/1n5RiRvnI53J0HXFGlJos27TvMPK1Bnj4LR+EUElwbj/5kbaLMKC7ynma8
DBqi00PC8rPScx6Ai7MzxuNs1bRBPlJwqawI2MvqW/t3os8hBj/dem1J2gQn+4JdvH2zky/UdpFU
Gqh9CK67vYFgPdbosKjzzUo+DnnhZ466kbjAcvqXxVRwuRcZQ6+pERE3mGYHcbsbJZEQpc/5pdVR
6jtZQxMmvbsH0xiFmYHn/T2S65uGRXAwEYmzw4MfaitJ0AHP5K7X1g8XyeSwqRksdCYNCl2Oba6j
KmZERFKTsMADz2hvKuvFJx0qRoPpeHPLJF1muwi0h2ZGKZ6UuAolHYyyeN3Aqejo5ECQ0foTx6ja
Ihacw+ECkIHrZlqvRSiSlO6zVy0rGhkTUqd8skD1L4qDaQQCn7QEV5GUfwpWx7n7KPOD4WxifLje
L3IBZk5pyTALqJAh4YuA7kt9TxWrlC9uj9udKVqQt+Fzb/etXqwBOcJs3O9VUdeBxgDbi5MB7I7h
SvcVqLgnuSYs35mpoc2ex4sqvWGPN7amaol0aDiABvsGGqKVzZx+gPZBR47I7tTgiWttA1OxKmzX
byfPUGQb0KX86N3rFLG+DrRBXsfIYcnEGxeTg7AD1AOhWiKTOE+CKM/U5Z3owVO/p4tz6ITRIgAo
zvZE8dWuX7vs4qXzD5RHx8D89gTkHZtCfF8Wx/6dVAKpeYg0PcBWDCXlbMlo7abW4j4OT6/0PCS+
MaJ99R0zjhUq8ZIObqxOYLxL1HTgLVqE3TZOYJHFS+Iw8z1h13Cu30qFtTmre6q+B9cb+x974Mtn
8yG6Q96tXNPwZyB8z2OjTd2jsRKj6UfKkQehWLdcaVLXl4wjhax33csiJaSHnTuvVkfnmvDiaLtQ
mQONmTUCuRLBBNWS3UJzsWu7r+oXVq5eb9rHOZ1/TNS+9ouBy0L11OcJ/j4Xnhe6MfzKP7GAKMqx
yFaCVMFgz6Uh4MQaYwlcOzK+WLbVXWae3qEl1nRm5pFzmaqasmNety3CCTwe9TJQJmbsGfZHuCjz
B4+qht4geOz5QoTckc7kP5GpDHxawjoi50ovh0ZUlCDauW1gqJ8hpwFC3nokxDdhggPz+gP+Tkwb
XLpG61vrq4e7krEZfUaLmnGB1kE2AkfcpxR9hVfLszxxEmRV9fg+uvXA9MM0e8jMdqAftk8hy0ME
Cc7HQ9hch5nR9ui0iwa2ng68KFzknOdzOzFiJbZStHM3GOkBg2uVzB+j0LNn/ZDH2iHP3NuACiq0
Bir41/6K7MHuldf9b6JiXs/I0QVF5sj3hxoJJlWkNDcsHdO2kAdlcTU6UZmInF30uiIEpqPev6bz
347bu3cl7KzvJyA/ME2ASImIoKIUIUbOR766wOo3dFDPG+hWFdWnuoFkbjie5OtbsvvESiT2Yesv
DU5inJBO571XhyMH7oMlL6o1gJ3A2XiHs7RKlpQSeNmeAt2vuccUnUDQlGJbChJpBUEQPRY5TJxK
B7IqwZQS6/PdHKRjB9c7KaPq2LnyYueIjv3ip7Ca6E8fSWCy9Bz8q5/2iyNnZlBRxGgc4a6F7EeT
f89nHQrbIJ2fjaK9YTUKm1roRUAD3iZHuJuxOVkBAeNgc9XbVrWeDunUpyQDWHGiCXYyiu5A1FFN
Ht76vLOigZFdzrv+XqQmRQ3PvS3Aza3xhf0/NcuJvqG6Dk29TRE25IOXir3ib0/lXK4u/FAJK0ZA
+c+PVTWnFXtJFh2tZAZKurD2AEfFDyum5HoddbolVWOKK+XP01Z/O/cfNKL1+DVyz4oZXEo3go0b
U+34yC4IMOZTq4MH+BFmjr7V4AbGsEZwiTaCkE8THM0hll8X4QTR34D5nwUZJ1kHMBJMVPUQAUK2
CNkZwTgdIGZv4+CYMgu5HtgJqIOnj0KXk6gzYGfa2EBGKSTFUpYxebnS2QuYEz3mTpD+xHltqrPr
2KomlRLRsgCjbj3xTBDtOsReuCpEug6vzgMt74y5mb9kbXRws2Mh6vqD8eMUAg6+OoF/7Kjcijvw
2qCJTMZirGL+pn/uFZCGFLrsWpax7T8GTM+f8R8mbjDuSJy654Cxcm8jO/4QuSgzUxEhMlv8fxGE
fDf+/QBHn0h+yBqPrOQUsICcb/jnEOoq8UbB6oUlWak6aPYA/37xhwP3rAvZW8a1w6nlCiOmFqK2
l9Fuy7pexNMkW6g1wUvcAZdV/ZUgF41xtr9DShVM0xt4be3HhHZfl/pMypjhe6h0XfvuLtRofBGe
yXf1rgTpThhJRz8zheOTcJJt9XoWGFpKdgthnD++8tmry+XM1cL1ekYlNumSEPs87Y2O41q4BNXd
KE3mulfSma5jnyxdI3OPWx/jUzYyP0b0x5boMdDJFJl3OpmzFvPO9nTE/MBeiJBsHTeb5UXtGn+6
TwLl+OamTQptDdb3H9tcWHz+vPHNuk+vJPcXjYM+wQ5uR5sba3i6gvVEfxrRy7YQaXDPDGn/zqyh
hBWeUCdYGwJD5mbqavO1Q3gj1p5/DtufYOK9O67b5LMtZGCspBz8oMhBUmEKS0VCeKAR4Zx1ZsYd
lnAeXEqgYQmWUD0UcuzIJHg+eBBz0cxmKCwcvbfUZ9yHrLVqFuPKCfJS+SdJ4+/qu68MEXm5jrsF
XT1n3W2vQMt1HxhaY8KrU8wwgti7Q0YOhSzlBmZIMjRZAWaMDzdaZzPO5Z7jlIkvklzi2MK8+41X
9U8FtkAdD7cUW04EevN6BEAcqu5eT9MN+eLoxm9ZutY5ZePpXqt80PwJZd0qnBgkllOgfn+eHvBc
gLzO+sUpkk0je5YZ+TpAoJGBJROQrDE2FpgciS+p9zlWxeteip73lSkgJ87Q9JBscSPBhG+VBr6O
tJU+MeAlzgvWWyL9U21qQdFTUa2y9k0UVNP7a4TsIRkPYJSKuUOSI3bZrYtsw0Pam3z+yNr6Kmf/
3algtEEsIQCAiNwzD49JQUmz7719lW7/ihUXsrt6NCMGYQgTDQbhFR7meZOLad17wBGc3bb4NrMh
Zq9phFnMU3E1ZERPqSnPZJs1kucRFgDXNMsKiIE6VeN3fZ4AhfW/JdcVl6Iw159btGA9xaC0rrt8
Br27sK8nsF9OQJe6CZ3ql+5nxilFbAErEyq8g08XteIOfMuP53hBjs9qnxGETVOKJt4D5namVcG3
fdHWYePUcqFlNe1qs4uWsFH6tU5TuK2xZ6VBSku3R7fAX8/gs9n7CgpS6iDWG1tBAIe7FvkmdycV
jGO9J8TPC2QSYlptzwC2aZ1c9QcQqXbgdZaIwZnAdAFk0z6oSxC3ky9a72HrZIIZwpUENf5ZXDo6
jbkcaent62RB2Slj9RYaOBYj+H4mdKCpJh2YO5O5WLIA1kWzKodwQKlWFT6OfZxhaHk47Ocw9ClS
nRWRFeYRbvgwxQCXM8SaVFh62gT7NSDcQNtby/crD93F1rSLbdKCnp3Qvz3c+FWQcIZCOAB6MZ85
JNQJ8afRnhlQba/iXIADHISiWWGa0oiZtlOOqtELKZxyGMBU4iecKbacYQgDjrGg6q20zDOWfyia
DbYqKqEeEsatkhHtCy2ooqzP2bDJwxX3J8njRc3/wCCmglxYiPG427H5ndRuj0tNtDa8UBs850xc
Z4B0O+cqMTPiCQW+dNGSAGkOnuxY5RiyVoGUXm3ANeSMRYiOWAC8LJRNKCBRGww3v8FjiKNddsnL
G2mLxMTr246WU5TZ14iZbUi9rVtCkkFu8XwH/tgHx3JJWX73VLU1mqlT4ekqPEk9BAogsGjlviTf
I81FOiPqf62kj1BNf3FDIM83ylUPcdVPONjdkzx8rAEQxsUw5TdHJ3dtofxCqa0uqLKBvXxZqFib
srDTfgY/qQOIOBwGhMFAmcna7h5rV2Lr/SCFJEjAlMhDlaRGkMpSTj+1M4/O8e1lrRa12VyTqw4I
HQEFNKtyagHojvWWmMAZQKJGFZmnk48ql+1bycvjdXaPQ2x/R9OdNAwQnb7qm9WZ0HAOxQFosZlF
neIeYgA5GDfS1KXLoX/OeZYjEFHJOye6qMqmHwAeDsgwRcdan4IvKaS14LfpLxZxPS0apSmhrR8x
6CuQrvVTasr+hZ1avM2iKZqA7sfLbbpXu47P1DDEcDfptEh3TPBMkuygIuGTih6SP8dkV/2nSuUx
KQvLZoMbIu7BT0l1ft9SzTont9XTIlvbKN3sgvhIl44R2GU0DO101kzUdT/XmBvUnwTE+7mmPDiq
H5XTDY/mbiaKCQNGc891IPY4wBFsVrQEyBBu5nzUpLm3VH49dPXvZymC+xjywEn5JFZJ8vxnjtVL
u+o8jifoWKMAi8jDXGsZzniWLhQQC3kKRoveYh4lxthAqRtVnr+gp48KBD77rKtsjzfZQY9+ea97
0h1OPYwA91kwhWBHotrLuJ1i73UAjmJIhhyMl8skFlPgPEEeBRtlvupoZpmUN9eu31K2hqlP0Egi
azI200mvEMstd0ZSXi81PUedcJE0N/ZmS1K3e7gn6AiMlz324qYnml58Npt68SUN+4t/3nAng79b
3qmLTTuHr0pkO23JE+YAnond7s/BvHJMSAIATRLwxvuvVgaCj1p+kS0ikK31m1z3SN3SugGhAfGR
alsPPCZGEfmDWQVoXKsP7cihtbipGcgIobhFVOTMu8oG9umSdQKVOSN834Ryql03+2/IyewyB37H
v6YKmz3p/AMTc93ewSFyhCaGOaLpAnDtfWXNvEkBwTtyFRhURUdnefDAhB3a4KDHNzEDv+5QzRva
75ONho3V5nNOdqo8TeGGi6mBFQtTT5W9ReZ0Thi6v5L54vbnOoM/Q8jbCbPh8rZEtKe8U/AbUwnZ
qfhN7rqVbaNlw/VewJ0Gh3RI4vcBsvKYGp37D+jpiwfA7NT7PChrLaP9uHI0g5xrxh24VHiRs9sr
wCxUFXwa9M+ouydwt/HcqFLtcEXgComf+nkULdxahC4rcgzghwKho6R2zFkXdCgGxrw+8WWFF/fP
t114bTh5cKhbSPhoWwR+MKcygqKyRhfHo26Ve0iL62Gdk+5AwNrGByqDnHCHbuHP0/lyLF3xamSb
m7Z9LstYSqTxXTteOUw+yzfFGmtWYNerZAQmpOnhBTSWMy/Fv7hfy5rvoPcX4N8AfwBfD+5Epcmu
D89oI1KOkkQhgiIHWLked/ggNEcyyAEobVuModOdfwNNYoidMhzCI2b3ouxpSHemITwRq6ec2pSd
St53+nFdf6y41aiL+zrYb9tiDvb31LYLsv3NjbXF/dZ0W84dP/14H+61ogWCa0lMO5zGL9NBUCxm
3U7yoEAiSz4uTTOISAyIFdyJuWiIBdoaggOGYGeCOzs+UJPKkvGJ2lEMYKKozcZat21P40mL+Opm
icioG148/aeh6Sx+8DUSTnR6jyR2xtOqQ/qXEfwjyK0nFvwxFG5KiR6cznHT5U7ZM0Jm30uRSX18
8qTsm1zsclF6gCouarGuK2l3oMjFbXW9XYP4o/B3h2eqAqIOZ2pJ02k5+Q6F0qaNhhw/KcCQvCAH
gDJZrtdb5WzgJNagL+ODf2eimFUN4zO4UMbxdLXbIDZ0rsu9UCeltauqj52aoX+MTyzpBY85DsPa
httDA9SsgS/QZZpb9jap6GvY8xepOIzH/T92FKRvVj+dofejurUXpg0Y0rCaa/JAOtVHE3rGCH26
tR0CkiHef7thmKobNsm4HFd5rvvdMMANGdRz+Gi6SrZWHCv3Z8LxF3YxMzpLt4yRM6L5dayTWTs+
9xJ3qy4PHhNWcuQ5nF+62aTsunRdIh0rJ+iDRjAYXw5YSEpC8f7dAmXHQlx7ERQ51OgtnmFA8S+y
hiYvJ8s9s9z/hiehXWOL/QQS895OqC1h/XeDHjg29m6WjnZ/MQ8/J7Y7ixxwUzF2b3WndfSEb2le
a3AuLfaZq/T3IEEYFe4DfbNlVkQC4LwoMAPDlhrOzdcLXrxRUxL7Vm5FOgUhXfOPszazjb4jItpz
B4PSbv5zi4icupihGixb+JF4PjDyEz2MGv3qS5SMwix6mmEWOk1RlTEBsqca8ByAhqmz1LZx42kv
bFilWgcJVZpBK4u8QLwoIwG3KaGAMRQhbHGyfNivXG98oi3WglVVZ1gh1ez4uHsXIlg+wmkc9ItM
NQHfVxj4qoMMXBYi4y2ffyfadPxbmUvW8z4Tt42eili7tJBRbX+J88plfQFYGHGP3YxPa+Ooi5yP
2ZKBjRWhC9i5lpEZWfw/Ygcb1W3mjrXVigVt9uZ3HPXb/yiDOvSzcVRL+0tKCNpFvViVKk/PR0VS
BU5Ndm/pBE3H9iTPgpEDK0bHkH9OgcafhAf8n0G3RXeT97AuAMG9hAaCWH49yB/0Bf5eqVB0m/Qm
7LPEWMKl3RTBAcaTOOaXxbottBau/DE+Yax8TvGMhcEjEGeDzOs9bde5bmBDUEBM2/EInzv5Ov/Q
4hfyHLcu/O4K4Ehist/a9jKx/2B1etN++SUdH+HzoKnB7rdjuEj+RUEUZGGmsY6OaBj8S5bWaG9H
msIPGFSnBhzkaZkLyZdTGdfID/a3gURbZOpJDxVcVXsma/ifm7mfjIp6I3M3Asn/zPqHcTluPCxP
FulxTH2M+CC/D4LnuMDpZo5MfKfzsUV92eUgYPl5RIJy3jw2Efp+wAOo0qQMLGYLzV+Nu7puSAMo
QxqBugVy/n9R15A+1lUFhcUNX1VFbgVvUMYUjimDWLlSIfQMfSGAfKbmzzvB3c9Ba5bY+Ap+9SWx
1MfaTMGldQm59S4TJeHhvl9Q+GeIS3BaSt3rGtxI69Rqd2M2QsusKFBSepRi8a8Tth2X0rSDo2w0
LBpvK+INBkWDgqMihP4Wqlcm4+eYYrncden9qpRhMovSB6rBZA+gi7j043YsE1QLhRWn5ozvMnrD
5vPyvIS7VzVj5U3bmm/l2u81JvbleH6UB5Ygizr1TaoZMf75eaSWQl5Hi+tZIKAWM30vJugLvy0X
9Pk5HirFp2npfVBT27NmJJGRXfTMDvhXgxXtH6aAZId+noigGR8UafsytlG2EPOCarEvYoLex4LR
x9mUaFFxvfKRsr9Bne1LvLmS5BZfg7RVTid83RKE6b1FNlEDFzFknKRc4IxJroOBUJhUWp5ZF4HH
d/fC7FZXoe8L1/O8VCyPrFLaCgt5fHhC7lPFp5BxTbzOTNQBI4sNQsLRSd+poExV4bFjSnMt/kyg
psfS2HMws9ees4sOZhKaoXEia8uoIvU/sKQwFaeELllfPSCq995Atg23fkgGt/+UiOBo7NCKkNbp
VJ8BK22KQ2O1+oL7+zhBt0/KCgkz7/7MH6X4ifJn5AItZ86hnu/RSUXuKm1W/uCWXgaWLbfvcvAH
b9NiL+r5x4BKXmoGga0EfEYWoQY79DjtWO8t2jq6yXfrBqTE/HSJ9ZKyPyqtAwnMqIU4cLcIzEQg
vBBhF8oyPtjKngR2hxB5BRUIEZxkZ8P+PDhUvCxrGkEAawb4bfvQqbhRAXFMmoXLtPOanmq05U/2
ORQB77PDwmUYRpfLZx8lFdjQzE6LF8bxmOxzFu8LxZIDfckjqFw2VTBoD7fWTIBkXNaKvmjyCph0
7wUBly6cPncReOoR8tlVA5chvduY0aJuXmzm4Vn9CC6OGJ3/x1JSa+gDM1DDwCUmvNh31ptmdM5l
pIDG2KGZThfA/OhJZq2D8YuqjAG/XzF+pvqclJVCRgjRkaVQvJF21NXAsrk4kvFSwlmpwYrCVOCb
OaoYCp/9JOAYH5VTjHSMIEsMxWxrBAfXqza6z5wqFAlC5zFRp7sP7J5UuhDaI25CeU1C3LRXjc6h
YYD6RY3Qel7vWxsqAh8M4ehy9m9OPTvzYukzlDSwswfHtILZFo7KFnohOdCuShIHwVhwKGErhrEw
/kLgT4DVUJwgDtzUUIvjUO9q826++B3ujtxO6XksrIwyzFm7HjJizmlEQRSCuqKEgu5q2jzGGEBk
s0rJmHxEzolAnLytiQlNK37NIeQgh6mG9vFBfo709bidVc9a1bUyObyo0C5kVwZuBGjF0oj0Zh+9
fIGKaA+KNBoFYYKz5AXfTwbntmYzlt28NLEvbAovK/AJlPYy98SpkqzdjtIYEhoXJQgMLekOYi+b
gaXF95JL8Jgx/fqD6fSyTCF8HnBHyhDqtWaC6EPKjaLyK9BHkGpq7qG94zUpRlxYXZVUlyys3Hsa
ypl6SEMR3DlnEuAioQlzd5J2M9oasyi87i23LO5iO/gfsjhdbWSErhECiZGNZf0FQp4tt0Dmp3FE
pFLlfYFj9qKhx7P+l2z4ai7pRJS3BynNAvuWB8SHElRXcMvTJ45bu0GZvZ/8V/EpjNzfwWBXMz1j
XJCUk8GpBOjkXKOW5TLcJosQuEAiTdTenVLGhWWRHlDj3AVEaGvhzEZ0ymiSUSvbekmFUPIyC3Hg
XtB1Lal/gFg5iw7+TNaZL4iUVIspleB9xT6p71A1ywJbW9HjHVOyOUeHQjJJe+Iis2lWl215El1v
eqvDNoK0ujZo6XihPHoJnR5s77hMWDx5uE9aZW99vCDI3JvxTmDTwFn/xFDrvuFj+xJsK/wPOc3V
QtEgQOt/P33LQVD1ducZhR1bZBoeinQz8Mjr0bTSoL1M6z73B+IZWjxCn1VCdLndVSGrqUR9wNmh
+qlAbReGmLSBP/ab0txBuz8KQF2Sqb9sjLRBpM1Rai+Mbtg20QQg4/HZpIyWXKUFCsq0Wyjc9g5C
0ANf9v+V5V7wM8npWQHtn8nroEAWkxI0wYIZuDk6Kz3vMCspeV16dj72J2tsGxIktN237AL/p9Vm
bOIFZNFkjMTrc+PogSAqCrx6pRuiDQ1ZMX0XXitoj39XGNaIZfGLeLCw9EwDFY2fZGkWTJWIwjLP
p+vgWMTiYk2vYWztwk0mBtxG3Y2RoSRHLYy1anIQBTcRZajbDuDmHg4lOwhrf+gCCeW0PONXmA0y
bsTYkOzT+UeN9BX4JRsUjkQUvj6SS6Hrq3f3bxJdInzN0JJls7vLUZqjZadXeiOQWE5tCAZOu4LS
G1zbPzyLH9XvZt9Vv9zAz/zdMVTk1xvsTIPcrxcxUf/hVeCDsEnMkxCjw19w+4GZY5XfYk7J4jxD
x2G4k3+LHKgflbr0+mzIqs9Nb9LehEx3kpy/nH9EZFL2Wd9uaQ9RHQsJgRS+MHjCdWoE7vdgcxjt
nNQm733Zd0uHZ5CZnd2E4ony16XXGhY8wODpzRdqf6JGdbRRAK0zRUCjMpmmYyY1wcpyV09YCNGU
iDhci3yo8OTG1QI8rzqM54gz1K4qQd3i1RKlc50t8O+NVk3YKNVjPU1qemNaWy/kMowcICMfegAk
zfvv4WIWAW6e/2fjthaVObWHmGSa8iECUrZizOCx9EVpxoUTbHbPnoM7Vzi2b55JoQmyjKVncGHh
3bIgS9t0FlDfmMiJZspsO10CbTnPs4H6PEGoO6K3o8sdhbBQNBW7zC8e0YV7OXK390c6iJ0VHTy+
f1QCX8dYoqbgk7jbYfAsvNpS+uZW8EftkiS0n51+j8PNQSDYjc8HrbzyiCctxASg9zjA+CFiwPSB
GgQxxVVPNbaW8Z2eOcXrmsO/OC7uwvNjdUzY0cEy/WcSVTsSEsSv5BR8uilZLV4E7S0RccXBwoID
0UsmWrBB+noDS/EaN1nYoOpbAD8ur6wpJSx/2HJHszol2WlZ+eA9OQ6M154R55+mN4rHVQesOGc0
0FgLcKW+MIRknPhoTpYULKK4Lf4B2TuKY1pf+nwZtVwNHfHgmCNvpbFsxESVabcexcDGdocZZSxq
Jk3WpV6Axct4+MkLGuRY0pfvUroyxeF0LYElMLFULihKkVLvnk1A/KP8mM1TLOB0O0F0VztTtVpy
++YrXFp3Yum+LJQqE0iGSoFrsgwYYN9zTin/8WMlcMt0+N82nJmsqx7GggUTBKdXTfLwr9UsSNSb
H9D8YZEVYc0tvj0L3hIOc4wejlK0oy7biv1KBZQIXzG0kWLKIhwpH0sa7YGSs2KVgGnjHMQKmCD8
3CzurnYJ5qrzLQKj6zpFCiykMPc/+pniv/LIiMKJxbHy32JUlm7n2fKjTSW9c22N50lCuAup1wX/
23Cj8MfybDpA74Bt8BtKi0o9207jIGSUDMtn2hPCqq3XOf8MhGqGLsl0OQZRak/3BSHei2UeZrf5
ypQ+4np4YWV/qrcMCEfWBYSB8hYXLOO60NpgETnNlJ7FG3ZWSyqfImEln3WvLZzLccwW5ryU4FLl
5TBlNosDEh/9FHeg3VAWeesnWtIwpmQTuhAWEVDOx9FgY42gj5L7oOiTk6PhqYI1UQWd6MDot8jT
XsWPAXlTbYPeGhLgCUNy2nFALlMytFHbn86sxpmnTqtMbB3gtxuHMGVqVnQB7ioC+tAn5ukXLM9u
sF2/MjhRd3uLayMhNC2x2rWovsDt07Lwsh0N2bN7J+Ca0yMdg/SCbfFtHzVJHoyQv0sB41eFkWU6
blaJfyhTBOKQShyIosIGImWgNPtQMIN2EdA7MFZafGUg9ZDSfq+Ai1v9St6TvWEly5ORBoehbZtc
ddEFSZ+g4tCTzRPIeblX0Mil8MRCKo4O0Ij+a0mZTrL67DXetBZv8IlXqnjjYYwRVCQM58kjtqxr
mmH2bnOfjg9QVmahprVBVh8vhwGM2tpX//8CfmlGHE3nDeVMxPcHlTUVO6RTnvqOoLj8Kouj0Ek9
GPwTPJFzk3psK/Ddfu3NrU1Sc5lV2ABMTu6cBbMECbTAn/W4Jr9CUOXwG0/aWK8ZrR3TWGxT8lWQ
HLgv+GFi6r7WwISgtAvxCv5UuWFtoDhaMWVJh+Ws5n/lFwUhQ4vqbkUHSyzdaUsHybQs2Sl4eila
xkA/iJEK+Q27etQmRoLPs8iOb/Kp/fqAmil9yHwDPSFCjzIVA6qg1P8EVm/aSd1B89OKbeehZWND
IQAvYiz/0tRPod+uu36bDN7UCsbTkD4H2bOXbwpmwMO0EnwNdMPsnvRyUYedMq+dS0TLv52Kf0KJ
hGQfj6M82Ojgb+1IfJH+5BtFsOD8aiZx20M9ZRm8IkqzYIvIRF/jKkffGmKsJ98tBmWdchBmnfL/
uiblVHTigG/ukwhlrOagWep4rO6t94ljxQxnXlG63cVx3irp63cEbbYm7D0PslDbgpe6Rq5uwZ+n
qrjU5psfWkdS/T9FLXxMzgzASD5VADvncI4qOUMg7/6NE2DTBL4BhXGokRmYYmg5GmtqAkpzusp6
C1Hp95gmKrSONtLTPO/LvZ1SCUyf0Lejq3qgFi9O0Er4ha19Ns7X5WNF5USxTj5oXRAsrHafQluY
OkpD00kByuPTY/x62YiPabRdPn8NaTDowgNsZ5OEkd6jQ7SEzmwPFyeI9E4/YLNQ/B4m1b9ImwRk
HNcpiY+o9soIQuoULd/2+ueiLBBUcJT8t6t0fSsRTx8tNkb2xdazr9mefe5w2/oJrQfbbWps4pnm
lPpqovVeEARgb1qcgJk6kyjGq6hkEb8mNSOJjLCQfCgo3LDPR8hJo+rfbDt0sDWG9ROGcDRfbvho
WOF/hgPMK8/KEC7gDZBDrdFwF0vaCjogYq2/6pFKzxd2Qsq+rl9cjH2XvBKg7E5ZKQNz2zAk3vVs
SctbVMe2cfqnmtGa46z4gdQO9YETZq//+iqggO3IjQZ9OeSYt+gbyXl2J+sy3MnDOWEyNXcCBY0b
aSDqgRDrQL5TA+xsb3vYVnrYeagbXukVa132ssKg/tI+m/lXv40rgayexXQ3tBLQ1xzqN1biAk3S
5uYV2SAQJxPHpOj9kAe19K6dNrlMCKIW/9OBSiGjklIFSBtvmstZXoblUqzurLVYwCR+Ht4ie/Uv
Y/jMToIs1F1snxlBl99p1493YkgMtZZ0aV7KB1Rq0zWlDcL3XjtXRxogz9bINAYdFbtJqQ9zZqES
1DTUSiHA2euPPT4a20b+hRzMAPxmkm/3TxYAElVBCPBQHbQXbn7VyO+GFKc+TCK/p4WqbUwQOYNy
e86TcYjta1wJk/tEs1tZma38j9dOTi2GkJ/FWWkQzs/8qQwg097ZWlbjK6qzLmyGszN1SHkh8+aR
6YcFs2T1w3ZwqQEfTgJhy31ctMxIWTPOt6tGq8xSWupvxlqO5oMusaAcT+vL4qbZgsxm7UMgR21R
+uy7Tpra3CbQQXhVf95GO/pfrI3QfwwscyOGLFPUMhYJU1GnxOtQGRII/OR9seoJdrRvNU8gs8ee
DmnayuQqgnrsZxMHQucL2A8hVQL40HtIufUMp76xqqZOcipEtpIcEoD/SCUA6TJghedk1RHM0N4b
3TZgYbFl2LJNbuuLp/H1RnVD8h9RbWAFjrBfadTgFjbfN9kHkF0DnumTOaajQXHYgGgCjcEKq3Ns
Q8bNIj5oW0vsqQzbLlUAOZGaa9M5+YTHSNDBIY0DeoPjLcCF1IVmcWVQ4LBr6ftQcs3dNm9zcPTt
j8JXaN5reYnKlQWDJ3x+MHvj3VB+tdCKcm8sskPqmIh3pUQwvXkuFrvMJcQn8g8E8dK4GFVgj/FX
vD7Jqlpe/WVnrx7fe76FSozDhK9DRgxJszpnk5FO94/1UoXKd4afZG1n+bSYwlQkUO8vX7Y4fiBP
7GOZUZExk6D++LLDa+PTsKmpfGhw1WTIcn+l7DRGsrdVH0k/Yohx3oDkwrnBelgZFlArk8Ll5vVM
oIdYfAdrbgptYFzK9CBMPaq2IWOSE4vAKG8uBr1K/gHxLxns3l5IRY2FSe7epuDfBYnuPAJvhIzD
Q3+HGbZLkAymARWI/NKZhO2OGr6YMiqIAvrg/F8Uz29yFMLYKfHo/cMGWbBTxAbfmCVSjcmbOYe6
54Dlw+BJCOir22aL0VSw+oZPREeRn01T500W++zKfe1LkU1Rb36rT4wRXl+1vvXytHpiPCDCzS2b
Pt9YnS+z53oqwmedQmIKliNYnVk0CEgngQFUyFTuy8r723YlN54q8/c+3WBJJAaCHoV7pQoRgU9k
VVFvlliiazYs5bDOyEZyoWlSsFa3zIKqpZg/zbpOAuzfad5kRDlQShDxMlMj3hdXsLTAWLLWaeD5
BwXUC281OOna9VZIdBNcuDOWvluyw+0dHC9RYk/42oMsK7+SM/KpQwTyL15L9gnc4xaJFDfQHAlE
HLAlfpKiMlWPTFRd2NinehEVjFZnKINY3QkMIH+w4AP0MkXqovV01iz0BA6KTjBOotVfvKeIQ+og
LPlyxRorZ0BNe2bE0BLb9hOxxwM3UJlJ+Mn6o2CLxvTYpLButrcAw3+9/OuH3nFcvCRpTGQ4W277
R17JuD3otzypVNgkJKYedI3Hly/eqjZx5AJuOBVVWNxrvmW6U2C8c0IhRa36HVsvUke5/QrKvnrP
KF/KLMa3Vra7wUxPPSUjNwAVvIAP+kPf2Ez0W8a7emzCoB0g7AAN7DcZlg/1ycsIJNd+ZpUew/Nz
+0Be4+DsqPRuQTfr289L1LqfTQwNiOiqsCAFEpLVlBEhJMfG0B45Tn3JvUvRwjNXDOrHDa4R9zWp
Evyb50k7rW31DhtAaHBtCjHVnkOudt0G/KEnj4xucw/AoQ403xrWBbgUcDPgZaYscuiNv53728Y9
fuv7B8j9KwwqPQsEhb/ZAUKekmYIhPJKQIdxfUEta+vPyiF9YkFaa2od7WIDBRDZO7i+n63K06oU
Cke4IxLB6R12Fc2sJ4I4/OB+x3cRv61XsTblhG/xdA9DdQTG9JSyCPW2KIIMMJ57/qM0Sji+Fi1W
HNeocRAYP1CIzydDUKUlNO2694pABcQpQYMJH+ja/qpf5XtJGn0DaiLxTHIDKO852tnhf3kpNVa7
HDDdkIX94fyKMjg40lYfnK6RXwIl67BBO6wziMEhXdY0sF4PE0D2ZJzhXxENA9njl7U2ZA1+HyK7
ktvThTp/YJ2VXkFYkmTeNzqhswZ2adC7YjXz07HZE0wA85delbrQJFy4f2MNR5YtCoZ/arjNJPOJ
xZfqmwMJ01DbwBCglm6UKFXDXKe6XlDGp6spCNBMDg72KM75T/WcwS7byUZ77CtmBo3dK15jF/HH
JYI8UzDClj1nOrBIJ5YUpLlZF0LWuWx8MtReBrRFwry2t7Ke2Vg747aKZsWa+iX8xUGJ4Vv8Rtju
bazUMNmpCe1NVFde+q/0KzgoKYkHrct7x3VoUVIaF3wvmjEhIEjz0bSeGvjshgs2E/oNpfosF/m4
i++OtwOgS7ChVF5CwybuBJngl2m+scRLFnj4kD7RyIZ7KtZmQDavx5rNppI9HdyrcM4yofy4GsTE
uEhPOu4EDhCx0pFl1OBneF6Y7hPjdf81RXyz/eZ8/fbWI1RfeElGkJ0al+MSI1YlXtsM+z6dhu2r
9X8ij+BWF6+mmmR50qrUO3IokwGu0ZnntI3Vmyi2DqicXYNkXrNlsKT1HoHGCL1vC6Kggu8IGY+J
LJEXEj35ien6SZl+T2XQKajS5LS+O78e3wrBoW0agomB8U99d1HRo0zUL6NPgERc5io9oFmDrHir
7AgBVeGRTWTaaZ1CKMGFoQBDCiqVAldHFLlpdWuqnJx32opQznVWIsnUTub9fMoe7p6XpxqhJP9q
UfO/CMyG8usX5ddwPPcvSgfAQu1DMVz5/dE/GQd72hb7tRcQR3QEvP0vvae5mC/ZrG8h8lPtlW1v
DSOwcKQzgIRK/uPx7Sz47Siyq0N7q3RDJHKjSwR7aER4NmffN2lr2dIUyVpg/wuh1XHkD3KumqKE
H5KjVMeot2jaDBlnX4K+SF0wGh2//KaZE8ZhTsR0wkzXz/V0J3P0CzK5Akkqp7z/4/m4u9aP5O13
OzPigV5MyaWGdyVnJRRQk3KEkyUR+dLpOu0xuXJJicHwDnemhyB3xb1OC6jZpJsVhu+GQYp1yr3R
Qb976QjD5LjzTYeqCKvuv13b3BFjiJZLHKFuy6vB1c4bCx580XntrhT1PGv7CDIIPR19JuxbQwjT
QQiGfMsSqI3Hf+FLYeyl8EsRIxf1T/i2f38OSv8Keq1RkYodo4f0kuD2mIN5CaMcsfTSMKV0U3Y1
qkmAIgS0tWM4lEnu8rO2xTssQagetRilFwR6PxzUD5mc/saFkqvhx6ZtbWzeAklekuoSvAlQn8OV
OILmDPy7zkPrQHEdb+kyTx8qCtcz+KhEEhA/iuMtFOLyLFyKz9V3QNS4chP1q7dM3zgp3OEZ+6mE
2UR3Z5OU1F8zWjGbnTnVqQ2Zcdye/QSaBwe00vLqrJQH9npYZ7UfZOAu43+q+m0sW4p+RqVZfnub
1tS14MqbVd8rYVA00Bqxn+KplrmerjIINsJFSdc3EdJ+SueRjMZDOXwPPKRCZhCKUsSdcajkYqb6
1IUfpSTsR94MJuLQOP8A7LkOMfFFj4N6h4PQiCphS9AVpsRgxLm67QAHClAtc+7/A52TEgwxl7YR
XH5QBiE4eknzfzZrBe9FJaDdh8n8q1pzyHsAWIMTXyZV8J/JRpIjgqwAN5m39fReCBioaKruI4Mu
Oj49okv9nMmDX2Pkq2yO9DfQhT4KMZhxtiWVbWbUjV0FOpiRqxIpFJtfVSHZuYykab08qvrgvO2m
8NhcirZmNZQTLjPYGQ1BLKW0wQvMNaYsco/gX0Ako0czS4+EbPOLi7N+M/ZdlBidSQxxrWL1d+tO
VrdK8B9hSCDXwyhx8t1iEspecodpdIeIPxl/UFZsIqEi7lMBJ4qDebykb4CvnRRNS+XRTlfU5WWB
z8dIuvalXkM0SmkC+ewu5mXDl01FWL6y/XBxk6ovFQY8YMTicI90ek3avkFXav6whbYuUpJpsx5i
Sy5ANxXSs7pADsg7iyZPu8sUefSJufpkWw6Mp1Uc7Nh2xOteHxFyaeV+S/CujtbCtsNIhrsY7TLP
qZEXpp5WpPR6+IjWr3HxrlE4SU1AeAFjZ/KfQSeIn12VYQJslHPXR5Ge2BAA3B3gGycaM2AWNgIq
5OGmA7cRN2DQavrLsfqKfNwgY/xGWyO6yAiuQQAoasNsCySqKl2joS4Uz/Sb2I3ap2sny0FHAkft
LhuzgAyr+PgwFjVCbMpgI6A8G8dMEY6a28sfjiIb9VevkM0gga5sd5eFQifgrAC2bzC7tIqDr5fv
FwRoXWFRdtTLOe32NXfiuj1khFXCSdihnwNYWjr9K2BQ9tiaQKOMOYgaPRK9ERN4sImkrucVniVI
bYzNgR/2RFZe2rrQfUVl2CWogEErNSjd+i0uv5KIDdRSCwN4G2ppUA8GBgh1T1D+rJynaK0RIUPu
3Xy7Rk67JJ6lkbabLy7nWVs+s10PsM+f21Mg9qrjkyQ7MikdJYWQkjR5UGtWnqK7P/uaDrpoDy/g
dN3UypmV2qXu0Ll3834HMFb99eauiHz8MKVoyZ4fhIIHXgSYJN5Vfvu/+oRC12soIwla6D8WSB0m
vbqXnHYTE6OiTCuKCDAavF333Aen/M5zAWKpTHV8g4M4uDAxFHt/iyxatBtUg+GIly5vcjNZmPy5
u9QwQ97NuKH0SZjopngJm254NDp6r15uHY7DJhVu8PCqhUWg9Hu02MFyaUkamZ2i+Mp6TaEUBtgP
/3cdVgm2CCb3OswGIHAQrgGpFkmlav2h0E31RS2X115UtO8/2BEGqwCWiejHiucCGdyZ1WjdNwID
X5aMkszliXJy1tl3+/Ky3njHk/eSPLforLNEf2w6D9rh8gwvT49Fm1LWQtH98dI3P7ATxuoESuCD
1D3ghMfTgJaqVQzFNKb+06pbXpN2DrTQtVjC1cKflb/+2zAFqtTrOFfXKbZV9IByfrZ9ibf44FCC
wWTvUhBLj3khqqJSP5ZIpUCQJXKi5K6l1IzqDRiWHJSidHwOW9ba4kizIrf8Gl2WMl+34JzUZSE3
hChm4aUWcA+ihOMZM9xAGgm8jCS1bxaiGzP6Ah+tKkVNYx2Nhqrocqlk9Y7/uYbfwazTDqww38Ow
v255G/z4jx0m/imr2X7ee3HgY9+6EJxrmRgSTuSgC0eiixv5/0eTHV25z7lsnNC9iBPi33+EXmh6
CLYeJ+jHcB/avnWjFK0BBam0mDiSFpb9kD8YWpguGEpJke+W8tvlg0LlP8Qrg309GknQoImncVxG
W8HZy8BoPbJ6kuiI5C8nlitwpAJKkjQ3xaM75sF75kVrzeSEUytEDuo00ZL7Y3daw9qArDCrW/D+
+rcu8IhCuFtcWrar9qXrqonn9PONyHVyE3AwlZjmZYQWXmgZvV4Ekoa2H4JscCO1AsxZjxSOcDDD
br48L4BjlINuNImcM9nw73bDPH23CUa+3t3vdg5vPtK6//QF/OEqyKFW3TyCFI1rOEMChlSMgAR7
KBCsFXSLd53/YQW4x/bBavz1Rk+GIegXcnxnZMk+Xq0stdhvK78xTw7xFe8e2v6eRAflE6nuZs5c
rSx26Dz94mF4H8nVB+HXgN8WSeM/evy68eqm36MM5dag6pwoTZ3eSO3itFsRf1LeZvWlbquONF+Y
erW2uFxmAY56J0MSVCjTZB7oszyn3yRgKv+Nk3s1qsul1Z5QqJQjwDTQMxZwWDYSWJb3lDhc9Tzg
lYwI1/t75zhltO8DadJTcohqngUxtlVFYIzvVOr+zTLe4tkMXQ6YEKP3ZX/yFne40TutVeY5Y5gD
huN0UKE5VApDbJ3nwUjb4UG4+MaGjjBvWiwmk9XGf9oWGo1HETFkIBxNUxqRQGESkqJIzq/KPqkW
IttsXSTD0GTr6+BgqpKX49HPNIO4xSz13cfeqZKjn+mX+b05LRZ+GlgfD6fKpx1UhdX7ZV3dChWK
36ZeSADDnoGSYe9NRn6yLklxmIFDIMSnW1NQCaYk8B42mSk5X9E/LyNbOONAMb9nUlNTpxHfFz9l
FamrmlHyEqPfu/aWL1DcU4vqRZdzwkLVKrw3jDOTQnOWysX48//V4KPxO5UZURi09xFbk5c3diF4
Hah9EkDFPEvas0jbJpetQvII3YqfAV4wYtPb/JzrJUqef8k6syHVKukmqzDI3dUZE35qO8eTYu/l
9yUKgYmgZONOhazn8GqTHJz/CX5NLRFfsCQOfBGlG6efkoJQmpr4nmoMpZBoELW3sWIF7OsTo1Aj
u/7uEwpWvwR0lzfE5mjUx3kIW/T3APDmCsxfjWXEvfjPpGJwAstTqDASx0zowHeulSaOthUnaRRj
MQ7lhwkMMYkZNyc3FpchV36F+nWoMLcpL9awOGmepBbAucmoBwOjFKwy48MsyLVQhNow3r+Qqyub
bi+RWNRxBmGApFLmgFLonN4vhbQSty06sXtS7BZ26/whlOj4O1mmUKLbbHSz2WOft5/Pt5jrxup4
qFM+fhiYDKDWmg+LbQvgJY8944BT7I5HVgCjWtX4aNo++orSzQuDKw2xUDHahZF3rU5+rfUA/dmN
r/ZKjT9NU2KSaI8V4yrE7xiC1Ppb1v5Yz/rLlk1mQRnTM9tSiAGLaKiQS9UR/DRtQlyZuj40nIMs
ZAzeMYLBiHCBsl9O9YcNpQdqWbbASJUc2vuSU6OyGJ2arW+Uifj43KZHooZF+6u7unC22MP4Dcnd
kspQ8GUwhWFQUAigfrO9HNGk8gDZHzpLJjbLhyrudD8YgKHRGByvGrXNzlP3+RepwrtG5uLZEiCA
8g/FizZmELezovGrXHPDYcMa20fFu7USoPlvU7pMU43ffsnJfIwynvD9LAGmosAUbzoQHdCH4LSk
xpsG5SUn3rJ5/N7Fn1QzIJPaiE/1v19PU5ZR9MU1K6JheGRVcTY4vt4Din+0K0Qpzn5E9XCoSG0p
cca062c4g9kgo9qmLQ8QYebnEph7Toi+d30pR7iZq4sxPQ83W3eRt5nmGx4PoWI8KajwCiX62lnW
PGA5/t8+QiAOLnuLQuyONZ2XgMH8XLBUC43JjJAZPXG7E99kCCpXWl7NFU83HJVXK10kLrhX7GhB
B1EgBLjst0sxGhlm8tR4kcIgIXoNGJ6Y6vgAESPKbqbOOZoyZLZ/C81zTLJ1Fy71CMEbAFZBOm6J
8lNJkQH7xrAlrPHRTMLQhKzUZ9f3sm+6JMMFLdZuQx8ggahxQVFjXObsIG1u1Cco+ZvQkpfCX0cj
k8+JHQ22RZg3BqJ3bi17TBEzj2dUewta69KDNQZ0vcFh1pA6dbvPmNdDGkRvCjX9VGDsquM2fPEO
D2XVHcnhY8GYl6jRIF0PQiV/5eyjlR9e1G0GekrAV/AVzWjz6hBQgqjbIy1p3FFEy/J6ydVSaA2m
zwf7WII5nChC3OlrN+9svpdPypVuSPTXCFsDVEHZM5XLiqAgQzYaAUOjWRDKc+nptBdCbDtxHHPt
ivFjhvBM/1nic4Ta0KSuqiD9t/yfYZdv5Wkmgx66Do7jhH0gckE6C9Fiticyv+lGS+eRkEOBuVYl
0AKQysyNEpZIsYEJbhPwTPYaGONq+oB/V+PU6uNQWPmak1QT8GZQKhAWTdb3bR/StXvSMIY03hdv
C0Y1YOAOV9Cd8I+BTEZvPSuoldI1IUXkmyXiAG9YQMP7Nqarbj3kjosTGNZAEEv1WRxHilJ0BBFz
prlU4dUuRCDmu10MtkWWOjjNqvL8svj76vL0KgX/LzqmeSg2EoWSVnu6c3CNWv/NZiEcQuM4/4FN
AOQFAcmGPuk3NgLiaug9xmP3Ew3vGQrbkQL9oBXE7ca98TUdATJrpFC3Jwh5Rd86R/0bBtQk16Ec
ONJeBgk07ZcvkZpJg9JaRCxd1PNcCEynRHYjyj7sL8ig7rPp+5O2LvOKaziUU0egQot6qwzTR0sL
RPftTRAHefek1qUUAA/j3/WhmGz7q48N8KLqynR8oOBrlxcPtF4xJh0dE3gEvVU7oXoEnzK5hTMJ
//UqhvdYaN4i8kfX3wC2cdKEhFsNL4O1K8EuJzE7W8X6ZJyovvfWrYEl9kzBPd1Vz3JBT6YelHaP
8NfAFeVuEYMzkTXHkI+ZJPrgEHtdYS4JmkiirguL94shsn+erThyU3/0xsIQZqm0WhvwiMCiJZOh
HDm1yjJwePh10xwL8I2CwdeD7rducDhapsA1mNdBFnId9Sg3VciCzVVxscMdNC2qPNoxQ0R1rx6H
eUyZbApsN71eyj2/wrhxtdH105mRxUY5jWt5oDpuZLaJO+dHZvaQ1WwjigBHeFDLmBk55UNgS49s
Gz44XRvChmaG12Qcm/3+no4L2Ffq544czvz1YOiz6y/bqbgVW+ffabhiAbyvN54wOfkQmVagj5U8
X9n3vawew+1SLtTfTF1ODFruEMmo7o+pVP714wFTzTaNyQ7ng9KvL6EA8/PT8R3GdHdjAy7QE78T
58GUR8+Opum6Fx/++rDzG6fhnIKFvV6HzU+gPL10kpufP8Ma0c2++k8nPd98bvxMQjwF/SNjg/XH
qKHrkGIflp/ldD2wyoYxbyWSMq6xAg5qHJYlKsiabrEterUm9CtW8DE2DRgkjH/RrEdgCNKDTluD
3AKANhDGdA4x5W8bscOq3J2xtLU73Q5IaFqYeXtcp6iSuA1rJl1Rrg5TDckJVZtkznbHG8z6IM1J
cG2OtyhiIHBuHHzuFgNwX8XoZZzU6stz7D9FbYPYwf752/RL2BkdU74L0MSVhwCfK9ibnTYRyLXw
U4c6i7cPdwIphP6z3mfPYm7vtwBGyp4svdhss8RU+x35k3Txllg5ZDnwZPcTzOkBWShXjQjGZ4+k
uVw4xKi4rwYDhdKgl3gOfIyPg8j1ijIiWJZYCbIOPmqN/5ixjVIAvvsLWQfJixuWn1FiIT3nShEk
f4EYecVNO7BxQoEFNUUomrZROiUaWMmuXp7LNGKrDzFVBNOPhwHNcAW9hnVvMa1h9RlqF8julIXG
Y1EPjNg/RCuB0rQ6nnoGlX86O9IQ3EgWTdJIX9p0iBMc85v8os2aczs67xRcEnMv4qX5z6RWsZtU
R++ollgbRzK1vuSnD1GaqQ2jWu/RrsQyi756kFCq860bRAHBMRXaIonTVGQYs1ZD8CaZVvHRMbTX
GjLzZbETtUWj7MsrnYyzZjaaRgP1Yv/d4jEQ2/MKpsBj7WTZ5l+movnpk3GP8BKKI2IACLv40uRF
zY05viK8VhGPjqJ1xcLO81GeNUfgLddGWJgiLEIPkqhZtInVZVbbb9F7DMLytO5WJw8A09PZaqYP
3PhELuJ8uDM7qTm2Lr7HM5Po6g0nQsK6qaraklLX2UCiw8kraZVDK2frBEl0Tb1f12VbPXFDig63
XwPzybUpapMLuoDEjq8HM0l1O5YLFJFOYXmCD5oZuqf4kjW1AnzgITW8OtrcDUbMo2eYIwTeM5NY
0nDbwyfkkOwiA7/QqKqig/Wdpxi5rKLhRRb8uY1tp2/zern+r5ZapH9YG5/+KROjpkFSsE84wjIh
b3XvN4KFFeweI+iz7UXq/ZUQ1QLdOOCYeQTK4qilscnNFPIIHMDBc0aGe9Rk5x2l5W8AQab/psjD
vi4x9k5oWzey+ekHK+CS2+fKvm7LlRjRkt8uJSHrEas/qVtIXLQYGuoqFdTlOAnX1+xPeNfOwKo2
jMNydyBbpUIu+VoIqaoJ415WukWoe0DzeoE1yT05cOISHJIpC9PW6Kh5RxqtFEmp0nrRuuNQC9Ic
FN7a3kk1oDFz9/j66iLp9/ZW618WMBRpu1Ve7kWzgAIF/GEb1VH0i79w30ekOIH5qkhFbnltCKeu
fRankCszRVkPnYBDts3mHjg4Y1agrhetnl/hu11lQhgZeNXoqMlNygl2KHz4dlSCLZ0hP0FGb4cE
c068CHgk8Sv8+g0l3tIwAZMdUds48MrQjso44v78Qb+fEJfMcCYPh8gv+oCE3NH7LKnK4W/EitZX
dIGmOzr/11lp4IunaWmyrL6boQpRJUyRnWd/jeN0dX0e0tM1abWmfdbW1OZBgHsMyz4d/rfJU2ph
7O5SyAgrXz6Ry1SqgLnumY3XIeMz9LFQ0GClyxY+C+QepY5YIQFcjfYSxrw0A5TWEjHxmFQOPjm8
Nv6o1t9pQUFA9PbzuRUFReZJt6XCfPg+AXf8yUPpHGdf4SqZoAwyZnZF+3VKVpmB+Rlzdl4uQ+N3
IV5VUKnI0t9Yim3ddIulppLOjx6vfoLE5J+oeNS0coLWunJ7ay9LZaiZA4v5judhwoU3zKacjSIS
3OoXo+kZ2ZpugnOMzOQhI/Nwji77nlUxdPVQtOHEBL3surpYe+Kbt/68MDdxVIH7oIKQnmidhrJq
hCc3vh8eBGc2XVkUIES0AVYW6OrYUOq2fkRfRn8++6fQzBKtNaPzUGJLaHWP4+XGfCdsu+D6Rf9l
zbIcCgizCZq7XKUW6aHT1dn+qpLycUdFdaaqxI6/FLuyLB5w0hI4F/QWl08DmQoA9F7wLUjJkzd+
1UuX0ZMZMx8PmFJQFJk7o9FsfX04A680vygJNa9PfVFUKSTisUKjfnsodXxw+XA5Ipw2sUhZ7E2a
cqInBfvaN/MAx52i89+5723pLRTweOU872Ks8mWdCzOdX2YKIrVa8Wi3Kf9x3/DdGLG57cBDQ6+D
fXlP9q1l7+LtrjI/mESbz/ltbzi7WUIEOufvbf2u2I4/YI1fPbWAEtS6jVllbw2LZZOv+M58eVpM
SiGAJ5Aww2cW7SEI3SFWcWCTeBYpfFS0I5X38LSj6RsAhp49kK/oUcvDBBXH3Ot7Zv0zdIocKGzV
vED55vUFRZR0bfiAeNBoeKyg4EU48Wl6LXsEhfDvqgN71ZWZ/HddpB8IWVRdM+gxYvYt91Rh4iJB
al5K782+YaAnn3vwDMenma6ymATR7EJ05eZRT8mH2DF+mpnusZSko9tXbwnOw1Rw3sul5i1KwtTQ
NlJsF/JECbqD7ww2WENsd65Z4BTURp15k2JY/mhkv60dBLzCJH2P35FEJ2zrIj9SWTujgy5105Uf
OuD/0gz/e0GS69ukmB/vCBjffJeuLryikIw7+JVtpbcZA5ReuoIW4MeapZxyfmBbFmEo9RBLMCA+
0qDCtDuYeAuhbrvVMZZ7Wm8CozI0O0m/HFWUL04NNgkhYY9UiS6tCbCE4WQWpQa4zRz4qRl1EHkP
OPWCig6+aPelpOZEjbAqpCiqAeWmcC9KHAQHDAWLVASPqzEGF+VHw+WGLX49HKfkZmTxFikMHpLk
pnoGQCBt+dwGLSdOgbqlQG1UhXmAxjdRn+c4MAEQxvJ0qrQ+mKMI9spGEuaYi+oyhjzijyeZdb7n
bzDU5fprBMOiryGC/zT+hswj+bA4qs4YtLvRC7TfriampvrmRHWuP+5wubVZmNSP1rDep9bsHmWD
rYcJmBgeKYuoqSvqlURpOBYtIRDMuJ+eWrqeI08p6SlSVaTm3sVn38Me3UX7xowfiUfnRal1UBaC
h2oJ9vyfqu173aIl+xVYN0WN88krWbEZGAhN5OYkiXsDHl8YNWrYbETH+r6kS9sTQhV69B/Q4Nty
q0tn8LFFuQ8A/oBwBS552iZmea//uvFKXJDb08+uzFvkTD6tedIKTKGP1vWy6cxVZ38ewNxL+Jo8
A54THcfBLMdUJE7lj1WzpInClDBPIZNGRNiPVMWw5HMKIVT+IRx8oAgwJB5IrzWHmJbdTVMMLmk4
msQRK+fx5zXYSBrBA4iFRZQLY9+ndV4H6PN1miyvPpKyEcts4GHogKNy0SOEJTbRgqXJPYoEc4Yi
fd3E3BYsdUXUu6sQaCziNb6FZ8PEMmOhzhaWcmJOj6yqC0Mf4qjp28HvnNrQ4pubyDX+swzOtfyt
pErjinsP+MxOXGzM+5EM0I1t+vq20TdfrhD81hF8GTmVkUTudKliAEIMz/70Vj7T0o16YVv/H6aM
kBkX4k7pBxl/LtHHqZ802WmLJVt7sF8iGGT6bXRhR1xYhrjHQSwrrEtDxOHW+8FafBRYnibx9e77
brlx18eYjuAMLMer6Sk9urhaqi/KAzVtg9aG+DQQOXMG5JQ1SCOPCRikdUwQEzgrFqNcyifgJPeg
pnQ3DlxxnxqwST7z9K7qXsOF9R5L6sYZQCfTuqjfTGEgaVLCY1GwuG06ERxqbG/M+YmoPNzDqgEm
l8Dhj7YwSVkc61eFyEzDlPOULxod5lfBAUy5TaCZASq2+FJb98sHjKoV+uGq0H812fNYm4unJIFk
5iRwZkRwgQHuEEAwjwswMj9lcE06e8KFFvMDRTAIeVBskBt+8cQeQIDIsmy0g8FthauGWeTnlwA9
os5XqCfWTMnkqwzKqYLme09hylpsJc9Qad40fXonainC7MecXPKkseKkrBgwpkfITycTrf/fkvqy
Icdr8h1rJTSKSP0ctLbzyvhR0jMD0zwmgJoOmHkOpmEe6D8cHAuwVP7i6ylrOh9fvwHPbreyVTTe
RD531XhGyo3Z89Zu4BQX196AC2Q9h0+Y+fR48AS5Xap3aTAdetoLGAekRkQByG69QO7sUym7kA5u
20GrFMjCja0+TyVy8C6NPs6KOBZRElVD2/ed1zYQ7lsWbayvz4I3aeNirxihhWLC7oGFfA8nxscE
7iImsEr3g0TgCCoD1K8HNjxOaFrw9PWNaNcSzySfJym7oz9d8FvtN/pz8ptpiPQSrnims3p5JPQQ
4pxPULtngMuQ0qmzsyzgCrhNBqMXg/iJzbO+QKbL9mt7qlkFsblPg8esU9cFUpPWrPICTNKRoHuR
M0QpcoKYIFecb7BazwhSwbOFe89D8MKlzVAi8o9Q5rCwhvmncSVUzsrD5sVv9xhv8o/BeosrDK0W
0QHTic7iWYVaeJNm7bPRMt5YkzSy99TncNh+9H/TTAbu7bR9UFj3ml0w8wgm/trnHa5sn55sLy0D
MMr6zJ2Ulh1P2sCRK8r9q50onzx5wNAeOs+UxfATLCM1+fJHo89j31ywr0Fxe3sGyFWzwSEujTbv
N4daVj93wlfDzGSrHsvsppLQAc27jTgo1JP/8GPduYuC1NkTUAYnWzgH8/0WfQazQDa3wqBaku2r
s0cWyPFHqEh2OZIZb+JHiyCXkrlqep30Q31oUH7HEUDIEz9lnVf7vvOEPdlZbFJ8KAgFLVzlFKv3
94BuLM2IYqf/xH/YqPUOSw/7um1ydilr29n8y1Qzw5w8MLvrZ2jk/1ameyqQtgI9rc4J57EdpZhN
lu+PP8mlG9JhzzCfmCPA20JoJpYShPSQ4RVM6FlIZXwmxdQ8da/sEWT5VxNM0dD/OpjdvLRApcj2
eKug/tUxn3iwjyLazRuAX7DBxS/+kSSg1awBwfWP/wUqW12e1/1+wYIveEdi/lhUcDHyhZmPaHeD
M0xi3n0S8XnPzvoh61SaYb4wEaSmAQHG9Zjm3oII9TY4FArdD85r96q90MGo5xGu0syolr1Zq1a+
JAWnyjRbRSYH56Nl9d1MRog0YzYUDsjfM2sKnGD+0S7zomiprGrDFMRpzXX4zUXe7KHlPk7xWLyw
L8G2WR6u7hcgA7W1qHKT05mtc5ZhzvMkYrCwy6IG5WiV+RRQYpfv0Ut+hchAG5ZDQB10t7DZUWIZ
fS2QoBGBH+4SAGnUOSkI7UdAXcuwFUQt+4E9Ng9m5WvraIkHVceAIjlx9kiAfsB6IqFMK3MAjFwS
9/j8AARiqA9L65A56/4ldx8yCSugiGCqQhpebhl06vFqbEK7RMDOWQ3KBDivQPM1YsFoMKtqxtvg
U2PydT1tYHsRfZ0kUvC7Z+9lfwBJmWwDBmYu69cpiKShG2+OjDUuSnAuciNHuH4F/pnX6gK92un2
8tzwUw8g/Y9NLYM3EenU+aSHK6N6xJObYP2Td7ADa6t0cDH3GwGkmv/7VorDAmy50oQNiTukqBJC
oW7ia1f5nbUvisLk3soQ1VVdZWIVbfWpdSxFqJvhhUzGjrG99qe+6GTzZxdTXvTpqmuJNaZp5016
1+9kggkvG2yH7rkVl/JcfXcLfkEVVibTDE4QOz3188ZxLO+kol5HZ7416ETnKP3YDe5Y4zGVihcR
2dTb7RWe+lUkFEN3lJAPmFzNJIFEYDqryOYtoO/uHtXNQc/LdoS0G7gPLSMeizbxjL8NQN06Qf9V
qotZK8NoYbMfga+axKmA2PUYlHrkvOQcpB6qW1GfDe5KTuRN/FrAzJtO8puK9ssDXbaP0V65PkCe
C7Mvfolm6h25O3CFREdvT4UC+uyEgF8j0E/olZOMqLR/ZyihYjgCe4Jya/1sxj7XB45vruXb9O3k
fnk6YT78/6EbTxtzQgVTtxyQ8ioBslIC0PyABswPwtbKq6jrM44DCSVB4W0MDsrZ4p0Pu6LUkJc3
1lP9Kk3pnPABUG2aAr+wyBp72DcuNyDNj9Gl2ZDLo8r9VBCYMfuEpsO1nBf2Ud9bgjlRym3+prYj
ANDum717Q9jP0p5lYC++0Uzh9d1RF6ogOyel16T2DltupBbehwT78QrLUIYPwsZIi3CrT1qrCJoR
dOgPDrFn/sZJXTu8HZrF39tUKp2A3Bn7U1ZVlm+WdL964OPOvvQo86KjBImCQB04BygkS4MeB2w0
waD6iPxUTNvvoEpxAo4MYDTfMA3zz92CV5yFua6AeOTwnpETSexfUXmTEoKMSoq+laclnLRh/drV
lgRfkArmIFTecNvuahf5afqVgkO28hAm+WTYB5w7fxOeNtmjjjHAuOI8p7i3aDSYl3szq7KmNVM+
A9H1OM7PG053myAizCvdeLOYQ7t1AbbxW5McxE2SndA7BHEv+fXNFcCu2jqMMk/VWIgMc7sh50pR
YEc2i9njC3Qcrk4ZmWG6RXbr7x1GrLOrJPrTtZQsM2W0xaUmNkP3NrcR3pS5x33HtbN83ti9yHH2
M+fLkbgm6Vuuq50uhCRA/hL8TBOGSxGX8jrXuJO8xKAgFRPkUscvkIXkES253DLAn+Ke9Np8myz1
DMRtW0Blf7ujWXnk/QPVdTd8yjWSScuZu3pHmxmOamkabt7ZZies5P4jgn26Bd73kxKa47nllUkG
3Z9XTIzp0vJmJI5UTleY3cOYn8BZFmAAr4uCv8/cKcyix49Teb0B/3qOa/KP1mNSr5sIoFNTHW4D
4ynIln/I1sRvNuF9MWUGHKw+Dd+WNEYJMyS8funiIgbEIO5XhMkiaM5ol7VsPuGk83A1GBXXQga0
DxlYdhvpHWItaKiusNg7zdtDQCOElpC9AplK2fbN2BSXJkSIqPNse6+0bpLfKJl/ecFWnfjL6x5J
VTz6n+J1bIqPk6yxzuXOh3kG77axJ0n2JkKIddq5E0E23Sgb/Yz6LBiosA6xFGdeYKEhHDBYDPQ2
iq+ytza36fMqbICXYf80YTvBtot9to+C8KlBBMoaoWV3x/PrQHkorZSUEZRhWvKhRfecImWtc3l+
P0yVbIbJZiP9MojIJQeuDqI+S9vSXHbZPPYh6d1Cuelhj9EF/Z02KcHQfMJqkZgMCV+o/q12vifK
6aDXD8Dka7bx8yy0LLUCpVPxDRmYYUGrpRnaX0l2E1UqRsR1PQZjvJHPk2a4z4QbD7BCR/2gb5XB
ysWBNOh3Q9v5Z+6sGGQn19jwamRSXtEGWAm0/RiYeoNfQfDcBVezvOL86gQblaU7jSNH6g4w/Laa
L0nbUoIV9lt8lt+ePvIa3fkQWGbqYBiX/O/AKBBVBzgIh943kRunlolyt/eeI+2WyullZaGw/u6w
EOCwP5LspMyvNRov6dF6rDHRuN+9JfF6TSqzZ+Nh0l0erxef0FTsCrPi9a8C+ZP35mGH+kvIoi81
76YDNucAj3YGZ4WCrzNs19svvcHQcSa4+YKFZAswNs96eRsorTu6+FlYmsdi+KEiF82GYvb7XTfS
1WX6wqtX72rAMYZ6ra4xDzjvkOxBFL/NQlkmS5AVKGZuwieW6q/FIwZFQhjnKc6J1q7Svhk0SVQM
13KSpQ8q5jzpr6Y4NRWEpOAKo570p2JRM8Td/tPTEcqrngwslUL8XNMB5yZTGxpYDIk5cxDpLd15
WGaeomeA0B6L+eKdD7SZLCJWrAvy9xKX2z016qjzli84uU3JcW2BOfGnYVfPsxesabFXq8XRYuul
aaqSsO4pHDVF+RzskJ87RQdugnfY8XvJnruXxBE6uqTE/dTQVrofRt9HVodBTynfAd1NraOz6XfG
qs7eXpPnrfctWUSzGgZSfT+HSV2ekPjFTJdzWNQ6tOr1ckQeXeF438ZFlL8lb+haldaQlih8YxAT
cKCoxVhuFvBsUIP8TMcsLBPVbljqDiud1L+zVIlZ+ea7+mg+sew3FCu5RTDsYDSiv0RmaHgQ0rhi
eRHemR1WbgCNLrEXVJ3kdGrdiyiyTLRiylg/Hh5Z2mxg2q3OZLkFg9HpLrkoQiwDQkeQLLOPaJ2m
Q9hV3lwXFtcnSP0eQGt5Om6JtGj8YjZU5KGeivx1oIfKddj1wvK6Kf0WuUMdNlDO2mKpOkZBH5EP
YPc2k1NbkpI2Pp9dgVXIHU+eyaBL41ngfCrpY5GC7YPga23B/zP/5Lr9A7B22Of/r2EvXl6DfopV
agv9vWP+zjdOAUaDGdVXSMQb1vDy2zhUn7RDRg/l6GCGwzbf7jwEPyjmQDEg0hQsZgL8/Dqjm5Qb
5So7GAWovmpjltxy/IxoP6y8zuax4sKroGmih4I4C014oPyaem8E5h9Wx0e7KAxkVzkf+pyeeNhH
OLju5WnbIZ8hmQwgW26oSo0hAEC99iezijm4NKK2R52kuwYWD+0TK5xE0fhNZ8gXDmRtz+UDoXXq
BaqB8po6i2EB1ocYRxmMVB/x9zokOmkz6bMw2D+RsghODojhdLIH+DWRy3ZMKtDzDdqF6bicN0T0
bxFaeUBAdxrGB3wBhtRGC1G5frmk3ACPC4VVHeVJhbZ2IuAzr6od5Gp5b4fKgQd4uhxOaBaO5djX
FRqvtU/Inqd8OV3RGxokRMrucwkZ8ctgclL8j39xU7b4jp8jiGNc8rJXcmDQ17jZQEszm1UGs87w
Mtlga5Ww/R+ekATQAX6kmJrjcDKTb5pwvaD2GoPtwCw6Wqvi0Kcfw8CqUhunsn3HyVmSm6Gp/6NC
BP+fpWjoXKpcE7S6sfTMlZ9r0gyoO4Ecbve3pf/i3Bi2zz5GwaCpbp+mdyan/3IFHvwXBwOVWU1G
K4P8dGpDoEYlbyYZdbP2adJkObqKz6yYqUIwcto7Lx+IHC6rMR0Zd18PRsA4OubCYlhPIaVZ7qUG
IeBZDV3tpWPzwudPkcaeP8SCNb2z53xxUlYnL0qrs8cuh8nmsdnLVOM9c1xOLWBfGIRPQcduiaj/
IgV0u9vl6bOKjji5zDHg+k4iPITKU6G4TUFGzWIdXB4EpDE9yKrTJDD1roXlSOnBNvAtxJ4i1Ed+
kRmr2SKLTtT3dVhssYVrRwQLYUWsKihHzZwJO5T5VFXMgODpK1V3TYNgJkMztq3vFAnItCnEFu5i
5AIbunVj/5PCFeps95107Pc25WqcJYLGT+OBbahJCYfFbEIT9LfunCnNdePmsmV8wiagh8h5oBqM
RSl6CV6YH/ebsbcKb9GAMJrIsR3TGon9aTyWGyKhx3KXjv2gAjmb9sa34CnWnhT6I4cUMVT460YC
eECZW1wzbMtSt6I+zjL0F8czd4atmRBSwSSnuVCxj5DhaU3BMQ1JSeoNNfJ0pq9EelyuxdWCizEI
oGEF8ybQYetVniKBtXvcJ+to3D+C/55I4FyQCohpbbpb8mpeqEy1kwuFKbrFify67Q9YnvTKIOoK
tKPk675So+ApGnDw1wL7oQAoUYKmElxktxFnNXVJoHSI2RTcKEo+bhUNQ0FGBagVB/LFjzjuNhRz
FzvTvBZr29NHkvMIA4IXfQ0hBTCnU7uHyJ8QxtzHBFtfkEZA+D2ulrawhJFxnW4ryT3NcWt4OUEv
G9pT9eaVry1kEKir0JKifz2NPDeDyzaAGEu3sgjTzYM2Zzv7w2kXN+KQ/M6l2ONuf/40ChlV1GFR
kkvIkqDA4ucrE+NTVeA+k1FdvwSPBBy/M0oQ7iGnHy35QGqXl6dcdurMy1tTlY3NBz633Vn71QyY
VVrbj5JC1qHl7xFnajbP+ICsmt03n42BVjN6gHEVKRgeWd5iusN2ulA9GUEMMbQfa1zXnrioPIzw
h49JTrP6HfAvzsl+15XjYKXQS/6cyTDn42vzw2LQRfKPMHDP/9pAW3EK1rt05dgS0AkBIUqV5bOh
OfdN4HlnJBLr3E3N+257nEJ0hJCgzKRQIM6M2R7ZqMsS1uxt5UXo1U5QUwA6IAm6Dt1MXVfe7zdV
NQYtI0aqopMmqRJhD6B7EbCicF1XK0pFVAzbZyWPaDOAbajDvAXkzn6vZmsJ7wrn+MhydOcq2Zkz
ZKZ40dpThzDiQVjQfORqjAA4gKK6FoAAufdx4OXdOomAyisQqr31ceGQhDyRVbR4G49BvCDQSRnN
AZ4J21ARYmne3EziN3LFEN5C63T0jHAv3vxdwtZ6u+xHKXrOikqhWBZoni/IMcLAV02qtkqg6afw
gJWYejlM7Qr5+pkBCO2ksYiRHm9QSY072hl82U/wcfuP3AMiAHx5WCzqgetQQdsdpar/qRdK5hbq
+FKyEUxBiAYwUH7OZzyX7yAPAmJQGewzrMnXdm/e4ZrW0Dhf1eicNTHn2m7VL3HxGRQN5r0GKeSV
c13+p2JfPrS1NLClbhLVKYY2GgmQzQ9ECr3IquRYCDSD5KcuBpGV3CdDB2iOLNQJMHIhPZv+7uNO
CxdOm9mzPzcHCsXM8MNW2Q+1yazy3WZFYHD4LTJidOQUTMxdOiSepsWYaxvBmMo3o+J96S52uKd/
+qgXjg5Uth+uBGBG3Kx1Rme62CENnjjiOfa4VnfL2GM8kWUr6ptwUWUYF8qMaaFnoZGmGvHE/H6L
P5fjoUrdB/eGSSTMsvuXeLKK8i6hYnXmcgfi+2SeFHuaDQOyMEm5A6GgGBJzScn2l3DloQBENoDk
LG/KDGipdfmwExf/wHetLfQARbgkYkgCi/GBsGozzQB9DDQIBZjlvIFWWw3u+8MgPV10L7t2ijbV
Bjj7cIad6svP/2aCGoEB+cle1ptI6/GdwUYLAkZ7UzAzjwGrQYvrjQxxTHCyprigJQN2uPwsNrMe
iHlGViudpUeGSsU0SQU8lUq6zPJ13h67kgcYsGZs+zQz10ocuaYTpJ2z+X2uLZm+LKLwSRYWkt/j
275lpxs6rutkV/y9gCR7J44hXEq2sWhHz4rFb6qI/sDLtJEx1Mmy35nGLgJ4Hcjci4emde/FYnew
M6vm5w4Cb62r6uQNHMJbUP1Bns9A3Fi2aV2ps2p6FcdCGkJPKZa6lQNZB1KASg93AwiZAQcFUtho
+yHGTQH1VurzdV+qko/2CWC0eL4NQHJ8+fH65IY+7f0qMHXq32t9Kdpp3+Jrth9Nfl+0KTIoIKgf
/63nEFq+tHteqe+T9H1qabnz5LtGW9Czl2WtrRbCPaYNUrBu4rVpSxZgxMKdct8o10477BsXdv6L
qApO8SL9X10Uu1pXrpgmdRpRblqSl6QGGgi3hsNQ1qOvrMvAixQ28zyP2a975/0cGWubye28Bfip
dpUHGvfYNqH0EY8wEMHKa9yZWzzOA+MD6e2/azPF6IVM+ZDUoVLoHVR9AWn7yn2eprQ1rvyZH6sS
jeBAPaj0Y7kAdky3qmfUglSRsk+K9tniMpQKuaMJiQisbYyd4DDpSHsZmlVI7/xkR20y19qWlvmj
MD7LzAixYp9EIHlQAfvjEWebVLhbn2on5dxZn/I/vpqktir3tlqcnwBYBBKdG+Eds9Scurp4+DZy
rOtGaIFNNh1SUlC+Edgh8QEWnsMLTKjvTqSUl7Teby6fzi/yFJ/o31qD7z66wiIxFh4TjHbvaaZ/
TGqaRTNoHZRx7KOzlt3sP2JoaDxl83wBtGJcYycpF6FLQUuVSiulCRb0hrnj1vdJ9H6JrDPa+MRI
CiEByf4J9xYLRq/SZCThEGjOK5cL4+qh8ssNwt8artFnGONn2aorxYKyfg+1I8Wc2IYbbkcq9CQB
+OoK9jsTsGWE+OPYyCRPPV8WkNtEp892a0QDULoOhqYIEoqrsE43k3Y/Yzqp9esHwDlH0pd4Qj9G
ywdtMvSVL/QtGSuZGxqFRfjPyzm9Loh6spvvP78IA7/1qZKBlq76AlSvLsOW+XgLpZ3Tpa0syM1R
YIKRYliEO/0XC4juM7mK68vzEXjdbYV/m1DAla/R2zJMqm6o8r6Vrf5CiMtPwiaBhboOCp5SS1R/
dZsabC1CAgrqFP8rOKxZJ+9omyAH+6DwH3Q2BnfodZdDJVonBNoZtZVnDqpmI02t9IFGIjSpcQab
l/PvZ2FtVAeRxVXr8KecMo57fs/3aiYmxTVbnJnO9BlxYSC7NEiWdktNqTAJGKTjVf0zaPXehC+A
74zQdZFgnRr0uvKQ1y0wzxoOuu6diPw057pnGu6HQjrBjDPq41oahRnQ0VbdTHf6BDij/HoXC4mh
8IoA1IWUnuss68U+VURAQSRUo2BKK94mj1g/rOrPf8h9glFma3n8qjbkzjXPHbTBTw682q2iTZMx
sCBpYWlxLo8LT0dIv+1mDzVXvJPMtii61P4httKuGIKuFCVGc4fmy7lMdfQ1el+haESgHxqzX0Jp
LnFIKR4vsFXSgn+T3GnVH99736Y1QztjGQNG2FclvlPNOsyJc7cS+oMS3w+0eJtbxeQzVSCfyFhi
U6uNqy9Sudo2ApYxKIrVd9Bytx+H/ZB3xbXphgGkP+zZ0NifKmSpNRa2Hz2xU/GB6rMNMvb1/mOZ
YYX0bRC+gCYIBsgMnZQgHsAlL8HSuj+kWSUeRKXkqJIn9XXpSDHATVvzPi2Fi+p/NUL84bEvkIQR
EJkyRSstKEK23e76XX8asY4ytUFNscQwSijaJ+3xPYJxF9j6OE4lOud6mzgwV5CIWb3QSYXatiae
LCeZrf+8uXehc21dtR6GRYMlK5q93+4Lug2oF94HUk1+g6xgpjfc7AyHH9Ngx+86pf1TghEYtO25
YEFzE1YZoXi+dNHgnoA6yWUsv5RrVAouAJePX7gmo+087bO6+RlN/syjIZSYWKrnOgIjTTPKXDig
yQI+xULz9FVxy++T183OHcb9Hlzg42q18Q62tfyrPdkhkM5km109ivWNKsc6E79Bx79Vt/0aklq4
Q8eU6HfuIxvfXHxyakbZcM6JoTh8jNyDuixfsMT0U2rfQza4ZwpfNS84oprvSs/9QfIkH1/rogFo
96AuTaj4ItGiAxpPQTKT3XSycmMZlctG1lreplg/PUSVlmpKd5eK5clYT5ILMp4IU2dn+rZZoMq4
cmlZopOlyBVFMHzKr6fTVgt6J7Fi4zPybMalLxFLpos1JL1LnU5+bDYAvKIVW+AE0glmr3CkZD7k
StRt74c5qUyHJ0tZIpac3JfG8Y8zGu+a+vSQ1CB8Z7644t39b+9X452wNhr9E0Le5uVbgBsQF7ly
l7nP8Rs5/ABUAgSBvCCqDicSCalreoJscI11mJTh5toO5SQD8OA3azbHk/RE5OBgv4QKbW/VyvQU
28bWclC2b9hjkwKF5zK/WHNrRQ0YfKJA6pbN9it5PPz0qwYhN/s49RJpFin07+SBPCi8uUyyBYjb
Nxt3Ffgd3RgJYiuHUlLsRvd8tjTypuesUDYB4jPO11oh8JT9z8Nbla+9ro6Yjuo/2KhU33SSUo7t
4C93OQvM3so/JykRLtmgHVEUS+T9tsJkJeuyYyA5A69z8ap8PDpg4oopGUuh30XGo32dZn/Zrt3f
cEtC6SMMDmkx2EwaA6mVX6BAbZuDhltGx7rfkO+UAMvyX2OeQDcZTxFHNGgs8RiyLpsqg75f5Rk3
cRHye10M1bSFLipjOAOtyim3tRXq8nFpEPx8tG89Iu8vrWMrYeH6I47K+weS+lvgt+I5tJuMKitW
fQA7X2tIVJt6gHaSDXpbUUqz/UyypWo11eJcpmYvm0iLyXjSN41TWOdWhQ7tWvbv6pmiVIctPFG2
gE8R3NdZpEvks7YjRDSXbzaDKf+f+0QMR0397xHFGP95/VJX3iSjVu07xcpDlJxoJp4z9dwbny10
J3SBGgJMMQ81+OCr6GAnnUsZEWnSagwud6DFoIVAHWXzIR6ghx3vQdXi/KNCf5Qf7/VuOaU4XIl3
uXG+msMiqkXt/uxV49eEFIga93RQK7CJ1zJbK56sQwYcje/gVoNOXYAE4MXqucH/nCY1oaJmQYTg
ugRAtdT6Waqwz+3pRZzPxo+sCPr1n6hnILFR9s9p6spj5T6iLsOVYu0YzpCkvRKm6aWVFax4LlJh
4lcggCE9aQYUi3TMllgJomLn6kNW7BLuDfmd0WlieAN7x6RsVqu6w59kZeCEM83FW7tpSrsxTwW4
8hTf4+D86gLJt/ug7hhSpN+SV9OZ3k2gBre9VxI8vmvgMTvaWfrWP2wBiR81aZ3Ic6lfazX+Xz4c
RufGdwnZKj8ynhdpV12nFEDL/4ELMtMh3IfwaRjSSaC3nAOmPh28SlCVGw/Va0igx+0Mv3/qOLiF
9A/YJ2FHWLgPbaD97aaFfru8mw41gMGQxvUHSXfTM6gLIvnpViLdsAcEQb3r2ZN7DHoFwTC8qwPv
bPTb+NALutXz0PmWOuzoDJBRkFlDOlIc8auqL/4KLJN2DQUqDVZq2Mv+sHGZpjVAlTMGek8ZJLdV
VPfmoXrF8J0fz5fOsOcHsTQs+3wPFfzXyJz1mtNLqG2T43EQDI6dEkkREjBkTYypR2nF/viDU46V
b47ja0N64D4Z/iwt5vdILsEMqvmJKZwGu550dT38QTSB/X+1aMdILP6PJAw2PNSuVr48bup45r9p
x2s/AkO4THhkCotQPF7KXVsIGwnl2j/z0bHIryLJ9Tx/GJh0iAAuvi7MpbHbNLpIfllQLR3IR4ms
ogJmV79iJ2K4PhfgdwyUG/mKzbBr6/U7ERdueBaq5pwTeUyAlriMVAUEwodJ+Nvz9LVXH3rHLqzl
1sJVNLvW71VAS1x9r3CMf7Xf8nWsdZ39QJvaZpeuKfD1ytBV904HjXNPS8Ofe39xiTK7vWbTtsHC
NK735tgMoGZl5JXyPR4fj3NMDM1GL4hveg8d0cWEQlpzaV7MqrRpQYL3uDKmbAwAV2Hf7SwvFfY6
w/aip+hb5X6H078qvQnktoyW1WVgFqJiRJGGGLCqtYuo9tzF4WlvTK96Wg3zoke8/z8NLYYtNf4J
HwQhgJXEK6mdMHFAbxREYNc1vK4A7gnlVAhwNOUg+XgyzN7p58o2ILpOSJQ5CQ0Tuex2QWEi3hfc
icyTKX9xLoGD07DpSEoat8IT7VFqM96Gz8kFRDu9aDGNNU7xKYjksRjDDD45qOvDKDUK6XnbacIn
wuAzEaZGLp7v/CzDr+pcu81t/ysNypszVV8OqT7/iu7ibgStlciyeO7XQUzlOsTPAd2oIRxtwxGY
g9iB6tPjs1dnjNKjJeQBYVIZ7OThNh+tBrNHzToZVhmhpWzBaw7q9UJUqd1axyFXMFFo105y9kRe
G0T1r6+YiWUdPY5OPpTWzHUSv1spz6xt1B0ZKyWa6E80ymEKUkhaYG+3SC1k3kAi8VzeCZ0t9fFu
wxoLiYz5/DHN+nNfVja15kAFFyuz7P4XIuRF3zCBSrzdn0nTayT/i1RTeDycLDPdZq8DTTTi+Mhh
dAecfKPksktIfCu7c6bBjMNfiJGzG9ybWUrpsTU5qtSKuLpR7EknT37CxyBYafpv6ZtwQbUWI5ar
+n2c3gAdqApn1tBLPT/ZoXcJCqUAHyketg12lbLNUx7I9TizthcAJ3bIvDPo10zf2l9e0Tdku9T9
sQ3E/FOyC0Nie/8kN7v/YqIlqiBtbJO9ZgfTq5aC+Xx/OD3IEzM7mYeEzMRkGloPm+6OhJYlIi5y
OK2398SEYmX2Ufm+8IxyHCd2ct5Bp7DsB3erteCEHcBQWUYP1EB+dg9fwnHcsPYRC6C7C6sMzdEE
eJiZmXNyDXddIUXu+EbHdAIwDnpsZe3QM6T/QUGlX/MyJz7v0wl1eIRms2mATr4Ob4khHa8yK6S5
zPJESd4UWaBYzApykfIgg5vnz+HXw1+BsB7jx9wiWcvnYDPFCGBv9fQ/oE6B1eX4yvJvjkjvfFWf
jCBdatHsIHMhzVfD8aqD2QSTR42j4FYADCNBQLMEBTDnEDFChP0yBthwR8TboMeuqvpgBJOzy7qj
IV1rsO5Wr7YBntkiJ0Fz0wGDoi38hCxozkqiDEMw5wlYJ5Ax/NlA4VPVZ18C6i+zmlAMsC+4/0gE
73p7uPSpTaotcL9phZ8vRs1sbQR30utzN3DMLO8l4B2Ux8JFPFl1KSjNYgASLPucIkCeZBb73Z1z
ddzp/9ZZk0Amu3QmhaGQqseIv9+M05rrNcZDTmAfO3AIV9KSx+a26FZoyAjpCiIEhtr9QZmmOmT6
Cfg6Th32lbXlm2NBGBZG/fWT3h5VdpHiDZt8GlXNCR+MyXZEy782HmxyyhH2R875+G1FCSj1Ydjg
hpVNuxf7HPeq1TKJoNFWNg2N1NNdzV1ejwzuJq/slea6glX7FMANIJ9ol58jUaWWVGEbe0dzrpHQ
khhwoUbiMxdfZoc91ZEshAIdW+aTqoXqsydy3ahMTdTr57P8zVWRr2fpYfYSOucrOSgaHXN662sh
dIa9v9gSpp3uIHZkRBzgqIW/Hww2dntfBV2+zUpv5iS5OvnQxycvFF/oMDAVyb63FlDDXwH1IbPu
SED2vuzXOyTYFHMWOdqFv70Nt0glA/jvWPXgvcqVxAV7G5JaBJ5yQ45tAazbekTkjAS9E1OSTFP6
bsk910Z3jrJnIUHibBKEgfOR29fRxOqJKBAgqY/2ChPmmrCf9aTg/cesFaiGUxc7mDfLBln/xyip
0/8ZuoYfDStyrH2hJekbnmjlR7xBQthGqtAs3DD35TEUyzX5NA2SmVSuQVWa0JQxEHzBjOKWdHF9
vkRrDct1wW24h7pzmr8VpLaz0YmYbFYhbTJiHS/+u4ajfZoVD9aBOq0faHGL4KCibHoSIAAciY3P
U6ZmvKOtkiDOygXnFdvcCCndaqmLC+7jdFKu+b9KFdvad2BF5qcfk34tEHVCUXf/7DX8ek5DuEyt
Mt+6pRsBTKMNt8NsBXcV1Flom90GU+ZZ8XR0t54xG0K/o/fnuvHd+DtuCT9UeW8SYHHqdLxzkFUE
kUdYzeOnsyRum2huaffOESpi27uHl8EJBzL0wGB/zwhgqqqOCXn5TG2PLYcyojDdCLXs+0wlj6lO
MGwgPJUcj0l3NnYrB6qqXPpH6YE2xhGht56/Fqlhli2OQfGWAihCge73qdqQiLNf09puyeuhgmqw
8zF6y3bT8Wycon0NMENb3bKYGrv/Tx/V5Hecc6LXxeABAo02b7KrtUPgrYQPHAXGma55pRPTUY5P
9E+6y6NIu9zJgjdoAhsMTorpyBEiGLohJ+UmwFmiZdKVa7DVQlyYr+hTG8CWUe+qpcOaEJE/sDgz
CCrrLFXV4+sWIm1pPwWSPJrOEcO+KtmUm5HnWs1kPKEfgdLjyD0xbBEwgIzbV/pmRB7heOnw50t5
Cjgteisexu4mHjQjgxtHhMvhKvH36HFPD5zAq5NHNcRwG9k9levdyxzZb3cdwB+Gar39yFK16eBn
gxfJMWRcbStsbz9izNhRHFjlu4N+1MIpByDYnDbj0jBSRbtyJhXKaewAQCNCMCIReFVRZGXTBm+W
0ImDpG/6xXrJ/kp8uhO3erPlNGkYVzg3rR099H97ziaxIXKBqLA/4OyfPX/DWm8jEGOhmmSV78hS
yKiygMf3tx8cNRbMcJmhWyZKoXSMLU4wUXDGwR3j6PzpSnXw9V5eCTRJnl9RLHQFiU9u1NZTa3XJ
XkhD/yOutTm4Kol0Do9MjmIwgwvyJWd2iib5c7BBE67AftFdH8bIPG2h4amWFA/n7tB3E0jEHcPe
5SNRbjFwb2Np+K2XhQJ+rF+8swvYpAI21v2UyW6s65h308A9ybH9DkJ4j+PfRIif8YX2cI7pbaCL
suNSbVP0OcoNUCMEKL7Mk5hc8uW8lv5hVA6OdAkxpZZxNtFHYVLTB+c/vmDpYNtzm/igMgk4yNbo
OsVWp9VQBGe+RBNOHatA7+Cs6PzPYmcKvPyLD3v8D5W2cfRDk0dt14AI8zqHBcgNxnJc3UoRqmYr
6Hqa+Sd6UDxt6297L3rfBAeV2gUvBNKaspuBnpNnIneYuiuW0W7WxmW6Of2i5LEVDmKKXFNL+9Fy
Qf2i3zPVUeYKHp/Zu/DPAQ+64noB+jc31Uavwpwok2iDJuKXczIIFUgWFEIjO/F6V4wsMjLk2h1f
Dvcx9G1LKyEQ4YEXzN1Ry7vv7gdh8TGAEPilH7doNpG8mT4I7pufS8uotZVSinpVySPDb3YXwDX7
NjRnj6MHu9j2xXqFwLJkhXIwGM41FxIWdq8hKHCgV8GSSuwUQut9WAHVVrdWb8FRDhtR1dGje1xQ
FWV8o2T/OhMxTO9wOBexhXbN2eK8hpfULlZxpjxLTWHFOooOb8d7grPKrp74DRI9y9pCoaAt7wjR
HQUZofkvk7Y6YpFZK3Rk2xbf7oixUBPJPVm2nMyky7yn5fTun+5ahDu7o+aMxhZTXZzAgU58nT/s
6c6Nqc/Y3YQ2jOQFdnMudYNiolWAVuCfHRqF3R/RtfRo80HwMbxoFLpvvO82BhllhV4vL6bJ8+EY
gDQZrR+OEcIEugXOoCwHnkYl3Gz4u6E0keHY9couHluXRBF0Ymrxv4DeOa4D1L4/YFmKwGjbeOcY
JRqWVGqQhCSygCyd6ToEKZ1SyOGLCWAZd4hGJEhHeIrTmMyL2dYX75DJgg8gaJ4BY6iRwvvpeo0v
IuHjPFn2gLWAdr1ZVx937lp4F9autsQjizvGyC2tbvhiJkJu9XellekUoWgv0LoNR43qxmVIjWRS
zOFw2aGSvq+2uVyu69GjQk9EVvvi8hOCAt0e6VlkI8986MLSMq+4+/FQ9lonylCaONvs0exw33Ud
Stcd1gPT98yWFQEJrHM0BA496PDvlyAZX1jrDUTZD7QKErQGc4odq9ZnIlQl9WvJnObpCalsWY3b
w0p1wknZoluS+h/GDlufInLvSHRqnzidaTv+b0ss7c9YDsRje2jdJ1AmE9ugk341rzZU5u45wIo0
4syhSnEyx0th6AmJljoPw3vNpbs9XsvEAmmCbupBNbG/quUcbV2bWlcadj44F7duj0aLLrmXZrMD
pnp6UswcW5w4s6FlpL8UU4CDnK/6tFM0uCnBuJG8T8QxABIjP9PnSY7ii4kSU5tZsn9ucm6GF8Ur
Ydp6AQhV1hGqvEfxUwWXeV8bPv8e94Yzmx6Nj0B82/rOO8aq7CeRY9wnSnRhMroIYGD9T0N7vFLe
r+TchsJ+ftH2TFh5uL5s+ivuUT5TzNJGTZ4wZdStnIziCfNzB+RdUzI09wzBvNE9vfS6hV5eSJGE
BQVwBUEEsqkzHrmT8RzkVZsfziwPgrsYwbrT8eo2xjyCTtNWzYnZqysfWwN1d78mFK17xRXzbslP
HyB416scD88jRAlgDTHEIghViLGnNHt2mz89bJGMjjru4NPaYCeKeel9pjLZ0Ac0b04ItkIoxNb5
DoVYdIfofBClgYr1s2nJEm5YCKAx9Vqu0XtESd2X1NkzWeSlTyob4TUdVhR009yoRQL2JD/aJVhy
DM9kRxN4ap3his25DAkDYSdNl1rcbodykUpjH4cIx5R+JGF00y3wIF1c08Fp3j/ghaWgP4ta949u
GZPdkpuoYJIx7KRYQP+SzLZX4g1rb2sNmS5426mdz4BFVLu95lUu/m5/GNQTPaEISBfdm3yizEqk
0v/9iIWiedcmKh8rxzt2a9PwMaKPShvNo5eb7eW5m/rxDxOYamz8lx1BnVOa0dF1fxt6i4zxiRf5
ApxGaZvkPIQaorLfBq8V3xf+odrdtpIs8rsQVI7TvizKrnDB1EydRjyq19a3W5ueS9XJtwUJnncX
PndEg5f7xEWtCL5HlX1spyS2IkSvFnRrMOHTYQF97yEaOCs4QIFop6NMFbvPt5SBPFz/kAoqjaVi
dU55mEs3ewtDpAsQu9OqfIISbr7GdCHpJfWaS2lq34+NeACTcq0xWQmoJpaVkbhEwp0Bv7cttzJ+
eR9GvDwkCVJeIyLyG0F1+tshuru4a3cThlkTe8pDhCDUwo8h1lIk/BVAAkzPJKnwdZSzFY8tFLwf
QuExdTT+hOSmxLe2UweFCNDP/T8Bvmjo85agdx1AV/IeVxisVTQm3TC8OmIJs1b3W3Qcaoj9Hqle
82M5N1UJsVpSV51UyYyicX0xTS360AkA4cl3iD1mNH+RZBi+qomYow883vwUiFgM0jbY9suwzxR4
FWzABKBb5G/RVmMlCwXRTHpx+M2+9ZHoGBNjFM+MkDNXlbqHq6/KruoVVnve0oi6lLwRRdQRBTpl
s5Oyn3bnZLINAqBmuEaQIiTg0xf+JZlAAcyLEDAi1zUTel7JxYvmbxQ9uYsfWVBgn00MTIXFJKTd
drsSuipp/gFigWjxRdsN6Pet2MWX5H1hidqGCmh2fib8nfleKJ3B6FS4mvZbUUNThER+qAGXYYIR
fTFVZKVpl4xsbNWUqq3Fem4B/EaCXTYnl8O9VlENtbbkN+xa7qlohTvh88R46x/M+2GV0b3/QYRW
ArNdfMuOE5sav895WSSJx6Tp4biFVs93eMe5O1sts+M5TP46aPL/6QlWauDvF38Sh6+pGq2hS5ci
GqWIdlVVHxtFhL8yeWlyf3onZpPkF1BSzaVgeKcS49riO6FNVebzEzp79f/pxBposo5dmqQ7XvkW
cABrTLX3wikwi01saQQBI7XIWnZXLfSAyS4qYEXpTnnnGX0ug3S84zJ9RMG+YOXnxTzrrq/Na8nA
5Qcwip/3HIGFoHv1TmAMxNaupf+2Rjn2OYTGEw7wTspnFymLM8vT76T2JsJuAwB5BdfdPbeP6iz5
gWwxGVbnikvzsvuz6GVIHOU6OgkxEqaHMJAS+GLJsHw7KV7uF7QaL5alqXMtq0OkRWOjJJGPPzcv
84LOO96oqAxmpO+M3adx/VW+2ISLNXLT0tRRACq/WL+UNKlBLFtNAqu3a4xAX2rEAQ4Bpi8yrxfN
99jV6Dkgji8vgsRJwlDGf1YWd5JfX3wCOvwBBf1+qs9b21ltdjbIqmdn8Fk0EIge/mN5piTYQ3yh
Ur5krRqVxRfnuhhO4oGmD1dTUVaIib4N2VWqvcsSN9fbXuisdjKJxqkIfXRMj7tLukVDk0VAAuxM
ZysUVWyefbBYlfrtid9Hk3RSEqtWBIrlf/PJ/bpHG+ghqxSmsmQlXFQC/v1p4unQVbNG6PoEgVyt
/hEfDx1XL57V+RC9YqFfrJdrQu5We6STKOpX55IVjwGdSTyvG9WkCkDe6/p2ATfRwAeK0r+k0IpQ
+goBl7YxNzLNCx6/mmWbikzTAXyxS/FTDhQkmqPa+RfEfwEEVPv3PXke8N3ZECtzd/d1a8DDNDSa
xP9weHgQq8dXjPUlitYFt2FVsa4SAUC2B1OdmAP9qnroiYVP0TnFKg9G0TjWGiG39gDZzGpBLTOO
hcr/YQ4ESxv8mK74vpa8sMd5idLgsbrTGYWqQCB3rofU4VSXUdqqHBhxaQvZuQMbwpCgOxyVU0Sj
nCiwBStR/o2+sHeKw0XxpewPjVWYU6fhpH9IG4GAA/NFRox7yVYbQYXeRul/jUGCkBYlUoloDFd3
88LgvqFv/uKacviqd4V3zt7Bp9ZoU2fOcWiAt2KiwyqmWje4EkmuGCIeQJMz3FHYGvC4lUP/BPQL
bmjSlOZXPnFAwMqIIl1OsaqwENQ9MunPJrIHRBNLCHnQOllAbGT3sy2bUwHAv9Pg8fCA4Bg/4L/H
6wYhjtDxgBwfKZqMoXubj2rJ/XBVYn3Wpb37fIxZwgkXsrQMQpc1d8bmP09Rz1ZT8A2BE2IxfOPd
K6aOib6HM7I9EKZYt84vCqgWBdw+BAPBwbiRxxuvSFFl1voPocI7CKMS2WdyE4gq0KQLMI1qn3eO
xwTVP9uBCZvHzYkhn0HMtH8NypXQphgxslsbHvntMDzzDPxNtiHIBBm6PeV83cRAbuQvClCQXAYj
u4DeXG1uZMwW9P6UPmg/kxHgxRnrkGp3s2jpaL6yK7Z2Kr9wav3ysQ7MH9bEA2ydDfNuBQvCaqaf
4xDiGfIWtSimvKlke/x8kdjQGis61u25hTM8JfRfN16Kn6xtSXJvYbRF2nFxHgA24mFrAIUjrqTi
lRtn29ogxSdV5IWaGkmybBIx+yvF8V9stEoOJd06nJmnWRI9kaokCRcbynIomUcUKl+vSbHUV6st
3kS9DSjfq+T0RIs1Cq4gKtutGwG+bane1WYSN8VTw9l3cuRhPbvI9vSoj5YcmpR2hZDYPG4IxVEM
aiHyOdnkcAHogP48sgOdvt1J1wQ43czFbMe8dEfqZgaQuaJAHhRRRHyZ5ijPXrzmfoPpMLauBtWP
8ndPx9CPU5w9vvIrnWffuNC36GeppJi5tAfKyPbcXRuoUJIUaq4JtmM8w9BUEyCTFJQaRdq1r5/Z
iZSyQnJqI65kSYC9+U/7i2rNp8ZiMPzqHWX1b2xiY5cIPOL6ro7Z1/Vd8evux7Il37tS+CzX7346
KZWmMSTRuJWGaAyp2ois61wmTlIUF1pyIst9TkSBG06sU7zV2Y/RqCprU+skqtE0h2/ajh7TCNHA
b48kCzezdDEjIiU7irwDLuN0ALo2gYSvfcGdNn1lyvsp90eXnna1f12a4NLocPU0d/NBnP07u5Cl
qWLaCFQylqsAOX0KUozCjP3EB3+Bv3j66+7v4LaJOvB4Zc5FB74q8+3KsUeMyJLRW0I0uvmGv/Vn
22nET1qtz2QCV6AXy5TpjAbL4yMzqfkNcm4rB2DRIZQ1rFcy5JZEeXQAav/mJVOdy5g1RXDWo+ek
Dfo4VNMiFTtAUEntit/BDdbngx6yywE4tEa1i0ZpNZbex9tFPUUJTutNMQJauB1Y2kQYHn2prHtf
4yMpCIwJMGW1ukc6px5GvA5VTHDXsIYMyp3YGlDZqgwDt9v3vBbGmC9yzV/gwrUdKBQWB+22AAk3
hMfKRE2XRKj90WYclwrQ86qx9ZY5Q2Fo0H8iq+Q7x1m2b+D6haBLLJ1rfWbNQC/ia0xuvayf4c2m
P5MpAnji4lUgLq3VXcz1k5RTPortnbCsSk9nZRL3pCdMHAwwZn0mx9SlR5z6orEYwv891qTo07YG
1HRcOXnpmTc9ensYuCtZ4obTXgu5nQlXBd1Je/HEluLDCKX5cuHjT7KVz7oFpDcWqJbHbIRG7xH0
iZ6RajNgJItcCPbINQ87Yz7yWOoozW4QLXepzkEQC1/Bd+HLH5i8wN8uKo1aRRMl1YFeQBzqJyiy
J0Af8pn0YkyXy+757rBhssKFBRboQ1nIW1CGhaueDnhIqPnLxqUyRKc/WnqqZM89swmNrhU+m1zq
41ME81Vo+GYJZGOKKDZiJew+l8x7N9v8avCg8KEA/CCVTsooDGBN4iI42jn4f89U93tXEXeELJqQ
/FHoiltmERfRYpsKNTB4jsE1+Nx28PmrcuxJyMdK5kgFW0FMiNAKiYpyjc/Z1uOFyR22zEa5dEo1
C17M6tmadq4f1gtDMG/N/kuwk1zor04B7/9TBrbQhHWTjtlltdfeiLN2dJc67ZXRITf45chyYVL3
LBmiGoztKxcqeitwAg2HbJccKDYwpQxG+ihk+vDTV8+7jUBHOjeiu4Dvd0Ew8k+HklKCE7x1MK8Y
Q9GkTW4E8u+eEHNv5iLmN6GVt2PA69JEi0/knioXHwjDMF+MtWSc1pI48Xz63ayYAm2NYVH9hqjP
DYIyK4bt/CsQoqThpKttalFxkVKc3ZfPBXYLnz+h5oRpULD+YS6qDheXI1Y/pGmLWjzFHKygZf0U
tc3ZtBz6ZfSg3Z/km5KlNqcZ6FgjH8LsI90pP/zJ1CUF828lUbsj3mpceGMj517QBDAmsS0IZX6t
vjqn9w6lH+r5rOOxeBkRsNwM6yGhvJA1XZrKGcci7Ra44qs8su5HDASFTrite4yHfejPNiK0gMC0
5q/lJIpQRBvy9othjxZ0MZew8hv3AqCYSXsO+QNaDVNkFWYQuKz/KKYu8RaUsiMwAVBNlnUv7bct
7vVssJZO9y+g6wJ+NAXY8wypuldFRlU8DRW+2Q3oK3llUjFhngEWoL8B0kLOaiU7EJkmYNbccccc
7ixpSuiBxJAxvrqmxMrlxIe4LuecBYg3RQ+CFkjXWdV+kqBHOJ6DtuKuQPnpeHs2j7Gj9xZbehej
/p4dltxYS3hmrh+uuagKjCv028PoME8Cdxr1Un946tA7JK12NIU5TV9/wj1qJO5ojuS2NAIe+xhU
i09WjcE+YsIJqsKVJUTPsMs67s+DYxY3CjoVbqxauiAWf6eRsEhvuLHxW5SvSPeN+EZrPg3Baqz1
Q3bdYHD+DIrO3IY/nOuZLcVOke69OqtVZiaZbxdH+HTFob2iPaj85DevC1g+MTl39h+9WJVs3+SS
9GtJ8TZYPYr2Dhbtf7HuD5QObVrLpa5FrqeTmAQ1VBcNrjX7v87XMJZaAPWplgMgUHqBlM6U23oi
j4mpdSMe7PTnAruxFzn0aP//q1i9Kjc1LVcOuOJY1KpASZ3wE7qm7/FO9sM8MuDFcmqTNQoc7XrD
O+lOpD/cK6lyo1Wbf1xBJ1aVldtv93AB6uZr0hXLveHfFzKNU0eRgUSy+bMagOhfcmeYJZs4Llta
XnFlDuB5wjz4IMRklZosVhoimuhZgUBKs1W15x4rYOzWvJDj47kgIgTUlXCBV6deVOQC8zQDuqUV
sd3Ucr36370IuOoZwQEQnakuQHfJFoCZIegVuldWLIDGqsNVpB89MJPQMqto4h9S0C1gN1fCmrMg
0EMY1DvpUFAZw2kAr4UegsMt/K42ajoJuV7K6J/ub23NttutIw88jhzUaezaN8rr/9RcjO8WoyF3
AvEI2z2JIu+8TcD4VKU9VdPsFKbes8tzrf+AviinQcgEa8XFabAnZtquTmelHGvcRMVnvUq91oNX
L9ZhwG6x8RqbnxZ5c48EXVFeHnzqFi/pXujayhSyt4ehqoNG+KZoyv5JB3XW/IUscfarBULl/lVI
zU46aKRPxZPKLW6RghBo0kOYv3kO+ePaK33ZM7uCLXGLThd/qIQHB4okpvkW+dYqV6cNQkLoEx8x
yhwLvSZFYfItDURwlCdWzngBGy/Zx7LBtUj0xAnBVA7oKKc9L3387tVf/03b/AgO1vifDeLvGzVM
cyNsdUZ7tAjhqtuFze45KkSpFf0nl/hO/eIk/qSmB4JY/mVaQtAwhlvMFVG8z6ux9lsq5tHK2jrJ
x2/qhV2yECTNKLbkCq3BoJAAjDmSzRUF6WgY5763iXJDkRiu0llIibhqarX30lrCXip/vRwW+31F
dPOPMuTuoERSxe8hbrU0yW47lk0QLEj+nZ8vMCzBTllkMjCUt6sER/oSKQf4EPtnwFclRWIlhC8u
BHxOe1tA0CO8QRoRhXmAlfnse7JARrHBGdM7nLCvT7CK8t7MRu9kATxvM3aghgKUt1paSyzlI9t7
XW2UM3QrQjU9PFQoR10WKSCUEGBGxDH82izrG/5b8wF8oLay4mRW4Hnq5Srpw6dw0ubeEiyBvl85
KFBUydmTuKJBAipQ0pA+lLlpsQISLnyvLWxWwiQ9iWNAwW0Y2BT5K+7dFahr1A6XN7qq0hYSHfxZ
EPkS4LUHwCDBbMEyXrthanuYUJoA85lLhx1l6GtAoU1qlo6IPcPXdpUcEapAHgNB5WhAuKPt3e/o
4u2cM/NcU7O0Mk7qIkidFHtp9AHKKy4QKSrntpfSMBpZEwZVZ6z2ud+eZTqnpezd0ulzt1W3C07C
89BbVUkIksrNB3qeoqs3oJSAO6i4d8SnkQcTdbZ2hNy6z8aUIlvo3vZX+OZv24Crlj0k2nKFIbWg
kTE5T4QsI9w3ftgnP40Ud7Pn0VVGSHl4mnsSIvx0DKB9ks/gL6qp9GmiZacUMEmzVvhGVJU6/Ao6
q/GmruTukfwW3xd8hiwaJiNfTkgfxxocm1YkDw0hzBR9RbSqimbs/kshCSlFeCxHKV24x6CYG3Xq
MByF+1TGKTVuvbFnPJF+pw2Rj0fx9CTKi42mybTKapWUI12XYPheKLhtkURw/OGXiB3qDDDIqc41
A2W2BFaI0MyzPjhJ20smkZQimJzx56dOmbA/5DhREQULmz0iyQdto31YBO2ZG6ZD874Ye6XlUPMg
JohEhdxloO771oY9IFDAcKGbu9gFzk8jD3V354Od5pZoa0BUaXPJNnjDQuxiERvIf+cR+oajEs+j
rgKlpLa9gTxPdOdr5iEfTqkDg83Nw4D/SjJrSEK9rr3EIBm+pzvk0c6CLud7ZCD7FWWzDf/Wh9Sn
yAjqY5Yk865HELk6scXLs9t4lEk2GlB58ogs+ZrXjt64HM3yG4EqfowYmAO0ms7RjuYpFQ/v9Gab
GEiLAmXuHBVzPpYr82MHrHJC2ZIM0Up7OeGF1xkWufEAul1+hBERZO7/UY/Pi6eFxSjBTnBqgrzq
wS1zmp3hvJWMx14+XvZv7KZVK4kbAY3JOzZtly7NLlYEYw9CR/03mE9ZP1A6gyLvISO/htoaThlf
x5ON3Mg9rVQ6gPOZEwe7sZsqvsjGB0mG/JWSvZcK2z15K0Yi5hXuH/ig3nPa+A3gc2O+8NBMG0a0
Mn55Bexf7GBecc8KxKw5ZjswR64LAUHFaC/BVXpWj9bPOht5MDqtDIR1/8Tj9BahNjk4OBurDEhC
6Yny0zyzXj3wE+MRdX8lJQ9O6t/kYyMYGRhJmEV6J8wWDFSSiI7CzxhhLfA1v8nzcIg6zTCefgGv
kcvHurCSmOKYc98OQdd7cS2w2itfCHU2UHBAf1kRArGJLit3IHGrbxcWfLAIUlaIpbBNI8CskLed
Zljv4tk3T4u+W2Hs6nCJPzkAJtBu505kF2FuMxhczjO/IBEq1ObmwT3ZwXiE+FayYnzihtom3GKv
6DgH/RwDBa/cbniC+EobssvzYTq3zqLZ2UWdvN4GQtRAUHhpl4n2bBn0bPyvDwQLtLFlaYuTmXcg
f+VtRC51gWk9ZR1gmpDCYOQJvoEjqJsg3nLn8R8jlahMnsK5X67YN9ndWeClC0sVtqAHkI/tlllC
CrmLoOMXMYqg9ibGaU837MkUR2Sfa23WSEHHcQ29eWumLYnRtwisy9Ukuniw0mXBpVu+arx2cKIu
X+eaHdKkPzWVUW2cHAO3VwxVor9x+KB9iqGzrKoys+ikOcNqEwVek/m5SnEAtGYsJmP+dD5dpxMI
DZpSlQMVz8kJYGQX0adYZZVfejNJlF40XMWXV/NqqT4EDSN6rZNUmaNF3/dJdLnyBFo633lv4qLO
vVbX5Rh//fgutvou/mgyDLPwAXHA8r/pP0f0DMmnVpKmL3tjnABY/tHP1qgo9nVb4qHqh+xiNtbP
GWBTr6D9X28y3jRvZ4da9KKsHOcwiuMmte7MQFnmGXW8HgxfhlMxAM3PKLDntFwp6E18W60hw72V
cbRzbyN9hzXwesQmhtDKlE2nEKeegOQUDpQyvTLpvzl9eHDhKY4IJ94z7XGiMcqiFCyXfYOs85qb
sZF/tInLlCXqmBHQDhcUjCUvCLUe8BhAopbIsFwSk2lx3fAKTbUUO/Q+JkB7PuAFUgGlAbuQMjf3
v5J7zG1Wk4rxpJL1Nk+McwPA6NZBnRHOCx1lzFl6To+gQrfxn7CV8Ja+e6JZqfNXmR6kZMmjblGa
92Iv3diKQjG/yALTn34aNpn24gjpQL4662qVM0RmHvZGGcF4ww+jGBcIyo+WgV1XhzSffgsKCNpM
LSADObd2Xeoyh3ot+P1k1VVq8Z3ieN23amTH/wzSmiNJE+c2ZpnX6iHO8My8KBtepamP77AFRoVZ
tkEOzbF937hdTyJu3OZN3jGN9CWQovFrEf5BcBJgtKOlDMbUOKGgTiD9BPSMtwVHPSPy8sVFlyof
rCJTlUVCCjL78owdfqfnM6ePB+zGx8yq+2TmtgaoIWzN4of4oGWn0/WcN+aWz62SrXQ8Mdu1ZQUL
Am6tOQBcK85bxlYBvHLKXma0z2jis2tineteA+9c9Z2trG6nWS9fnMUoHJ4YENCkvv0i8BSD+rWi
/zbAppxHuYL5YB5nryZGLkBpS3Knf7CeqAA4VJGLcr0Mmij7tFDHp6PBeRbADa+c/KDLWr1fbETm
/do+yTKfHswpnobWvOzjK1KI7fx/tdg0O5T4n47FZYlAxJwYPvh1MZVDjqv9LiCX9eCVubSc7EuS
kQIhm0Ypv2uoEebEb0Y/iwMTmlW67S+UfKQvhHWsUtnPWFfkKboP5NqJ4sDE3bztHTdOQtB1Ad2M
0jhLzO1P1WMzDW2EB2GV7JeDzd6Vn+n4EIiB4Ka9GOh4irLyVdub3PovrE4SyoJL2qKKuxA8slzK
C/0vQRPehIVkxGQ0yyKJH4tZKSEcV7a4eGWh+2hf1Ivif54Vle7quVPnpD4oaaZkU1XFwV9lEpY4
gLD6I/A4Olg0h2LxGZ++0FTXmAHIMyEOn3pfWT7R1sndWh8Lex+4Tj4f1rI7jXupD4bXbdpDvt3U
Qs9SGHT9Gp/+A91slPCFb4D0wHIrIEqQgRp1Sf2u82zNsMW6S4mrRVTLjT/cYo1oXbUfLIPpMamp
ZMqvXBCb5rsP0f14nwtk17fxi2dDoXXB5kD02JRini3tO4fVOB8yhun7C0d7USRpKq+RD9x/BdIf
pQonHBfLcLCf5xNipsKMHak6H90cKiAe2O4NLFvjW2mGXMiEZXRawpM/v1XwBls4d4dKNjcYaXRr
hEAIqp1qabQn870T13+wRtVnDZziAbDnue9Nr3wfkMIitF1oLRAlw3A5MPLLBHbf3n4uztZ3lGar
pHfcoB+OrO4cfl275kTN1QeZmcZOba/uvElcSlCjPd48TfaxA02ZuReLvNVcnjaobxJhMDs1euhP
k5m5+rygkKYcUvk91HpQ0blG20EYp7Z3GDeR3MaI0tujQO8D34QjVBGTvkq7tKX9LlCLpF8xpZOl
OOUO5QiY7EWZXaBGVLg+dnw1YdzPm66PVEhk91FHiFW2kJXQp59A3a4EWFjpAuownpMFQZdBpKlc
SQ40oPKKqydr/pe9Y3XIs3JMfiDBLzHtznCcq+2mjvLq/dX9sprvl486Oj1frAhuCUYe5Gl7Vg5E
GdV4ULsofYdadApzp+f/Hqku9YFhzaeP0E0+ifqS4Py7rfMkxVw+HKT9QjV2HTyWq0ndRlpqrKpT
vfnkWHPEQs0sxilZr8bbaHL5+W0FJrXjAWf6Glmsx0EZzh184soy18t0wgmVtsJwWej0OsS9KWey
JBB5ClNlcKnbyeYAgVze43Of/n68khCKg6cpRu4k23N8F+I3xr47YviZICFJq/PZ6k+cwqsLdM90
U8lx3H2m8jJdIskqcu/LbNZEsTCDA+rnbhLDa5JWR13zSUUjfNF/PNReFm/lMddC1l3FhumrNbO8
sOwn2MO4KDC6SPh0RX8S6ZGF77M/lCosYxP+62qJqgAmHmB1FWC2ZjgzDWtIiG/I+KL6OoUmAe95
KOn9Xg75t6SPtDG6oIfMZHIKlxm1t5eELo2Kyqd9Ha3/Fr8bNCCnYTzoBFOh13cfNCe8b0WDDwYD
3Ta7ks+S6zqmYMCLhf3LXg16jDyDC8+g7DQq1bUtIBSPzgov703TxeUJeVgCshBvNQrccoTr8V+j
gDA54UwfsjDjR0pr0uBq1DTaFzm2M0FMr702syvz2vLEYErHxSWIl3WMBNGX9kXS2H9JutFagvxD
ib6H1cmQ9sJSszONhfumCCKhl21uF/INwn2qzREnGDwC+zRSmwC2JU3huer5609oKBntmjmDTBCu
R+qh+I/HTDrhmwYsm9Eb7XgDNtD+j084Efz7m5wZ/k+6So7TH5dGCNL3a9boEA/mJdFRmouzgLV/
RD9UeeEt+shhR7uBB3euSiaG3XqCwAYCmVu92IXu8kmb7fBPq6kwEX4vh8MEk0xEwCGkoLYobiLw
VoaabQsL8eO4sLIJpxP6Syne7LryfLQSAXqc8OuAe1pKSukYPItPRFTbaF6NSXKwcGkzRhNJYx7D
NrYoW7zBRGeWZf3nPMl86Bz/2NR/8+2s3uQubG/xZmgw7wh2zYX/rSGNEylf1Dxd7AbXabvAuQuX
sAe7JZA87PpyekbZ04mjMcLua2Qj5QYprbzxcmu2ivBiiTxwzC6uirh1aRPuAJ3BHFkQYWm05CF5
zH/rNgZ0kk002ZZidsDEF5PmPSM6JaKoTjAgV5Zf/9d7QKcQT0vYw6a9/BW01mYEvVWHL1JILSmN
Gn3LQQdDe0/9mHYIQ3KrcVzxT/dBKcpqcFLaWS2K40Fjg5mo3wahkfGYd111+0FkYe4M81U34MvI
ZEissmGYjVPoSRXohIn3nJHqsil9slefWS2A1SwFnELb5ZXAZfUfLG6ALJ9gTcRbxFjbs9DsKu92
xkD/KAHqpRuA5aKmrEo8pzqtS02+hcLA7LeyisSmBaU0mnj/QHh3Fz/TvRYBYmgtyu6yZfawBctt
52HC4pnJcO1O+irJ87MgYbmd0xuE9K5Xj4w+CccMfDokSp8x8PDXG5MWOnPIwPYvBCBfcoSnTz6v
tUGigRksmc+LiNXwtlcrIJ9Qdhc4mq5oXn+tnWmV/RmoIjA9tSdoAUgxh2GhXGmhzwqJVrifspqM
IsQ7Oipp6rDkX3T9mkBpdGhNzYMF2HPhyqU+3HGMsn2PjHCYacmMKHAoBLbTgTUViWxha6lv8KIk
+YQH6b5S+AHgHy9zhNq9jcszQcaJ9YhvkIyMyLuomt9r3UnZ0ht2nIcGd1klpVqVToChS4Or6GwX
7N4BETt+xTcc2c/xcQIr3GFMNiWwYzxg9Y5NMQuQc/rzubuMuRWJNk/ssweO8snnNmWKoUn8tuP0
nDi9HXqZmcA1SOfD4LyP/jy9UGfvRf8OAupnMKWXRYD6aHNRGVK8NFGpZdPgL6SQNTQGC5zO0vVM
wJP59z6pvPY/WEtODa4tfif1RRFaYWkPTAHiHt7Jx1P6oRzodmPFVvjn4YFH1MjIWYMH4pU5eELk
+B0QAmDDZwvKkZbFkg9AWNmMeabgQPnbswXVFyn1QH8VDarQzscY1v6R+bRKSE2xp+N3lYRfTZUD
+qfLUvhMgC0xU8eAmqFrqffKz8QJaYK8FVWXIc0U95Mw9G1zINubuvD2Kq5CNgv4mxLtSXnneAOm
2/srLh2MxnroEafCnd/26F0KXglcdt7V/1E9RkzIMyE92MRPIBOOYzhxjeTuSMO8QTIC0FeCQ1/T
sL1rRQk5rcQk0aMWUte5govqhh0On+jKiksGtaIme++dacVqBxoBI0ajkPTGB/idsQR6tHcwLDXz
BYViiNKB812xpucaUIyeej9TLOpbywxIZcpXgzMQsoJF9XqeqU1P2+f5a93NgXBQxT9PiQdVN/wh
jQcsV6zYs9WRZ5JFKLxGAP/E+EtGKilkae2Q3bR0n9C1+mqlQO/eWfMFLAZjN/r5EmjN2iuHRK2p
amkJWadM7ZGLTH3ZJ+JxHgGqtclIykJ4NDVPWqUIWBe2ReSvGNFmyCDQf1WU9KauLmRSkMM+cCif
El50QJjyr/LecLKLtg0p4ekkDANywXOAZsGJHFCSWE9N5MscidQlJZKa4DqAsHciCk653jZRy0Xk
pQdRREzBlXczjfnsy01kgh1W6OAJZDP3CI+ukCP92Weu47gnSLZ3qgqTl+/T6lSZVt4v9ih3jObo
E5f/KNwKitHIaPvXb7MuiEl43EX0wQhE/qSQ5DY3qJx++wL8zeyMco3PKZvDsGBS7JC8+97mbGsM
S65s45dfBAOAd7fqL1Wyzmk9uy2FqSPeEB2L8B+M4Tf1rQ34m5DWI7UWyf7VAswILuAqNukP3iY5
Ny+tz4xTYrd0iSHwtiWAWXqXkpQSjkeNcyxvRqQxo7jJm9U3KmzCNh2wA62GviB90h8+XkrdEAko
2VXJWp2G4js0lJqj4adTaMbFFGSJablTKitGb7ZWGpB1pBFju/cW1wKdeZnYND/VwviNlITGvYey
QWPGczEL/C0SkFQuSRleRhk3rcKqbcUtV94asILnHrxNR/uPkkfftEUxZS+pGEoeOqmAqn8ezcUT
XBIq4iEd+4C5eo4iM8DwPVI2Zc0DNjfdi6+F5P5naA3g10PfKthRjOYM8sY6wyz+ZRrMnfxWRuzU
VKxLkKV0bvA9R8oATNHaC2SlnNEH5ck5nnTJludljEPQ6MkeTCfQrQhmJ+vtYSUEztCVGzc5WoYE
MtxYGHKyHCqZ6eNbyyYTNvMDOpln3DTyNuPf7lpcf+Jqvy57uAccGluL++ktFyimYuAq+EM/9XIr
/Rb6oGYRdU6/YcznfgriLyJYQZm9de/E2HUmoM5pZmMStuvOhs+z9ucagOnl8pfE1vLBmIQgjjai
qwVbjvdkHW79hpUMrBCwcn5JpFLq0CoKbxkscpRrccck+nJWHEhBxLG8rN8pgKEmopQfBX3Or8UG
ZszzJtmr+hi2VSKO/HV739d6LaPf5KGko4yCi52eqYlrLKKSH9N39ajIMP9MJl3X1ydYeuhXi5xa
HeC25oiyvZuGb50+Ck3GhVZ87FLiYbg7VDoodH+E/o0spK/mtm0Xe/k+EhFfq0T9sjswl0b4decv
10KOJmvR5hfn+dzcLbUatmcFNrfVPWsr9drwlYO04IjUF1oq4bx9IlRtRJO8YGv2FkeiYT0+CFqE
OB8X3Y0y/5FwLQoNRojc15WNheJQqS+n1JJFW6KwBaAcYgObJVt2c4Z2sdm/iuVycMGSxPviNtik
Qpwg8ndP8utbNZBKnQMDAs2CTcl0UMSO0h9JK/chFUAxr0iMZfGB0MHiQSTnjE/76Hzi8iHj9Nsb
DDj9fQRz6J907K+FVYMsTKriGOSKlaX9qqPONz9Xkzvp4zDTSJFZNLOlK2XBQftngU3TUQj1wM3R
O3MOWUgkNtLMabJ4A2CAyYy/X1tJZ9VBAmz6CTxJQOTmmsgBNvSwI6+zplPScCGds/Dk39NABTi0
bscw5DdiMHKE/O9WNWWZfDTUs45rNwJdtWDa+6hzZG02KX4AipQD22unkB+5RnOHUXgyCvfMQ3gK
f9zK4G1/YyJ4TU8zypz4r/W/G/VYKwml+wDxBLaB3WD1pSfEr7iji9F4x4JvhpykqOJDwoKi0oYJ
vzozE2ok0MfOQr8hXVt6/Zc/piiYVhJz4hv2IxgV1NAUbN/86LbOB4Cf0au2PKf1uhu5QfJXXWbk
7GEZDdPxUEypYnxHr3JNYgUiwR2/L8kCxSSb7N4reYg1bKbZqhDwOr0FKLZ4gOEWshcjT04GhISK
cTg6QGAedoHjv2KWacWzJERpDYdCNDTc/WbedkFXp30a0YE2kcoRMzZOL8Sthouf3XoxKO4JCbiA
jwPG1Sh/2AHGmx4lOnb+pGFQ+F19gcntgES5qofmbS68TULHClPSlCAAto8KhrT23Xl6mHz+NMTu
JGCseSbU/vlCSrk7fsN5BMbsLU/XKnc2ZumRjYUASFw95Mha5phONGxBjGAuuZHzeQiKR6dB6ScJ
PT0I60+2pXXHHeMG53UCAp+Zed7IHdvLwMbY4zwVZ5sCi21zVkPOEKhMwQXe5A9baCHY+ztMoO3j
CQLcoQRWiUyFHrfz4D34yoxfiBGfXXbUTrJimQQmGz8uIO7PlI2LayqLp6EfWrhtefuZ0OBWqSu0
9eIP5w2tWLiws/Iq5urBz7RJAtX+DO3UITiXpzHf/EsNHF18fqOxDeFf1WxtSk+Bi1sBWgsjWf64
0f5r2atCx1MeGTNWm4fHpzgWqCpCVMGssMCMVUgsh/o1apr6cZTm2AiC10LVy02jIbCRjsVRybe5
t4zjbU4CqNpmFx1tW6tejq/emjKLi/SYvJalvQhuiVfrHlXX2ujhOTAILZ3KkNnMqgQHhyhPIduf
l5ef5uxb5lnBqszO9uIjlpZ7V6bMyccA/Y1uWeh9JZDrOOtiObiiu0SMezL2xrUmnFImQQ0Ubqgb
1N0DxO/Qosk0r1VlcL5WBN2TgC7kiY1WuidT0vPIMIO+1o1bD5LvWwYN3ElzvAfmEajMiPQE44Oc
XI/CUGpz5HnmCfL7mMlv1/tj5bEJEuCnOokJqNG3iDlBHBdLSAerfmZfZ58gt0gTJM5hHa6GDCDj
K8b6J+3XfLSfvwhxVTGe/4ep2Gyl7rCKuz384+nYxSGKLcmvBcNgZjryAoSE+DJmomzeU75Fn7nW
hfaMaj+VFoki7Ou3EE84zydzEvJHYcLpx2Nfny71MmLtT0jUnwMKltBpP5/x2clKLlGfy4ovReCG
/PlZD6+Ro21Fzu9h92d/mxS/hQ95IsEVi9pywgAEooeWBl0xv8DMnFGyZkYlKaTYKMocuSxcSoog
PGeNaRJgLCFCK5XLJFbKFrj6xgHMcSGW48wCcZXUVmgz0z3+UiyYkYr3f8sPfQlgv1lJ9xJMGVqP
n+u5xqgpq97UlZVMWHj54zpm2Mrg/6PeoVGmYPCfZ7pnXCn58OlM6izNOTmT09Qwbx0XWgz2Dnh0
xzvrdcyTu+jrC0Gd7b/tUzf8crbyH0PwcwR3ixMOaOA8Y16RJUl/EHoT241EBY4BvufoZQncJHca
gKacnq8tbYogupDPWPp4nKc06P2R812a/e7FtfEP2w++br9Je4GxUB+fo0bZ63y+s7yYgmgSRz/p
bxzbPydqLvFwpRoXXieFF9OkVE0oyOWi5iaEtj3ARwtS7vz0vBW2/GT2vb28A5ocytHFXTS80yXp
NgzgYlY2UHAOFnIGR6h4z4pNsvT9xEJboh3Ga5iCCoWeQl2LHsAxQITvSYBGXlCVtIam5dpSt6x6
fpyqq+IGhrrIuSCcxrow8naXb9W3KDIIEikKSLa/GRuBXx6gqMxrLf5jGJ659BWXqAOsDzJZONN9
FEW5vLkWY5U0m8q4fsNt16S1S/jVlf8oy41IHzTK1Iv/S0YH0mvjiqFzpyIvOKdp1d3Ro2ytm4LQ
1HsqAfVaCrDrbj+kpCwvDSisxjFb1SHcrUrxS/HLYCFOmp7siBuHcgmH0uWABOTAXqf7rHUaq2r1
Z8G/WRjnIRmdd68K/aGzhsd6u9ygD2fUXIZODw8BbLhspq+IwZn0ohSs9mFSKrcdUydfhOkvrTkM
7RcPk4Ib5U2xYWriN+k1XdO78uEzSWuGQf69G/56HJ3A3gNce8lHpRzZZmdZXR+6xJ1K0tXLdDVp
UGbV7FMFxBm1BvXYyOfnRoID2lN6wurfmZ2AHnoZP8QAPeGV6tjaoT2RV/SY8xXe2pFDaxjECR7p
R3IPjNbOmBKDR/HBNDXoviIi5xX9TethyxReCbngtkZ/KOEdd5gbYbQFn4Njj/3sNE8l/SUo8Rve
B2qoB0WkrZeWy3Lg3pKXYp9KS8vSYXp5Pkf3qG2h13TyoEuT7X6/tWR6LNgzH6wShFY828sohOCS
vGiqaK4Rj/4HsU4Ft97avcVTo/A41A4XVIvgqNGfTfVy5GGi7hzSVMPMrkNKHxOCQln9EqQzt2qV
Y80o4Cv4ruLkguTjMx+YdWSMSDJY8w5WM/eB1v3YorZIVzZ1OpnmGK7LAv5KFzUtX6yCGHugllRo
6+aa1jdDwPK4bg9kTYVvJVnsTT7lZI4Plxa4xfQ0sKaDiZB606w+L2ku3OSGY4cbIKb9poNJ1iG6
EylcZUi+cRZRNMk0WCbWeu84qE3o5jVn1K5VN7mAwfEGN+CDbmWa+0wAYW1PnDbEiU5XMCilkzjf
MlYD22zGSAYda5kKSsMYOt5k5+hooyNTV0eDCTVKq1zl9UMpKxNU0JGxmosbiC4p3XLByV5IgpFT
mXh2IAVfV2h03zK2YnTwrAYFRp0dyJD1bTvvrh1L57eZSVaIfSNCoxwldqR8q4C5EH5oW+jssCZd
WuASyD97vYpnN/V6JlEXnJLSKs3Qjj0rTrx4y9knJB61nP4gsmGKFJSpaMql/AcUaOebHrFLi7EA
oivIMQvHQ2PIQKhfqfyNEvVk4+HYVl2DbQHWibRwMXXwFe2LDdxNzMzp3z/elEne7lpEbzus8C5i
iCvoRqyD3qc9JAXHVEmIinHSNgNe14YRoaP62evqx4ucs/LFEGSA2X56cJb4OMKdLm2YrBhDuQFG
bex1F8c7PXlUkidyeiMas4zhXEUlSi0VIVzqG3fmsUPZO7h2gtQkdYN8XRBbGxc/rJFunaEd7P/R
YMxwjuD3KmRVqIvt1UxCDlUc7nzbqU/fnYmonM9Je4yLLRrT6IHedU/dirLGm1Le+8U/YpGUYu8F
5tsRJLjZIsPoTko7928VoPU03zwmUT4qZ8skM7hf/z+fV3NNAwXLprvPQW9+BhSNGCVrTgtp9/ca
pxu5nBURzij0V8hEzRdEQvm0o1/vw2ag6RQE0O/+7duuzL855b3R+AGOBK4acwUZlFylnT3udGQF
ELmWDfZHVNg2x6w4v5yDTpTev2T9Rx/On3bS+i/zuNUls0hWYWK56PasSijhnChVQHEfdiX7BkNL
4m7ipsGVoCBGs8sS1WY/gA19SyOrKCEiIvo9xnkBxetARnyD7qph+qb1DFleHLGmrUlS0sm1WVMz
Hxs4L8Ey8ygj++JDacg9HjYLc7KTBKGy0x4zgu9DJ2143435T2l9/R2tv8MsBuf5CKR5tIIbz1fr
nZDrHSegnO9vTdc9zegBswBR5BPqL3/9KLszMKrXegxO17HZ9EwlFRFrudFREr8YhXjgj5qkg3+2
UjnFwRX96yKHqUdXDAktjtr2X0vavx5Y5dbyCP0LfjQiPJsn91Lbt5h2Oni8BKMbFrXQHe9luxiU
1dyINsWy4YlAPDd0JfiSliagjyaobBVvIl9gDAMNG3E54/PC/Pymy8drguACcdMbwlrwvRm3Txa9
OSvDU4kcZ0ijlH8ECiixCNnelkp0UB6nK4sknPKrCbAD1QPgkL55czVKFAfNe927aEM/SkPuAiT5
bjRfN+d4lDdT4rOELcPSHPEI9x4O1gwM3uVBeozk8/1GRFV38ZMRsGFDyhoSK1sEZ4/PQsTM7Rog
HVNYx9io1BaW2I74KGlSw9AwX3SMmOmAoZ38Qq/MWZLUhGVEMpnL0r+CXVSwA0QrUT99H3pPOWym
4SoT0EitKWW7v0kN1pifv78l/2uLnDj9NXTunAScnqmiuJ4ZaxgwevjWr5l5p3MOAINmawscDYOW
jJC6foYIP+kozuTQnfYXCTGXgBs1htJKDIhHOl0xqNV/teRoO1m9pW3To/J5yV0BVCaKGjrfTs30
Icydnds4HebsuiEuKHYKhcs5PN9II+hkp47g/rgnVR9T/AhfqfsoivDUrdG5yvgL5jueDXVcIRrt
A7Ve7tlapRP638AXc5EFBaD+a3wPoc3UmL3IybVJ3VauX+mxHvm7bKcpySGcj1Ky4vTjR+S5O7kC
jVgShGKlxa2j3aMBQXrRfa3ZpCDEpJyCM3YsDn5QJ1MQ+01jpExDVH8wittbKHr5EYN/O7JkrN/8
xD+x8N+hekklUl+kvHK2x9fy2xwCOXOL3mZcZoWZoa2zdSGh/KujjWc0ReMUiVXKKaAAa+tI8PUZ
nJwoJNj+tJ9aEUKSN6xzZAm0tF6NumeUbqn4kNjDhl9tSTbKTXEGgGRgZ9HQ560j9Btcd+9JrgM2
xruNFgLb52c7uLA7Hg5n5plVFXxB2pptESSwj+3Q6pn69tmr+ZWEEHWZyuHA5j0XV3e8EDMXQ37B
++InU8pS8VW67+3LJrBdvDf3f4VY1REYxWel00QEpmnEfi/ZDmeKyDEU85GlfPGCs+z+9eN4cow+
gsS1rSVowGiZKP95FEp8/9HxHxrcgBcS5dsTZwbzpqcAcMjbnnXwofVkw9dTVBTz2dxEJXenjrtv
Hewjns8Ylr2/zpTozi4NhCK4MP00Z6BXH8eFELjAOEndzL/M9Fn/s/uuRDWfiakewLlpl3eeRRiP
zzkpHE/FdCZUGBHpDTKo2VgX7/Rxv8sg6m9dZsXMPZUGkZW8B4TV+v/rnQ3hb4vW/Trvkv0ckOa6
2VvBY4V17odxxsCCbiHqfLwWfr/U1fP1tkjwrCOW/GYpsBmW6Yzlt4FHt2CAdYtPykqQ6ZOLkWpW
ibhZDlBM3WejuNzLX0ux3lr61pMOHNGu5DeqG5oVr8P7Xqzd3pNTbqXUY/Z4l4LjFao1a7j6sk//
D8zxf16H5DBNRV38idLhDOqHPOHAdNyfGd/BfSQboWIMOpSxBcVQdLv8Ua73rxLtSAmB1Q1796SG
HFH3CTA2CUOsUMDTMdoS9GEJNCy8AicxnmTda6E0KRLFx4POra6lEFHtJIVL55lzws3fXbMMah5/
FxkRg276uG+A5PCOlpMmeKNBA9lkkfpI8uAJqzePKRJ5Og5tJwHe/wbg8cf+Uj05id0pqPJBtYwB
aOsBMZqJ8AZKPFwvosB8vphKGfrufsTmJ8mC3BOtKlF+3s5XFnVpfzFZVqTJe3IeBA4TAHGtNVTx
uiT2jk71iKa2o9qSRExJTfUiDnjL22uj+qCNc13bz3OUlQTG4HeybMh8rOp/o5E7QIFJH7wAjFl9
OpsbQZ5wLRpyKsULHAgtUD2QGLYkb+8qQ/fkO5glyHHHK1q56/Moy+tIYc7qsbX2YhhKuuvfBfSs
ETqW0VxhbQwcXpE4VIm4vnkqjJpgPpLVag2H3GqL+maj/ib/DVA92mOXIZtxVOXOJEgNWmumlrPX
rq0cqdAcemmXGlOCQhoJpij1LTy8QaAnPmeX4+1xvcq5D/iYmG7pBL3NJeC9jx6l+660ozQHCplI
fVY/SHOUNZGEHLfjFPORkp653IiHIlQ0rRDZHOPjQE4JxWgSgmBHxsGVSfr5JJySIh3pocN0ztYL
71dZ1neBktmohAu8u0OhdbeiDVlm6/G5FKWRYNejlY+Xc4SZY8x3lyXQeW4cNTJ4OFGM+YvuUkT0
qnlT2tanxstWox2DZ22ngLMTWneUiyhl7gNb61Mh+630YJflYxs3aES0GM1i3nUXPP8oe7nxNWG2
9VHTX+jqNbpvvMBQSb6CPMCnjxuYzjkiLGjKFqS8qTa9e+Htpe7yvfZvY55M11fVdfzIzgVQ3oiA
J8m8qa98rywaOXOpzepXN1oxFA+hLRgouPJMllgTxId/dR8QOWAVKDE1RPo6CP9dTbsWW0iXwgS4
IY7JuzPUhtGENNf+NPSUDQNEVBI9s0hrA0+9dto5SzPCd8c4bkOd1brg21T8MWSs5KvirpycoIA+
RoMDANz3Ke0COEcswWsge/CjFt7woujk/cEKkNo7AqPranFaxZG2vfFfy6V8IoninsF1E1G6DxhK
GufzYTKbs9oEtOk7n5St4WJV6fK7IYrpiHB51J40SLIRJK5j6PDvQV1tvtjUd5HPB3CBW6DW4ey9
8dLFfD5ChFZfrDFPAPvxjsLEJfCW6B1053bBWpMPBHimIIje2BNyFcozztsUkZUIJlR8hIeu/M7s
nTRvYsjUFM5377ii9twkYgccDRYHCFin+XUu1nOSgdPg1EY8RIkw2BU8J9QuCjWwlLl45kJXW5Xr
ZAVdJZ4zDrmaLWvx5XPa7jDp2G51j45ugPGynAdTGVPT0qRblwTeps8tOYYjKMTZGYiHW6c9yuOK
Y1ldSaLIhTEyPL/zR4VJ7N4V59+fMVpPycBYRvJkMffDqeeAAPL/XyZcMb5Y3oxtfqZtT7xqKvN3
UbPKNuhGIqPK9Mb+n1y+lHP6vcj3lza1QwN7ryf27p3Kv6pQdua8/3Fj/6rA5uyJpbPfM//N7fLl
yB62SKGFZeJQSbVEIDm5Ou5FjKhT9CDytsrNcFq0ZNz5b9+5qCuf63d/59MH/Y0vHSKgxiXDw9YV
vYSube0y+8idHee+DP6L4aTI1iNojgC+VdbNHL6GsgUZ3pAcg87oWn9EdnTUvJdQX35edF932AWh
IAIE1P/XDon8LQ+rBildJt9N1u/nKhzbvM8RhEjMBEL5ZnDC8rdHWHfzvNfFQlvbYzWUJm1obl4h
2z828H/6Yt7TWM2YDQXMfQIvg/bNV7+EwZ6h5YZqC12m35WDvVpdpcn1oklztIcp/OzNOMsDzELo
nNYT3Gb9y3+8CDtJylmAIjXUeqOitVY5jzT/nnSnUb8c8Pr2lMpTEIJlSVibJ0EA5PBXPJtSerfw
OyZvamwEuEe9Jau1gtDO2znB6iVxxLeu+gzGHN8BUVIMhQ+an/pQJv+EsKXOanEA8ucqoFfGk1aj
CzWTwpnll+v62d8EpWMm3hCTDwHSq6LO8OnvPlTbmCJJRJyFcvF4Ip2f0V5yfWxcder5mc1VTUpP
RXPUH1hoW7l9XL7FfpgiUnQXJ37aRh+WkqxAquzW7Ey00cnQ+i57w0n0TBTq57w1MmvdYYirILNR
Cm8vb4x5mWE383n2ISs8xuTp2JZZDTDmq4lWQE2JrEE0TKNg0hf5ZTnUbRyRfC2P5yrDqRFvkeUx
MROBHWJoAOYnNW03E56aI/HRd3luMQQrGrWfVpC54FxcesGDr0we9RdWgFdcmzTzfmmUXuo2LQls
KwT1CZDBSxjW1D7ddjWtAPvhSlV9NuAZv3rEisqUkdmYqwiTcoFN/OlNlEtl0zogkM2GzLbuRODE
FLH5NPAKsixpV57ZIWipPPWIlLxoy9h51Y9+Ia7Roadn1rwpbH6ZY7miocbg//nz5Hrt+TTsoPoF
QiHnkJhsYze8QqHBPPgz6x7/h8U/XMJLro6MsK+5dtTEJ/1ZKMHFSOHHNMOLWwKUKjeveLUxnjMh
B+YPxK71grZK1gGyhvfvyTjunD3wgyB9wyW1hLNWqeV9Xg8AhGiWIbXXODRiG3qzgJwtLytcfMUT
IZv4lWnwfLPPvONC/Nv8J8lF5eVWUZcBHBRNTEcR9JW+9S9pf9iDq7gHwIO4/Ci0oUkqvo7JDRIh
QbCJeZsSNJB780vNsKL6toUzu79kmIqWOkfCVTyi6a3xjWEBpfphGx5p4ys7Tqno1FKztO/hb43t
rEOPNEFS2SArs4EvOEcYObVwQzmpFkd6qxUECaYRtFwGj8J+oRuPFS9XIdTfaya29esyrFu5OKHV
QWC3sea6QgY4ZqJTJzsaw4ioyd6kf8l6Yarg/QuOZQL3ZG/2lt9NOQzlTiGR4RuoN6jCNOaYQSdY
+Nladf76arYojH4tBYDxx/Etu2OCV7u/3CADSAt+dYKS/bYwTnqeROJwvAwLfdJwrgiGYww4+iko
OGf/fFD8s1sv13Rvp/tVK0CflX7TXJRtE26/L+oXpB8YUMLS+nDmhB3k+ETpc25Li22PqkRQs6I/
wilHpUy8Y/0aC/eKUGEaE0dLj5ECUIbeoZUu8nLBaoAN3CWgC/chb4I3++nVldAiHsQI2fBN1iqa
N5YeIdT/wAnf5LmGQQodexOKqrAVAX7lZN2NdRJlut7FQvEbiWEK8GTFxl7Hl5WI1X5B8mSrC9Nd
tFk/owyBGc2qfwqsvzOdvKq5LaBUX4Rm4QyxWO8nB8xD9XpCq/T2PsiqyW/jMPGcIXWxD+qCwDpc
GqE5P++A+0+8b0ykkdJn6+AJAwQuTjKeXRbn7qPEKQ1Ltsb2AS3ismBAv4GsFNuKS4bdCearhY2c
OLjTH8VwYrDvc7pLsbQEUR9Q6LumezgYpqd7hMgVx2D7T5+Txj832qnZLK4K/RQ/Tl1W+l/8uuXl
KFTV9XONTPpYcNMeKdBvsaiFRk9BqWz374l70dGkcKGo+ZAVorrSnhLrhfBjcD7YlwHStjFvxSeo
maUm0GTgQSjHuMxk/f3GXBam+aInYQJOcipDehd10gGO5m1PaIkEsd6dZu4YnFJj+9oQRrP8SLk/
uZltsokmOmMa93TJirkG0TY4mF3gnI8hM3Pj4NzDq7q7y7N6EqJiQcO3GFOCdkOClyZ/7EbBrPvc
6k+m90GHwumtb2Lxqa4h5IdzhF02WxettWEKSRoahM6as94PQxq7OtAPShDJOW+EMLcxIWxPZtiO
yAy8QZvQoWtbjZYIXQIDTukXIVJuMS1XDJwHoNTGoejSEgLP0w+dbtSO5N++TZM6lkEdk5mwt7mt
llyhhR855B0gjJYt5L+2iXyQAwF8himid3sQJI3ccR17tMT3xdxaly/bwCjBMULk6AHYbqywIj+H
hUnmvvwD97xrqXMtk3JzB1lhvQ4oCcFoGEwqRpvKTnWqj0CZQwFyxxJXHwvEjcgdVN0RhsudW6Hw
N/saPWAf1hRSEtcLAUiMNeX2tWXEXfLnt7OIBujAkgW/C0aPSYORpDV0MQdmixjeaiI0DR8dujW3
86qWSGTxL88vmDVGEA1mAGrAG0KxIV3OBIPOiJ7Yp6Xf0wkB25Py7znNMqzNDXFE1KWysBhTiT7t
vD3Aj5QJVRnvU6a1AxF5nFmS0ZlVYHNBTudr2e3Emx1Kl6kIEwKAlxW1s9XVJAoT4w3dh23kCwLS
0RzQrtDylYOHf5s89+IaD/8SdQ3hE4aS8t5UlhuhFYQ+Rne/AVLJpACElsB4AbUrq9onp23FlIJ/
eNuU3RLszjsaiPt9a+jPS3Axz0gbjp/JHU9iVQKFW3xFPqqcoc6Bma0VLsysiCMvDKuGrbVnU8rF
+3eKdHYyG3p+RG9ynui9dOJRtDMRdpvh2rkTJOi18+rIXfCq5KEY3Tf31vb0pk3XyLe7bg6DSu3M
iNjuc0mL9YW5ZKUEtsi8fsOG7eQEvU2vk/60rCPRxRDU1IM3CKnMPiCO1q0gh1ZsSQp493O3aNmu
ItUGCObaQ3cC2+fbxug5YdVm4etKgoRlAY3mG9xqbFCS5T7XxQofCHyCL+rhW7fHe+RPWx165jvj
HM2mmtiF6/c1AhUpd2ihHKi40a91BL7OMZaX4WM5F1f5hLLmZUH3iKAKDrgFUR1a3cS5SC1AfA+a
RIFac+/7LCy2HXlBtJLHgnu5jrstrK9QE9TZnXeDootqlOeSAeKZzsyS5y/VmDwYIErea/l1YZpu
DWvS27cx/pI7mjLLS/I183jbH1ccI7QonpewtHlK2hkfCdedle3QbRSFfsPvgM4igNs6sj72/B/B
/W/Bp4BArhhlBUzd81CsYnrRpJDc3sROhG+gmLmvDUZ+0aCbd0G3/jNDvAQaLlwGVDz5OXJaU5Oy
FgIlje1BA7jnw5BdXUaDxlevIbNgrQ8Kmdq8AkiapCw7ndH1+cuW4K2CDhqROYz/N87Rs/Cwv7Dt
GKerTq1RdYCToz/e8WygDi3TlHGrMav3nEzrBNwvwr2ekNnyf5wBW+l6g3ev4RQEZY4wh004oFfV
a2pyTbr7a81atXMf2djhuEjFPM10xEp7l/M4E1GbXkW1oD3GbP/0WzMCdJAjAl9sHT8XYw2af1Rx
lL2Il9iQ0uZjEfuFjJWXGnjkms6/hMUwT+AS+iPjOpY9STAr7f+hYKhoSOg3RzaLHVleV9NXI2wF
uv4gTu8pqVpX989zAJZTToVYJfc8EIb29Ou930ASECfprdrZHgpda1gOA5FaZNjYxFuaVuVH+Jn6
LEdhycUgTfaPXloUITOOyEEKSnzmdqU4Rs5ex9RpPv7G1Jw98gl/vkOC/yv0yfsFm2pZ4xccOy7E
9f7MW8TVmugc2rd+3+ZtZCqSrFrXABYDB/s2R5chQSB72M7hwqPSs48RANq3EdA2lxjqHd53OaKA
3b6Zd+iMjhloqdRU8wIPjF9A6PPb27DO8RdSZgGmfzVwcj2Tu+JL8GtKyIOeY2xEECZ4hWG+Bl9n
ub7+dtZSCtW2b0YBv2yaLmPj6Bj+g031bEEBJNmzMMdsPukhbzRa7pZLkx6KvWWmHxdZFL/Pced6
ysR7FprdYXP4Kgvm431Z/9dFAIKRmsWnxrLX0lhu1I5BjcL4YgVyusokemgkwLLFXa1Mxk8qPea9
Sec3FwG3AbMt6hCAEgjUDr5dnSGeZn0t/cyI1MhqZQqFTChVXr0aOfbi8cz4Jdm0Uzad+Q1nAy68
ne+FTmZL8467h5MC/qs8CXtBmROoiEHqsdsqF6hxa001z4OLBSURd9cboZhyfM+3xb6+eLFh74uR
M1fp4HnVYO4NG6RI2AmN1BtjuoWwtY2MIvHOAtFEaD+grPPsoxrykrnNXKv5BxzAOQ8kS6pcmd00
PveUPLZLP/4havzHrkpHpomB1vufyyidQtbL8FzGcFQ+4TjLfwp20ZWYGorCR3vOo+Ok8mkL0N9N
m0j05S9r6fJLu8aLOkjjszF9M35oQzF4RiOyF5eEH1mX0Eij/+sfVqoJbt74lSlnBYxedY5UbPt9
bFBpuPZNIYHCcd3o05/usBAOgDvKTxwLZe1gmba+CyOM1gA3qRi1TzZdJZ7s2ZQAIdfcNC5/Z2i8
VVcSTBaNmQqAxoNHsZn+477/KXzNiZpxGeOmEslu9N91BwLQdc/yoZuKfGSBok8y6JG2uqFa9yZW
9AjWGAlMwSFg2ocCNZq2wbHDvaP0st06sJKrEAP9LzCzJYk4HraHrCTRHDxo/Uk9Udah8md5WLIj
aOik0zahc5y0TIZSC8QBz46AJSB6IRM2JjgYIGMbh+WkR2fWKNACnTffuTKjBN1VJC9Gk0Ubz0oW
/T2n6J+oP9+bxnxHnRpuvtBQed8kM6sb/OXgWkDocVjH3FaUMX32iE3q2xbWXzCBX7an0hmslIG5
1IV8L3UHBbu9JAG8L0BVGgXrlgS8tC0DRAL+g4ZVQZYaKaLEQdnLonYpsYTTiJnz2Q36LAT2oYQB
duR/88ISdJNyUxZK894x+C47Uq2Fl/s8Mb3/Y5w8XWsc/rJNL97plQ8qdB+YiNDtKPyylBkMVCNd
VVgF2V0tej5OhT0t0ZWZw/+DgVxbxVU9gpZ31xE3Jl/VVAAYcXbs/kq8XbA4XGyqYNmy/bTTPuOC
TCz/s6ekLsN43Q9VTMXQuzt7bFGbF4yiOFzBSBkBIwwGiypTBCuSJ5/dc7ySsEI4naSFxzWFTElH
u+i9DbWVLmN7WzPchDM4VpuhmsR1ifxodMomK33+lYf/o7RKOgWl+B/aTrLJAzuEYOA2lyyZ0pu7
Q18tv2sjdCLxocG/ZiklPRSPbYjqi6lnpQAc4RGXvVtnyEPqC71rlXO1xt1l01JyR+s4FhAkvmO8
1gVpgu5VR9n35YQKTVZ23ATABCfzxIgCXF8QEapYyBUJmhr68cw9RKa8M9BT7d1vhCHDQ3T6Ihom
bZL1MjVG6tK0VQfWiePcLFcdQ+nGIUafgdLgr626uKCKLVIwcfERyYfw1JscNQ3jG7cwgjP7H2NN
qmNp1DOS/R+SUPUryfOsZxS7mun6WeTDXKK0GDcR+u/swkvv0+gdAPHem2LNp4pZHPJ42Bun/YQ1
NGGxwcnlKn34EYmg2Ka7YBVxGxqg9LCvlC760zLSHd51F3T/Qe0h/h2E602sdhpRvOK3pYoQcDN/
jgZbn/n8zbGUd2pnVNlkpf4LxGmzzkdL3CB4Uno8n+tRWr5d+vteRVBdlxHxX4wS8wRSwxPTeO4D
+/zyeUTWDZPK++bBMiZk8F3I1ZG/xs8zVefvR6qL7Cgo/pWmt84kRc8hmgWgAngugr6EHECQ9vzu
SPnzLgoedeGSBKD0nRsriZGJmg+8PSb8tk2SwNWMLQ7cO5LCFyJtvjLYsqgIXMNbN7YMZC3nkw7A
83WiI6c1ybQGzsIrLQKpr5dPZOUMG06RuXankDt747Eefr+jeGwPuRdYCV2ohboMvmnbI2Xcu+FF
fx14VHsj/lKn9X6Vdxh5G4wT2jUK4RSbX+4zdQ4mxN77AJQTGZFaDVplUoGY7diCkaA5zpC3u+s4
q5ox0RHR+y2d0CjLvbpG5wSP+RXBcFdlS0vATW/41w6VA1gSI3FiN0Qa3jJwMqu9F8+9XtFXT9CD
jKH0Xec2rsba9v3OEJ/rjD5iWJB35lP2kNpJQRJQV6VHynvC4cZt0tH1qFOmmmFGvESdUzbCrtXG
F3SIMm+LRERkGAGMqy0Ddx192hEiN0qCyrckrb4Aks+AyP0x0oxU5SfbJvwK8IhaHwT9vVFzns9I
hYs1hT9KUNgsvENb/Adv0NwtIEkAkM0oRtXoLPVNi1jvWJ+pomGWYmMkaHTYsIvBx8ttfu7NYQNQ
zxdWjbt3/+Ccysma+D4wW+/8uUL2D6f3cdgf7m8lYztBIT6Wvi/aq4noVUQ/TewEI1OfvK9LndGz
mB90WYeKIZfwGMN96R1+eZiAs5toonyxocMHwPXrZeqIJ0TgJnxEhaikMBi/hao2clmI0v6pX6hp
qoioVWTlvWtqvPuqYTb6cWq5gsbzKz7HT64PDLHbDtXdfTAxb1N5s+mEqH36n0q7Zioqdk8jW6wb
jMgESc4S+tJUnBuhg7x8prFHPqD/efNvwKe/fULuiSKG4wcivsu9MNNE34q1OCZ0JYqtnTIHBXtT
31qvDzt5hVX298V6FKfEt5INwehiOzsoW+GcQh3RHfoJUx658wNwvFWQWE5yNKeQjlTRdk9Kln/T
pelnwn/J80Avn3kS8iehz2CUWfJj9jEAkpngE0LADPUr6OB3Sl1VMFWtxBAPsclp1ditZrfH0mPO
hgdP+aN47QeQVEBsx7YdFIfLJ5me8RiKdn1/gSMccn4UYr0QBdo4kYxsx4OAtZvJRdMK0ZZJF7Ks
rruxKFyzTNaPD8Olwe8vvoJuXE/A+IOk1f0RSAP0BGjaY65DxfTPPcjTR1MbN0eSnp9RdERPYOgp
Sqh71Ls3PB3qbJrb6pqS3RzT4BKbItxPVZc7RjMqYHplM6nePFsNAmM1MFR9FJYloyjNzgB0hxvL
qACsA87yZ9eUVs4/h+sgujevhrZaJwiR9QyMRVjCJ4b790bmwefSetL0j30uBajW4rjg3KDhBqmT
vTDzcD6atzOqin9nLX2cZAhFDmDFbNmvhux5LT1pcMoRd9sVqdAONFN4AUcK4V0EwMrGB52b+py+
mjf8PQ8ElkzmOpgfck+3zuJ+OpAzxSdqk1YGCAZw8x6y8h0pTvwGu3neg9dPZmPypSdbciHkYm5x
q18H2ZwG/Lva+jq9//VSG4Lt8oc2djudEY8YsaYECHRf69tu3wHgIoss3JNX40+HRX1Irt9OJyUa
dX7ib4BS5VFNv6g2XAxK/xodal9hPWGXKHh8q4oFQiX4O98WGb7+Uqii3RvKozxjFS7v1Of4C662
qUfNFez/ULenKMdrQWEWYnARddDqqXlfY57MDxTcjgH29zkUP5umddIfx6rje8ZgaytXKTcUzNIa
LwQXRRJRh+54LJuH134v8plQLa1BOrYH5uD2PA0N0CAra8hFDyPTSDf1i4t2QGYXGybZcHTGS0Fh
tE8c8ufFYK1T3IIXuVqcnJcH2KdPstrLNZAQfVwx4zXIUGRvMnwe4PqVceYjKqKtTuoUk/z8S/X7
cLhLqrJXmxc41FAxPkHjkb8sjliTDuyjFGss8mjvcj6NRt+kjvYXc6LCTWY5D9jJKouH+6LQFnNs
Er4l9ZhQzXI84KwWDTdgdjf6SnwsHThRyYk4JpQLD3xV74aVwEl/Frzj+J4mH8e94vbtsq+9+/Bk
au28KWFqBythZIAVzYTYX1KMy/QJr26B8aeKEHXTJUiM7+ofyW/ENUNmuh2GnQF/D0Mo2xOrZtzR
NVEv3IeppgU7b3EULGMEFF+MqYFUWP+xm46tfLNPppNJ51s7ltY8fjyoeXdrYkdT0/zDgDBVq17d
YypsqcY/cJTB1SXiukIcrSsLgyT6cDNCfTnDVgM7W9XcLAJTkqAESGSbf7/KUL4O9v/oiYnm0miw
Rj6jbhuKM+wDit1z9ZTmpOYzzzv92jDvRassiQytqOnoNH3a8uk9NEI1pjWVLU6augojRG/0hGwg
JSTvicTGbBrsr3xWFlDCwrBt6goW2OVxT1HzJU+biosNyzpYxKr/FAFHxTmbFFg52vSqlseBBBoa
gtCEi0a+cFZotMVoU0NjL9GdTg27gICesmztzb2I45WMl/dXYSQUf0ccWQ+8283X5S20fiUHZETs
pc6mIVurjRtLytdCtk+74H/Qv1eY3BabPd0LvUKPsrxJE2WXqsQgBV4FOMkIYHqulO0pVHIQXvW3
wT7MCqYZV57J7odPHeRcOBHpJsNnbKezVTXU6CJVwbcudJmkTtP+aDb58ZOtLhn83//R5+iMJovm
S8t7uU6H/FDZBFWj1r+tH78b12sB2tBw6NfoH2gN6miyjhB3QMeRXHm1CDzhsbvoNp0nvANNQCWc
d8sEI1wRaW63KVhvdmPcSCs42wt/mTCyQPvnmZgAg/6Q7QLe0aqVWA62b5t533vACwCyEUJZ74L6
UWtZXxjpL9evY3YSQXT3AfTJKc1G56dQ2/j7iUFxbADlhbq7tknTsAkrz5uzI44Gju3SpFEnpmHL
Fc6hXnAa3zPiMW7ze9R9YCnZ+c8vtWTZ9JqEM7+jTjwM5pWAaBRWxInVUxGTW3PkQppyHYWx+vvl
Wswxiz3GYzuvF1J5FCXQIL1lK0I2enbaRVvqvuLP64yNX+W5M5kEQJe8ZqIE6RJmDpdbC1b1NUqD
NkraENx2Hux3ctMFk2AwohthZBaV779BL3+LIojW2BIqRxYdACLO1Na3yk2h7EO6qE5ksBbmWAb1
GE6rxmCNR3yMOjbWy1lCgUITTzxH/l+T7bACW1eyEmtBWPh6KcVkQyOFU/b/HBjDV+oqh3P0nFc2
duFw4UT9LPD9RI9VUJkonx/b8kv7Qlyqv2J/TMdgpbhwJBcIEFtkq2ed+F8dWb7ByFb5GiCAX82e
nmhKjac/wO9qEEhhHY8A3FubsrXtxxf2U/C7RKM/cotVHy9Xal14PjmyNjABTOkRCMFq4YFpofZ/
4OIrTXQDBLfbpBV+oEWkUO6ndiDlGWGE5Hdc1LFkCVv+qKia3rNugjo0kvtlaOqUn/WmXF02Gb0L
X74i1fOdskPRV+tmOO/68Ov9/uUI0ePe9WuXglyXY92s0Adcg96HIbzlIWSEO+strlz+SzhTJDVS
b6esmr4KT8gYfpa/E5Z88Bs/xI4ptC7aXldLshGubAAzikupCihqVx+WS9LLkEcvwJwptFIwiXc8
DFxALs8fg5z4P4CdMFgfPb+vbfdj8VR1Of52UViHT6DiSKrXOrA/xB7c4LRb+6nzSQPtCEg8ZM8Y
yS6yLVRt9ssNZ3WSFlAXRyPijG4s2JTBCqMhlZ/90qO13EKxH2mlXuW1xdn6goSnScofvNhNwRS3
DwUGKRom354oTAh6YlL7wD0pv9xvq9uCt1QQIW0c/cvj1v1viPi60RF2kFQCeI3jO4qwwOs+sJAb
QBbbccsg1yt5uHuPOrKD55m2ifWrneA4+2jefeWljqwnm2LJOvsy2z7/IbMjv2GODy2Q5zg6Bk1U
MSYVbrcySojZu7d1NBRzn4+6+RqVOLAzYJXIIQOIQM5TD+mhtJ1vRovagLuOIj33CjILzFXes5Zr
o3JbAC12d0G9H+4iYqQ8cPGCnftaU2WMHFDyT+jtwz5yielsZaLeQvgmkDPcCxOTt9M5W1ehN6hb
aVdhstdHpl+XtXUB1QCtx8L4A5JFvedqGl1Lc1cD41nHw+1wZCIe9iCI5P8OrkcwSI066C00mhcB
xeTOAG/vLGRxnSEAJs4Z7y6j3hwOVTviJDHs3l6zRVTss659n/7OtQbXDgAEyY2ec9/oTXId/GZU
HwuIl+lUP2QoXxQ+1JD4+fxcr4JS2vs+wr7kvnMUumJOvUHwALrQeTklrBdGvk0KqgTlV+omRVYY
Xi7y3VQKh2qpHpRMWwgcV/ho2EwoMvWNMnxI1JkoEblcGWZ652C3bJiorzrdYxmr3mzAeat69J0z
q/J6bq8UuRxMaV+Cn59fv70szyZS/FNaDXvGxUBQc27qktOPXlV1HCo5ypwDL09gD37KLh91sbOF
U0q4/eXqTXbeeWIfqP8xOr5PT75sPyQ34OAMKiyJ3GwvbXeo3X2ZlJb78B3pprnV1tuNM3Pb0rQ/
jN0DlMIvfPEBVCDdO0T9Rr96lXym6B4tnQlrtwQqOCdtFXuVHruuYGG1jZPdp1mJwY3zsHrj/3gP
vBi+/aiAO9+D6uv316zQZ0RIdAelBPkJ/BTLxDb3pJwnV84+EP59Zm1y8u83iwNPxUJeOI1Yzw/4
/ubN+9SNPMN0fSJwbYgYu9PHyHNXHZvatQ9I/mVShtVZoZCvRAidwK7xc9XOGLMh3XZPJ8n5P6DR
Rj39xXRG+0xBvjB9KhRMYYJPsgYsjyFwGaYt8ipnwfwMR5kuN+Nktyzs48v8yBtTRz8pKQ9jF8UE
xU2gxg7tZWInUl1mfYTQtgIh9SDXM0iBQU+kEj8O6+t7WYdf+RcWkhsQqhd566sO8BZmlqJPhDVs
m6PH5hzInKidFwTR+qg7K7vEDoehX0EHnIol+KT1oO8jgQpLwG3W8QpCzokagY9QI3QIe+R0M/+P
H+cC7Ak/7lq0lbyW8Gh718f5a6l+jJ2/rLrwYScv2UYuwu+5e8iNXHXmmDA/s+FUO4WyTs1KmJPD
GPuRkCvhxYsghKO41Sc3Txs9Smofz/305JU8ZU0BOpa4VD7oEEMZEh4b72axoUEczf1q64yhhwBL
zKI6iuIg2FK07U5Y2xbJ6OKKN/Vbw64QW/R3W0xedabx7v4QtylZyxdb15oMJUnXutwYQh6uNdzM
sp+Zlf/F+UQjD5NRg/9uK55PIGYMbR2T3TRzPb9Kn4CVs+5avKKNMMzItUBUKX7VWorazSOitcx5
i+7RHL+YKZgPAVx4B4fUNsZInHiJfpVISkBV1k8n4Uh4GTFxg2Y7rQbJkEqLpuzJBfcsHDTewD6l
YppI0uXZpZStnXpRejcpHA5250Ve1O2u5E1nbrjYNXQkVVzXCZ9Lci37+cKn8F37MrR21wm5wPwA
eNHs5MBAzbsPBNVYIF79RmbIcuTzBA5p2RTn/20yShVSWPOsEpAX0GTR78FdKtN3p85V6PYzzzDJ
HwWkGTHk5qb0vEyYTkjfS0td7u+jzeUwAybWKdMTx8hnbbqhTHrSGXo0+2aLrDnOjpFmDqFDmXzY
l2aPKXrbdojOt8m0A4W7GksJobaaHujLRoMEZQEFmz4JFaunmt/ZLqRxSzHNSiDgnwxLeGGdBSFv
u3QuEmdjaEM08SHR2EZMN/hiiGWXE+YqJ7Kgeep1ztfPynW7cLaT650nYmFGVPmjopRuUqrcNqgI
fx5+lZhUisFmt13A/xyMrQ5mnwxukvHl+1dtIEu1cBLW2M41KuqwlUPX2KArFLoR8VzMruM0FHqO
DIhFf5B6a0iqcfHlmrIsnf/CefzbsOx5vMnHBt0ZPB133EsIh1yi+Mg2qW+MlU7IvewxWAqBxGKL
qOjhdB95PD8G002NEsYkb3lpXXnEnRFNcC1Up+psZZ3JhvHHqzkb+zE2+XrazQWvI+Su2DnCiAVD
8CYMRfLq/HJoW8Gn0hxnLSdF90HoPR1nP1ALo8uCVQT9KJxzgG9LwHgTxJ56PAe+O56U3AkwqF3v
KUoFgkBkYHQz/LJgBL+vlq4PbcSOmyjGf09SAJMTkfQ8yywDzgQT2bB+RgfcHInwsZ9Myf46L9vQ
Nv5UYLQQgXSGsDSqY31b1HfVBhgEPX1dQLfgprrgklGcW7YN/b1Wfy2MnuCJA/f336zBydEHwaT1
LoOchLpJ40Z/wDVjcoVGjX7IyBrCm5APTU1Z5Tz6tp1+pQyXT54+/XY5go9fIyzVaOyhTVxruGL3
ERiBuJQg07cdy3iZjCjwikoDNSIQ95u2GECvMKpDs7G0iY3p9wBDERxSrZE5r8+IGhRIDAFjW0SP
+8cGW/tyEBRupr6WJTjZv0JNn4ynVf3GCgR7pjAoHL8tueMg7Rg2yAe0GElISZrTV6Ts4RDV0isI
fU8Q0OXGbQt0RRcd2+93/DWeU16nyU02HgEFlQKpF58VAJzVFJutgjeMg87ZGddjLLamkZ1FAkE7
ZQRLK5J0B0qz5uhTfaYONCI6ZkGKczZahaXmBG9dmoUb3c448z6cHeGIWWhTiu6LwPKSv5z80Afa
jxF0MM/dLkQlTCXMFn/07ErJMHclknw22Gk5T0+loXk7SWRURcuBOXIl/z8x6rhLJ5G7EU1moAt+
VI3kBonD4dbY3+X14Ya43PzG+azIGeKiHLloTW0/wppuqeTgTPUmV/QP6k5XOWDRO1TdzkKDzJmy
XDWYbJVGnq+g1dT1EY+AcNntCVO78QWRUNDxKGFyhgOuPopx6lcawbm9oDvyCyY7v5TprYxZisC8
9WdHlBaQwjw7EaWed0s5FfzVJCUsTIbjUwLYPHBUSwFb1dKPtQ3agh6Fw1HeA+PrVkjZIUpHCtvB
w5lzx/xNE7VfoOZH92OvzoFCiV5Enc23WhN3yA0zPtoI/u/o65o1N+aIDD0ULMv18y5Q3H7v8OTI
f9CxFXFQXbKa9AqNumxkONkNn5s/JnxzfnyM6DZ1Ruc7txH56spmrdh5xaCM8yMdWhihqf3pNwYv
tn/wmqwzfKTLispcyogzYMWaQbj4sE+C/91k+hfm6M+Il+MkyoMW3w5B6xNqcmPJfvyE153IbYBh
PR7yCIAaS7xxW0a9rn46LiASDsT29mpceIbWc8gYeJ096rqoD8bxjG5wOoghoAmrNdDgs7c+/cY4
mEY+KCh/aXqj+tqW7MmipsnHFWLIqh8OHj2ZL4QWFPShD4rX0kjvflh1/7yyiF5DNPExdTcJ+qDH
tlG9UhlHVY8hvYdLCotSavyIz6ycrWZrBFwZb21eRihXmWtDgEWaMFLagu86m5Iw0WMuTZh1uc7Z
8cz9ZTF+mg7IIY9N6E+DgMkQO/Rl4MCvpJKpjoPXrt3Qw5Tts3jmFh0L++Go9U6FlGWqbApXqmIP
rQH6QFMEugzT/WhjsHqggGe1jmdVL7NE0k4gETEida0FRBj76RfLXVReCBTXlwIIa0iwTxAqRgyP
cxVBS4lHZctABtrIxp5TmbsQ8S9hnM0ZYC1wVKUTmxcaQUAtdkrkXr5BdiaW50/BvOMEY7fTqxsM
e+BZlyT7smaITYf7BqRikaR6vdyQgGKs4fKxjVMJH+HtexC77gcgbzFo+YiDf1O08ItcFqUDe9ZZ
o9qaNmHevbDZQypXuF4l0MXpd78WX1BDYBGDY4+EONrXFNNekoA5H/hUhoxNYGw2nOKNEED0idqO
O8r44sciRLOE+ixBpsViXRAPwgNuzwbAIcaoVE8UtfLsS9J78dIctdSZ/TxyNYRChOslp/pPA3yw
qsma8z4nLTijqQYhKyvVG3V86z0vhkI9Rsi+HdqvSwPQJ88Clc9SwJfs6sfDjEotsBx4QR//yw6O
Q23RUVoxEACe3NYchMszd6wnBsYL4cMcM4WJRjd1i/sRVZkrsfmDcv8N51qYYjWOPY/T9+TgFjCa
KZcKTBwphCeyU+C1ygOL6OUBMNVfn4YBP2ACg1ML5h+XA97xNK0d2hFksrEZYErMAPckmeC2r4U0
Lkk2kYQdY4GGNnT3Q1b8qkIFHq5vrkUY5ClRbzTXzJcwFaxaDC+lTwrk1vzHANf+rhwZoqRDlk+t
nm/+qn+eWvfPzVRWAYvZgNmhqDyhz26dDjL7iSf1M/PWSq4orJP3oSLxueJWw2K24sdFRV1GS/bf
Sdm+Zk3D2q8/ajB3EdsaWLJyIU5A8kL2RtLapWqK4oPWcG5csrQnB8cxwPtW8kQ8WuHDQFd/esYh
WG2+0sTDDMsAVD0DOMYFYkJqv2+AE+eeu8C16H/jV9yO6duTgZ0Mx5+3vr0CrF9h/B/dw6FBSvQs
bbM6wNN7DHsembivB+hdMMFOnJddYTMtY0f/W+j3x40x/uYQrAaXOIfMHTn8YhPr0Vr3J6CK1dCE
y2qPkxR2oNO2W1tkTzV1i1Xgbm/UnI0KHPp1olFrpXfjMVP76160HTovTv12xeB9hworTvb4XLYc
+EEPRyc/dRT29QYvMVy6jgQCrMYmj+yh608BWPau0FeSnSHOrMAejexyrF0rjS0XsI7Fm9MfGGeM
phmcPI9mmGHaPpmi25IFnGRARQy6fKdj4szLfztWCAY8GZwxVEpakRj4S9NJwk7y+RA2TGPMSuXz
5pdKhueUh29ItKV9+rUVlGthNJXgF+43vOW5pk6cXH44Gpjglk5Ak4D1wBqZoW4qU3jl956KESM3
zQeA8i8joQzaXb9gRJbBJeOogggsXZxtwyba3oCjIOlcv9GlvabO/7Ypt5tDypP3mmO9kzJi85Sg
UMUmVsBndWYFCMPqbO756zaqVlB2fypl6xjY1+t/k5vIJYEYzgp0NMT5MAWiluExytU7NkDExZ/b
B973S+OwrWkjcg5xqREDFboKwYFpzmG23Pze1fmSwACBBmVBwjyNwAwH7H8HCFOhs5vHw11gXb2I
8m8a1rV37bifUo/IRhg+tYpaw8JvaVPNjtvc4bV1iHlKgIh06fsFrmx+Nh6ZR5Vq0Uz7bCNPEQr4
HR6C+LVEenKqsb5XeJakb2KHc0nsjOMbSPtyGdedwYCbCTRGyRlswmsfAPd9QUh5+oQplo4Sx1tF
voF1AWjSsmeGknZjGxguQ93rVmdibEifilOUHR3zAxASk6qVDoJnQI1puCURUvpwDkdee6S8MZ2M
0cdlpZtU+p7/G6zTKwhWS50nTPtgkEZ95PCQbO6Imrt7BeCsTOIkFkKL5AyTqalWAVQ4zENc4tUK
NiN34zo3j37lFsSrY8MgdrzaubCT5HytndGXiOODhPMgjzIfI7/4+dXrwaIB52pOo8yCJEP/PsuQ
UXeERTbwaU1vfCk2Kz7tIX4WB6hf8T2pDEYLzSDVz7IVu7oyyr/jknSCd46iV3g+UzZVyqX5HxLk
N2WEVT1DLlCKflyb0gKEG8FxiKNVz6AJqRUDMKpmp3/8jnj0yXbENGBo5s0J+V2Ur41MDz+kNykE
BInnva0ZZeJ59mxPTAkmApNf/0ELMHj0ofx0A9tegV5bB6gUV8dnaNE9uygTJy3TuYcvVMo+dkW2
UxfO+XML488tcReylz0nbCCY7FpIZSSoms7NryQxdCiswGZHmATbknqUJtvePJSP6ET1+Hlbrheq
4FiwJjbG/FZ1sk4LRgDCt0FUM1XU4+UI+5H0MJ1uY6+PS4QPhroGDgeTVF2iekAEDHfOA620Smuk
GmDhNxzVnL1Xc0v6xCznM7+KbxJbUJOMd4lV1dr6X/u1+3u/tbwbHZEPRZjolth2BFoErhF9nSBJ
JpDNCaO75uaoC2HqtnleVhPbX88puUTCPAtpv0zjc8NSs6hIsgOr70mkMBXLNqV1atymLza7yLvr
gvSKpZfi3CD9gYiZLIPbOdwOMDnu7OZOKkgWenP0pkNzAEpTxWbVp9lcCsTXv0UPXHwltknkDdbA
uVfxhZI0fDuBQGcDXGWEfy4PpJstEkXERKYz1wuqSDlTRg1RDYR50dQvzFg3OTR9+4Cr99bFZy1h
+rjAY6oD2mtRhvAxU98YopduHHsGmFvuj+8YcxWuv0ZsZDFeUliVRziiKglaD3jZoymzxleMoNr5
88P31cnMYTOEpRgBaS1Az5UXB1Mi/cp5N0OvXbGTrIYxgf1nLtn30569bMdjYyfgCV8aG42LRIE0
k5GCBDa4ovqugQKHVKnoPaiVZy1MK4B9BrxjAI7dZ/gx+D2BY885kfKLT+FUltSg5ClEwTZ5oBd7
LJJtsFKYHQdKSiPbtO+bRG3eOLntUleg3LApJdo0SGeLX8ASixtqC6hgMIqnbUCe6V42ZFal0NFz
jXQCDXlwHqSeMjdj+m9EKqPbSZCidvQet503GwRO37XDnM/ND/ZX1cDcJ1joCvfN3J1/7az4lnHS
IZ8eadjd+0QDJl3nMFQKUTphNWWcJNDX1+GCHknQbaizDDQB/SL6OaBUojRSTpS2lLPIFgo6y4Gq
tsWD1G2m+axeCbMRTgNc0RzqjcvdBGT+Hj1gXQ4DzLODU/VUyVIFnJuxdF5ftlnym1Q0fmo88PaA
Ih6bsk8vRwbiz3MO9fEbhq/Bx0aiF2vsEsdffCHfe/XkyaExyad932jvp5SwnedfsieXZT9aDGCz
U0ADbIJK9W0juw8I6GMLQo18yLFiB/1kLQsOrtY74PIuEL6ZAwDIaHdM5WOyj8PocZJwbmdZUN9j
vhaZC7G0mXFN5AjNRHbSo6+G/33wJnsQnVRImMIFNp+fw2VfROSXBRN68jX8L61lK7m6kjDFo7MI
YL434RRxmmezOKwasT3PD1hi3gRkK2r+IUktpwQE4rAzyBFZcdoXFgCON7aL5oLeq5ZlFq1ra7PR
B3VBw3wpIFn5nCy6ZqJCN1JPcpQqKVjvIYJr/Pgvkm8tv8wwXe1oAq68doMQWqt8SnXbYQR8HaaO
Uronftb7bI2EDPSd0qkf1OuUHJw3eO4N9ugw26mpemkq/HnPn2l3B+/8pAHAPzBJc4uWLYH2xxO/
ky1ttDtoqwOhcxzUrgiX3VVejyXhtssraFs1w8+ZVlC15Zwr1Hj6ZRvcNrP7Lbh+ij6npatI2UC2
W03v9s+yK5cBzVCeP4NB8hpfwuhBrCE6HrVYdj29LWkZAqaYIHAfYE28nflFHP+mfjLRweXyYU2E
OIDmtLqBMSSOwG6urbCQtRFkR5ra6ppuon5rDFL7Aj2tMyUFAE5P1JPUWEez1N/UxTzM0UuZBcOv
sElgC57Z7ED/jhCONEBHjewO4TOJwD8zgsf+4S+nS1sniAY/V6sADtH22/Kf2eVIAgdcCSKl+6ro
+Me6m2OtSyAJvn3yKQU6I4Db6fF65w0esIKkZShefnHWLXJ3tHate3Wy8wYpx5pTTm5bwZr/gALC
16b/gHPTQbYC8J2b0EPSa4n2Bn9bM0eJ3LPwq1wrkXdZk5FMFFGD1LMI9PBExIU21oqY2DiZGM83
dbXTM2mF1uNa2Ht8mraQ1vre+/akqRZ0u1JAJXxgfMnx3rjbnzKvtNMeRw12979gjglsUVDexs14
F717FgHNcw4Tv8zwYOA6yW+MPsreiOwkQyA2SMnqCzUaPuzfgowFZEZ7e2kXif29LMv+wGJyAt4t
CzDaIuFOCzzP2vTK7qvxIo9uxQ4Qi5L8+gf2ei0DE+18Y2SKyOjMgqxgOYvDUVVt6HyfRJTkq6Dq
unybu0c3NJg8tu7HihFJAxEDWE8MQEKe+s+pIwN2klimp/RV+4QsF8la+98dMOTy5EA4wTSMISvR
SUOKHXzP6nVh2SRRYbs3y1PyDCIf0ZjufZfrtGVE9B150NeEXe9T2atlqGzHQrYduMEjOGAwsXYq
lWXhljy1u1dLMCvoz/nAgGi3SJH0diJuPeD6s85w+IprsuyaAXeWOhftzQIrqgv7E/4LC7Zz424t
umMfz3nL/0QkTk2A8EWNeiEe1UhRuZj49A85IvWVTvh2f3Vcf+FBFfwOZXv2NnQeDcJTskFQ/hTZ
IsSDHTs0+lI23+1CCXXBBH6SiQb0sHvlmGZ7+hca38aIN3qIRMuMcKaS80YYxfMXzCv/21gwr5ej
8ntN9EZOkbhSJ65a3OYBQNWa/xkeuFU17hIMBK7y2Yzi9xuGa5TWjJLRv6pduNtGUfCFd3Na0/zs
Z/FN3RK80fnSWE/0b8QAnp9d9j7OkwsdGQEjKxxaDLVdOpuDEDkA7xtHfm6patQU7aQCCxrmGEO2
mOaSjzKoMvw4uffchvTRJn4AvZk6X66mFzzQS2mfst2RumRLTqiTwetB/CnlYCLaU/QdDv9zmze+
Jh0V7+fMCf0gYGikMnMADbELoJ9nY2LTsSY7UMwK96Z/LN9QkXBJXglpsP6GD6e0NnxHqGn6dupV
zUcJKixlqo94YKINAPAwEuCsohzrzoVifVYseOy/l2hvER5Kxd4IZoit/Xb9hAhQ0HgDWPeI8nHV
SxjnmYPudHJtXXn6Q+TTwYLqOOCGT4smp9xw2ok8I1U09xnFosLI6qRTdQNmWplxRWFpwNjwdyqW
14KvKkXP4IaiatJ26QJDDCdi7RQUnHjgzWMC18ir+c15GW95q614vnxzuTQq36OOi+MocW8xisYU
LRAEhvyUIT8A9EQmhk8wdl7K0XBrKyBIFe4/OM/0U8cLIsnLWjgZXy1a78spMpLbB9qG0MK6rCbd
T1ImuX0CQOqvcpUEnYSK+DErD/9i4COQ6IbM6S+4Cu9TtwWi8Mhl+EhrcrN/ffi7S/04GNnClLy5
KXpCAvBNMl+zihMFX3qzSxd3WW95mv/sGZWWLSLK1FkIqg7H4q8FzMP3KRX3KJPxC0TyYjztS3oj
LIpqrerqX/IwTx8HWzc+71F/cFh83ezlqQ4SZ4rrsAXNkleQqzQRCONVKbQ6vvPTd+HS8T8J+q4q
hIUGVPjkTTkxFYBgQXeZfqFbnuRCCy/FjZWpsMBxpzsOlNnLjYn/ou/YoHldHPFTeW9C5nlnzt32
iBPmRFZ9/OOvyahR2dIZ4Tk3cOlrYzLjlyznIBu3FjulKBC4u/UADpIKcs813HZGF5NgiYSEQzOU
4S7r3ZcBxqTUsfP0eUbk71QgF8PZz8oOoJ0vZdd5Oz6RzRc2OJKYXuHhgJJTtvMBzhFETNUh7K30
aIWGGnaXnEncN3whODej3BnDWgekvyO2XAh+pDEeoVQ6UTYDS7C+Up7hQNGVXy7iYi6A4kWTQKGM
R30xmzJ0OBkBMsGtF6k8MjR4I2s7D5O8iEekF1RIixUDRAb0xhI1sa9TfiSljrI9dAxvfUT2YjNq
HO55kq/4pSqUknmT0fItfGM5UugchRlQG7hIHHoMncL3s8IcWLpDwN7kitYQ0FaAzA49j7MPB8Zt
NqPdLoMWSklmcaEcWmt2S5RdPizyODTeZ+84yuKjWyDZ0+auk5mxVSZY9TkDJL5ikq5AudnmyOQD
GbbXs0q9p25ybRDCx+pp3aCaXE0nmWxGuKoVhXfDBKpaZJSleJr+u/x2D+DeN99PE+k8atac80EG
r7zJ4LVLW9HiLHrKUY0Q6GljuEdZho8EJWrB9tyKeh9FNjZGlFY/vsAnSjA6g5XWMWmjStzNTCyc
PIZohLR1ubYQL3aGyT6p3GogBjJibS/YFczGaErEAK9QLSfjcfwuTYxCyXqYgimpfLq40BRaQgxG
WE0gu5LjSjuDOODzKOZCmyetx6pIlTg24ctR2gHnotv9Um8uL8FfcPUzmEPk28QfvVcUYpvQYD58
rmoq1mT/FgJf0si7FyQ7KfhYi2zi75l991HB16fOSqAr5CrFyCH6K+Drm/3DGwOIdzKFAnWMr7v3
IPsMQZPZds1FCRaGL7XWPvW1/YeHd4KDLL38BluPdNTkpWVt6YlC+BzWUDsvgV0BYk8O2/Lm/xhK
DHqrHtBn9GnSGXbwK+5h2sl8J3zRbgrSdrVHWB3RHNnpBlsG2K/ucfZAwKtIUI53Ae2F0/xCPD6l
Vyua1HxtHZSNYY5O3gr8K3bKURyq12VEEUKfp36u+kXMOSavQttz5gOntvWLqxUmPKjGGRPHd4Ww
nsW7CrB0VlwiwriuwGcOHYub1Ize+ZvFE3kcYFMXPtxL8wkhQZttoB68/w9isC7vRSKPULvnNbWX
a9QFm8O5EQC1Ga6coaComXpywsloBaFGQK/kwOuAZosIOGyb7xzp22yC11dE3hj2e4ZXOeoo1wV8
m8eG/npnsdQhJt6byy/+kmKiDWKq65ZidQ5IsYMdxO8VYuPAtQAo2WPHWa9VHX+yeZYGykewvCSN
oos6qaueG1zCUq5VZpvIMG+Zf81SM996THQo4xZj5SYbGtYtSvA0DWpAKw3Wt+HKZh9IiH6dFWhv
p45UaXDicmFWk7oMo8N1mrHMhJBUkFisXL86FZ3Utm7SZU9lWWIwEJGpv3JnqrVZ5oKB9kSXOfY1
grGWvZHOd7B/dOiThrLadB+eltIaSMqRZ+lnjyA2FQkptHLGIUnEcbclKsC7dBddzeojEdI41f9G
s/+Y7L+7pCMpq8Fu6AMN1u1Vv88k0g5Ok4vMqlaEiZOP0+anTFX9XRib9zXI0qz/7j4y5Q6NgIzq
A18sPUjwx28LkcWwyrwBrbf3TPmNGxpmkGv17rec/RSE4hjpSQxwttCmlQC5cThiB++//EEEFyyo
oOKjKG2/+UQ9ujl2cCIoPRbj+xEzi64mLPkRkOqnEPenvkRrugzSYgMHRQsD2nX+a1QF7wylan2w
Gsxgd9gskpItNwJsB60B16nnjMh0lbC4sJEgNGx6zfSK59OLaOoibN7y8JWVsq34kjJuK5L/O/uT
3EO9KIVFSJXTL1k7Y2JIHp8fyI2yDPNOdZi/6wxGXkn1Jfu1PAw0sbg1xs4eV2KIYX+ioZQfdv1+
I7dtwSsr0/hc2b28Tura57LWYNgrypK/nQFggwSBDLR5uMZ4kH/NvBg1NRUc2Di0Gxr/22smsuLX
z2HBoK0P7pZAQ1ai8mQ2uelJcaa6Aa3jPL+mee60r/hZEFsezvzEwa2AyQPXMPr8ulqEXkUwT7Yu
4JT2qOTYKGx+3iG5HyPiaoxNho3vkKCJvwbdASrYS5UxKTmBfnGoqMZjZYuyX9sILobaxOd3+4Lb
OjKWMWvCjVtkkRhY0Wlb/RyM3t5C6r/Zd5xXHnaoJuOK2RYKZmklnwbio1iuQcbYwioPvvmPZc7N
xY7BiMpnEIXwHkWfhoqCSRF49ICnfPlI5CXbgOYOCAlvJt2GpQWGsusrxnZVyuLl7AQHpuTVvHnx
C8FcacZwX1a7e1psbcbKVsRtyiL5b4zxJ6jVIYqotTFe4Eh88Nl2wzQ7wZY/gcUCUnPsuXSqVgHX
Z11NzZmRZH14BGcIT1aFD2QqVC15X2m/Mqg1GdONR6sgwtlDRhQtsvtBAM3Z3Kmc3IfCJdk2TxXO
EQAuW/Cd0apSWF11tFOPkagDOdTh+1XBAgYeFIrB1A9qzLq8qwRuBTicqhPzBYw0dfIPAr2D+0D5
yzm84gUB7+CUIut9ZD6D3wtGoDvKn+X7C/Zy4mFKMdZozTLvRf9yyeKFm09PrGUwDcJslHO33efi
fEMerGjVUWLABKQHasFQ7743g+EvUp4s7Jq+pOwoQnwbVB3RUy401qnZkYj22yDXfN+Hl2juFDDN
kycVmC56wbaetdK+lqeCnhSlkOHdhVfZENyyIaOCLof6A7ekSSnXqQ+XgwEZJg6NbvinBzSUM19M
t3nNsGQCYphl8w6859R1RN1WvbtaGSrFi94ndfdVpPF59Bn+EC03AC/+NdHaQW2D39dY2wfJHX1+
W0JR6KUy9OeFoPvP+MCdeM5QO3ChMEsb16BDhklG7gskqXm8HyRddw/zdxSMKem0sdR9ICNmpm4I
b0qRYCO3hbqDF08fONAbl/kFBwcHWwkOxHVu94zKxWZp6VghFp0Mo8VNYGM2zzhy8qfO+mxlLGnk
A4L2cfHV29wAgai8feTwI22C3f53+9exgGP2FtO9ou51vk5Xg+6RBY6tR5TprsYCoN6WblbVpgaW
Upk2msW1n1bj2hnLq7uB9AwiS2QPWEnVT3/OwNb9+tqrqxnUpY382CTU27qdoQfBuGh4XyZHhI0H
6hXPGT2svWm9LOBu28+YWh7dK4IY26+vCYrKXtojQbtOiSex79FwB05JcP8soIhwlYywBFUOQuIp
bM9RghJHhioR6h0jQLeG/a7Kh8u1s6pz0BpGdh1SqWBDCzXkrPary7DfAkmRZ19/HS2QHhd25vXP
qXLow7pa1BFRSLY9nxIDxYwcsbrPh9cIZFBNk4DpeSkW3UuOCdn+vovHHx6hx4DAC7iqgrOoEzVi
17oREHozaQwxZRytLd+eUkK9eM83MVQcimKqSojcf389Plq2qjv4jMP3rypSGwDY69RmMC7Rz6Fy
TEeJCX0d3O6LdVRFKNKZiRW+ys0Wef0qlVVNJvg6vb4CZRA3tlWQWORmf7RAZG7HOYx7YL0Myz+f
8YGbZMuYPE1Sse8Myh7OLdP4uo3zBthP8Efhun3BNVDLt+TocUh9LPq2Hv90FVaAZ8SSMKdoR554
CoOAzC6LgY8mjUB7j1hD7CC6IGNSJhnGaVoxLCYFTCTPCnN1Rgpa0SqTemCz4U4HlIGZML9FSkag
/dqkguE9GOmiLkfGmHmrM71sMILQ9Dih/xU9f56OFoic9OZ3qWeOAD3EU/PYfsX4/efXk4IfDrEH
ILp/tercCUQth7UvEqjX9v8wws+diIhRFf4wfmuLyk55whfCVFRDl2a5IJ8OsGqNWe0N2mcocDrd
aAnVOeMWdOiBZ84eLdJdwA4kxcUZno/X9m32/GWRd8z1P2XorCzq8vsNp4KQN2SDjaq4i2Q9GJ24
qfmRYKxFtoAi7Y8FGqpXi2OC7hsunHFReYSMVIoYs/0SzPUyjIj6CQ7pWdZgk7hsrFsSYHKElQl+
WZ7wVLSrECaXB7rxWojTxlfyKc2iuB9gBylcBPunfUpkO3Zv3OFnQybOnBGkjyn1jyTPROY5HI5J
KiqsjpaBJEq9OTEbWQ2RXYjfj0zwTL6FrT2COp3APzdLzvmw6C4PoG/aBgRfM+VOh398b03t1ecU
72wd2uGVnEQ/igi1OOVSOi0HMuqb720bKOSiv6neeKI12lxP/S2pmdHHYZmKQStq/asPZr4OWmwO
VL05uT21j6p88BN9+pzigCm2xdm+id4CdpcqXaLncag+8onfykybL9w1wRy04OXJeA0Ro2POOgu/
U34xsJIOX3ymI0xrV+tBEUJmxw5LDXC3oFONai0teiaD6to4ZGw1RcjwYfMBieV4qexEQy89ursc
BSk/bSndbSSzQyvl+mKvxwA2fdcHLfwIW0SsefgM/+WLff081/lWsL6Wtce+UZipQcDtV50wOSyn
by48IGQ144o5dzlTEfq1PaBFZV/hxI2uTJLIozOMiKizsuvHh6elZCinCuPXoR6LWxfgFVYVpuSZ
wW8VA7CdhsA2VTochfjZD8x9juD9ke75qGOloBWjDUbwSwi74BXONXdhFC/L65GAoXYz/YVlvbTr
i6zUs2uc5+QFFB9Nhvy2+Qw4tn7lWYkgJB/b8nElNdIF/q+8TLjK14GzmrlgT3UPwm54ifNCgs7I
pLJ7nMBqafaIwWCleavU+R6wMAfStPskqdjqrPX1LaeKRSAMz09PPRZR8JtwS0Sp8tQvjG7lgCXp
Bkajpho8GPApzHGcdN7dd8oLN5BaUVwWYpqsOwpMCsB2PyRhNhHCgl7fMCpqTL99lfuzXxxZfR9L
/TGcmVv/1mFwMM1+TF+XI/+LzV7HAiZjZDn7SOsEl7swg1XttzsleHz711k2u2W1+OzM3Chmt9Sm
8m0jzhaa+qCpiFdj6n4NwR0F6P9Sdxe2Q4YnKmv1/lo0VyQSGZUGRk6tNETSfKnd3dwIsX7WabZM
P511aXnCISYmhT0LFcM23MwMaGWfu2XQGQir4oQ79fMw/d2V3iju2qPm5eMiTaKlsnq7m6qH4BUH
Hui9EdWlPzovC0LZCjQtTW1/FmLSv8WE06gDrd0vYASBNRGKgP+VEVc9UExdhPqLkR8wzytP6pF4
yFeVbmVxpdN8ccgfeJAIy00dnMGI0NJr4xO5SQmMxrVZn7jxyUpTHhtcut6xM9S8xMH4Z6EyKySi
daqt7U0aQSrIpEon3JmIBmxLxjnSIfkGEXJqjxtb//IYZpUgZb0wpJ8QStx0Sw11UP0mGWQgkDZR
+3VTR31JsVpL00nLTyLaxknQyw9P95qlLaEXv/LKV7c1oIuuBk24ViJs1pJjwFBnkaI+xIiVoFel
cgi2f52kCp7P4es+d0v5CyUuo2oTVgah1m6WheJqqH2IdFdzuzJ588eDWUNtxiS1ljRaUfVot99T
i9npxuhXWTWz5we1WcjknOkbwKTXKCozjZHsw0inuVEYaBPF16FpkTDKUyA/1+d/UgB7M0Foew/N
evB5bh9dtB2nCcUup4iQ+C/otHn1OLzt0u+s5e/NNlom9UruiqcLxcBo1KpnFiajB+vWFXApFOOP
56Om2NNHBQyy8fsr/adGu9GR5Mm7YapKmGgzFQx6DO9/5AP22m3lEc3VmYXIA+zUJxjnfZzlg+x7
2yHKZPN0dC2XB4aPOQop6oWlsJJdZoTic5IYn9QVZvroIKL62Lh/dbng4hLDUEGys/UifXWncDMt
G4SHKSttKRHGm20rZHMxJ+o45FLXvpI8H/oxbFt73iaTefYumR1BlBAKhH6EN6tHZp3yLMqIXEMc
XJrxAtiba5A9uoWv9PdOx4C8rRGEExF4/6zxtC0982/4tJcndymXFqpOA9CWWacSMavUI9hWcuI2
ouzyDY+ZckQkgBR3TqABS9yZ03bqlr5BwbaKc/bR94c+VdOutE5rqXkMOmtOiCSwHxwwz5ZDEZUU
FFo/pW6apNERGevHcP8ZKCMlqxDQvyrRQHxoXt5iLHn+M4///jOvewaBIJwyfMRrrCFAT+WrDHvg
a1TUUo/DNP6WX/LQC10ALzvCO0akltew6bG23dxPaC6/DaSa5c5dc02K+4AIn64rmKxz9Dtm5uMf
fEDCk9hpKP18KUsQz/Jgo9qzeKJoQbInfMvWtBHB0bbtSVPkpl+sgDy+fFLjCOweH+CCjMPlV6i/
JccCmmW3tXIGs6Jyy2ezh8Xdj5sQcmwv6viHVK+ZvQBKurNfqpIM0CeG/Wp0R3cztDyy8s0FDAV0
p7/8v9qFcE2iXT+rdGAMfGqWqZqzWkDfeDQdnHV0BxlZaldKyWbY51+ItMNOM/UbS4blpSQXA4Tg
Xyusfi8i+Xgr0lk4lLWm4FdfZsRhWSIY8qqvyLZ7CUwu/WrfxKapXOUPp4ti4+6gJ6yWsLgmx+eC
03rxxa3Fz/9Y4KVHibZAln5nPlKkN6V+YGDh7lBU8vpdBB/bbXvALlla2wgX1ltUhGyI/4rxvMn3
fKHHOXj1byleXIw0bPStjDhJZ58ZNZFmN1+fUlAgt/Flr7zfyvMhGuK1n90gRzSMxw4e0DI4w5Rj
5NX840d2tPiSEDxSjHj2cBDUxoOdtT9Lb0cDo4sBNH/L/x9h78Agch47zF7suQqegquxQNUQ1xOd
OI1jGn9SOfxodYaZbaQxmmSGFf26cUsJ9jYxFHN8Ha659iLcg23SmAxrsrVsuJGxh1/8BEduUl+C
8WsVfu9wDHbOjmucrIGoUE5M/7JkTEri7NEe2kE1MJPgKifmVByz5qnQ+siRQbR7BjfDhI00Ro4I
oc38wMr9xUml5+eoym9EsqjdjmEE2FeImM6/+UdxZzzgxzdyDa0v923TY2Y4O5goHMKf6jJjhStE
vmOAp9k4HTY9/LCTSWmyjYAVlqAUKpLrut+J2kFW2Eb9Yd6m+DsxBqoe26z3R0f+KgcT1SDgKv36
j9wYNcet2/UTjK/8Jng1B8Lby1WwhPPGnTDmmac8kKayzjJNYfGcqOL9PdZ04/PYXG7tUx0hx94C
FaDZExp+LVb9fxdZXzDfh3j/l7gdIJy7Ww9N3hrSkY/Il37gwGys4eldyvHa0+MohMKyJFwczZbR
4qBY69XugxBs9k53XgYao+ukMDP1yX+OQGDcZUfuCHFaBT7OMZOWwb6E7nG3L2WGcRLwVPbXkLhy
1obK8ZYa+ZcPihwm/APnHWepy4g81Qis+zh8bMQz8LzCP9PKkggN2LSRLdKbBMAKJxKzJdcgprm+
pIuYGh68AggV5WzZC3DBcSmOZfbo6S5znj349GEml8xGzTpNo//7bso5MCImrzVib1PM/w+v2Eh7
kPmkfs83UVHms/QJbYhDFvvdaYRXowXIMsO4aVh+jlYJLzchaVgBKPYjgIBRAYPUDZ+/C4SS/axT
xNd9wV29qYJEyZ+IzYMIiTMqeaL26VPWraiTKYBauJQlw+T7GUnqSMwjJQCsMkOCOh3If4EL9fNM
c0ouiiDu5A3vQUBwbKqoeqb3d+dwVJYN0RwwESNDnU3dmG4nSL1zM8DA+N46AbUMMNjSDDC84KVk
JUbM0CcHBOIUdU1wbjlJJ5dG84F81101cvqqosZfoUcNHGT8D8XGeBmQjN7yoShJSVLeUvjRC3AQ
i4VzRYloHrhEKXsaUvvS/5KLTu9NY09vrY1dxVhGyL3tkg/shPfEQyrwRFKVltt93CxCoOkmdnFI
m5I3AO9rbxa7RTm0mU85VK80M3iMMEy5VELGVCg1c/UtmSipMOfB5EXyUqNv2Oele39Cwi9PoDQc
TN6ZLc1z8j0Ncga0P9OTJ5Z73YeR6xahZo/UOyN0jsSE5C99KfGlx7+WRtvNiru/UVVNdvAd527t
YfGHx4lMwnoBGekQCLsY0Kv0DxDANAXO/AjKz/ySNZWN4dde4qsAWvotVEeA9ifEbw/uBcbcT9Eg
YZmTXM2RGXMAp9ZLGKMNXeNUySsgQDGqC3zjE2PyEo+Rr+RIIPp3pCIoEvDlGUna3YasQN8XjrYS
WYmwtPbV9RcOfcJwFuHGY8x0wffw3F7gTTL3mtuOizYv9WzAfI1CXHQdCf2asWa0yxaygOuQKruo
QVxxZ+C7HcBGWB6FVWaFPNCUzigCMMNORxeRnO/v0D7x4Gu/esbspoeogKJWn6T3votUTQfPLX5B
ptMKcTawjUPTJmm54pPZKZgym83wIzZkxGV5udtb6CdMPcv3+CiKKvxrR1RbeBiXklmEj3fknrZ4
YKLDmgvmq7Ac/ZWPnQ8cVX1yQZ/TlaEUqiZ+eZ6+HyxX97eLy1J6i0tydct+6j0KpIH30/NYCMMX
kMrPPEOEzDSiQcnaG+oe9vpH/2JLs8jvtFMYjI/WgzbrGSvvGz3x5XbL9yQs456uhFZpCUkkirHL
aWg9eOVPqeh2v2JJbCuCNFfgaiTa3HIPVkx5E9Pn4LSZ0lRGBXSaphPmZaF+DTdOvtfnQP7r0iGK
shZcUizf/A77jrh0CydLQXmLdffuPSFqY0z6US8VgFZSUQnECNG1Mm44yjA9oZGFTrB1uuFkCPyZ
gpEoa1XOgLi2eKmC3cj54gJGlIIQBJY93MwLR/4cO1UjPdJkTA4jh1jkWkssVz4SVWhD1G+JYYBg
Xv3UgLKKVZQMawPDo76UaCTUSO+62DapGOvCpBlGw+KHn8PgJ9Ujq8GZvRmqs/I4Z2UOrDShmuQM
Nk3xE3wBX4kOfmYml+/jm2mItmPQ9bk307WuWrfIcGPaMKKWAPnHshb9RCoxZffadqmLx/e7JsEm
M8K/hUz96nGz6L+m8E7lgNH/Wg3IsVPXulvALJanMCF7aAQfxPHFEEti9Ob7ifVNExihHcBhm6ty
tEcFgKKxamjk0q6aRNi8qFOXb7pfWZNeG4vfNXh/WWGcVWL4i09gL7saFdskktiVTr9sEZDdXuYk
D5VB4+nDZUCIUmJGtQOv7eIvylGQIe0BDa0if8frJUZyAa3dYw2OYG3dVBg60NNJj8pdAqQSZfUG
i0IeRjfwoUk4DlmuXz2nxBvNKmsVflllu8it9uzHDi4XNjterNkrV5RVQdBz5T9EK+VQaEMXFOOo
JDnz1NQ3XZSc4AS8qOhDBEsLZWFEozVTrWZNMBEBUwc6clGM0axSsE7edQJkEI0dMgXGU7+vWtQ2
pyWcjzfYaRhxymHeroPV9xplcLKFiKOxDynjO6mvHz/kbaohlwdOZ3LS0mljNauRCVEnM+Kz4jpu
NlaWz9queKmycaASBWWS0RUrzYTeOriw1ZKWAkIV7DqJyFxZ9vy5g0TbVmkKw3pC4p2F8PL3PFdG
rQpDtcmJrUET+5xFVqrEEeERC7lBGluiqj6ydcSD3llmBDXCnx1gfDb3/GfwFLHMruWUkDLpPc6b
VqMnyi/Lpt65czZGrDeQZIpRuRHcCBqwOTyuns4lkPanOjSBh31BZaOMbdmyhFn9BScxNS6Bi5XF
ffXJj+4/2id9u5t7b5TXn2p9039WtsOKXgYPdnbj5lEOiJnzmNi1XeMqq7iprNybWYfirwrsbR3C
VQ7kVcjoclZ+wLKXVDFmsdgjsFQaL7ZmZTzFBODBsUnlBXMSU/Wkc3s2BfwhfjMnXjGBJ5GOr7Ub
VY20wVvwp1HA46tzyWjlb+XlfG/g006B9+xi2bEHil+QWwjIH92faA6LwiYJxECDRCT8mzgGNmMf
6iAPf9DJt0DLQvqiDPNIHjM8D0OgqsewWmwlZeio+yt/Omn2BIO/e22N/u6Ga1TUYAmbYikJo1WV
hRyy0Q3cLJ7lJ88GFJc4QZFVDTCEhffcsyfQCzt9w59cozVbTQ3thB9eXqaTXPDgXPRLk/yxsZZ5
zs1bsUFq++KwHdWn3+36yGtCjjlFR/l9A1Lm9vcbsL2aOfQvcSlbiBWexTjz7BCxPKgq28ZQ1zNg
3YfsktL3Erx66zhU2PEkTmKBW2At0ErB9BeJ13PoDmcrsuWnkb8GshFF8RF4RKgqIpWKhey4fN2k
zswUQaJwngNdQKm73LO6jCH5CygKEuSN8rZx/UgBuNEAqY/spveHOURZ+SCq7ESjkKAAHl9OWDBQ
2g0596hhN8NxZH7r+gVPS2smIVPCYsx916mlgTbd99SowdNgKYKhCdCdMoi4KViDU2j95CSIq6Nr
tQ3CTMaTutfcMXw4R1+JHZGDzdxOJLbQu3fLivY2NkUvk2rz5qAoBOmdYzKnuXfS2hg18LWSB6YM
KzGo9V7a8oJLimyfB9veZqtLEY7Eqr+gaFqpE9ymZroWVbv1PZr76+U5Vgwz3oZGRkzQEAUuqaIw
I9XrXEuzXHxE748jcmoxqjN5ttcXZGo3Bxsups8WAcn7C1f5cJpd6dU8GsZvPZjMtfUp5XsqSd2A
ioeQOGvLdMFKGYqeX6AyGcuzZFz5vaYF9vpTCR0T/4xJPukYkRBaEfxAYylSBFjVWeDrxqUfvBKW
xv5gobXqC0pb1ttoS3jCYbc4dVJrNhIkfH73t0LcpulIbojMdfKes/6nb4VCoWuQvjvy7SiYUdX5
QlEYLX1Ua/WC/GUCBO+GukTF2KoimixqeMjLGy1u+lonaCgyOYYGBxouGNT6rF1vy9VvRZVl591O
2w0K43YYP7FlF++CWoZMKzhAQGzTXrE6B5khJz9BCD0DFZWYY5Qc5krqZYcfg1anXLg1aN78qB2/
7YblUGqtGyE6M5VUKwntGgjoioix/htAfZs1J7SwTP+XqvAb3Xf0Fyxq5xQ1rSMlxTge9Sgvi6FB
aQFDEWYQvFVW3PsAdCwEsW3zrFrBdZnUNYLCSQTEa3gWUEQ5ESkVpCAuCqSvAkk1PydR4AcQN1Ve
63FTQzkOzatnvUZxIPHltn7hlS1pUU1vLQjurwvffQ9J4xel3DsudkIFkn4bNSnxF7p1n8vN13Jf
1s5HQx2TNiwtxkMEJjJeJEgDe4l+vzVBKguZwHmo0aBVqGO+RQTjDgj/qKG7BfV/8Nku277O2GTo
KSr21YKvjjDLlNg56nDwbhiLhYhrjV1nc+uGOqmSijkBeyjFLWVpJdeenTYBXHBv/XGofuXo+Zut
P5Hl47oN5s0xzZWRye2Lgaeo2iBsBgCl2OQZ3fXoKyv7GyNgI3T5TdLNxBf2HhwcDDjLMPC4HFB3
BM+G5iSDTmIRBLPwUBZG0xPXXZ+K2Rj2bP5urWujR8LipoUcTKBcaNm8oWjxm566HmGz1VO9BPcN
B0RIcAz7LvAhW6+sgQfmudKtuhrXQXYKhxGixdl2BE4vqGpdCalWlkjlDL7+cGFExpmiwe8gfvUD
1wsuwqFKdI1Clt9pP1jt5ybhzLcLU/SljAph28IXgfw2RgeB+7PMsmdPYkYSZQ7nrzZGPIKeqKGJ
71qe6keoo2lhLjO8JE4PxpUD6quO6Lh6K5J+bwrSA9VxW7bNofSBmuHtKuVKJPTdm+9uhC0YrLeq
BrdZoUPmIQbz8EYSNzoMvg90CFTDtpeWJin1I0jTmEjr/hcoZLCsvfdQJR6DE8lcJCJLjVrfFQnY
k4J3x7575fMNPvWd6FYbXbMsCl9ofZL7FBPtE1i5DnjSb7BpPW72SzljkrqsttvJyA3wfHTx3zfg
YHPlVm1zlK35j77g/MpHNUd7NW1sp7Qi3QwdFGWvfVzaoMgtBPo2vOiyKFHK7qT5OnNp0p/29Ye1
ghS94hMSggJoDo6fb6eafz5hq55Iz8wcaCy4XaHtA9iki8TSnYN1CQTUwEuLHRhj4QWAruuWNmY0
RroG5Yvatuj1MLDm/3b010bD+n7bBpbBbZKleW/bJo+1oYLA1ukyDupDVzBt8YBEcyXSmYLUdCOm
tRy4OFaFPuWBuwpb3jitOngv9g+3ZzeMfU+79K9E4lq4yXxXNfVYYTqcIegW2DJGol+MnlVgkwnu
GA+CQwSaKUJoiAJNHwdMrwASir1HmcPXWeEBn9uFzBry8RjwkQtfkdgLSvVHHb3bgs+ZQ5tidCjJ
gwLOEQYF/Ujd96wjAfUItLtcSSSiPZTvdx24xkQITdbj2XHarwxqKYWr9dQGKngTF00CZ4lwwXs5
Fwn81PpclCJ75k17/Ib0W5q5nYwu6BHnEEDWL7Lt4P11YMzN5Rho/sYt/nBlG0gE1BfakkZs9cfx
NPwrG9/rCiDIAsHOJPv7yygAkJizPaT9D4unEqWlGYtOsxcExJqk8KjnJcw0bgCPnGtyByuHFsxE
fIfQfupmH5IdqEReK5QcTosNW5BJTNcDeu5BnMvki9FAD/Ar0pX+kZE2J1XrEl/SsIdbXtS9dEzP
2Q9PXdStEwppJuhHSXVlOAYk8EUcE8u4WeNF8q5M40yCvt7+Uk7X3M7tdNlszOayuZk6x+n9S+Xw
N2pnL9mYl9lRlrzXnS9PSK0WJ+sokbq63j4j0JO0s1sLrnSL3AOBGzzJAFZLRdnohnVtu7ccQ12a
TRAkbBIPP+8KFAuz32FaOM2n0riO4XMyr+mcEIaF3N0cYVrbYE9BWdWF3f7aKISkwMgfLThlGQuv
ppxXC1LWE+yEJ/9Pts/q4cvlN5OZN7fo+qVy4yMtrLi7IBWWdkwGaed74U5mGZa0Q0JK45GLxZ3e
QiHOR5Y2nYlXxh/Kxh6FdRHN0mkEE6Eh0UaAi/b19VTEjyY6b0uEQLiirF2A3raaEKuu4JAg87O5
4d1ZBCcsXVT+EYiXdlvGwawkJicgB27VNuaoNZiR5bh0bCKpqbGk+F3XSqcyUy+A36+GCl8TznmA
7jbop0pJd08YgrRKDvn/ba+MluatxYCDSQNP/bCbpzmYaQpIGLDWHKXXnSsYbMJ+ZnHjtA8QM8WZ
nJ+kILktciCWYdqw/ysmCsqVKAfzSpD7xWdWZTpTfYPKPQ6GOmo0RQkv4QZSIMhDfVpkCfLy/wGu
EPzBH7ROrM+zFLi2HpD81fYpojmDS4HrMvplktp12vNNBOPOdZiIeZd5LL/66gXJqmyfXHD5LwKN
W+hx5fwIyJdl5zfGTNgXC/Fp7q35fdaHuS2Tr5fVtOKEgy8405QZ1RA7P1pcxq18Bn3j+Lr7tm9z
kYh+nQM2WjN54Gqg4YrL64FT91Zu2bhwKlVAZ5iADCK/MTt/VpoN+b/sRbLq87iIqi+RA/TLLMr/
VcMlRFl2CmmX/cjF8ze+YxksQkHccdtaJVCA7as92w8Xar3TpEfOjDUjyfHs4uqOhvQfgD8YH0oA
i5dvm/HnijsF1TIFRa3U2bCuxarY3b1pevVtiJaMNH0VZv00iwzjUctFER0dnDty0KRhg2z4pimS
kBxfB6w6ueUcn9Ul7oPB5itDY6tbLhF9fbnYyZPEQ2Cd3YYYbDp8L7iHBwWRqLbow8C1/MHlbbCG
pul8lUnUjFpzhSYwQqf0vgu5By1xI4Iz4TlbEdpRb0uJFoRji1z02wkba44hOAY1RMEkI/oxhEzT
/QCJofY22egxXedaZ2qYMxfb55Qg8AzkiYrJAsm62kCXbd9eSNMKGHMyfbt0bH+mgQhEIQLMmsxz
mxduJ5gnun6xZb335gnHeu1umVzck2SjfjyW8hUK5PHj9lHaqj5QWid1dbS8G+mfihJNXIs8WbD7
mH3XwKpkg9upf5UY12NctJjlBAWnkS11TSif6rHqUFnEi9AdGrrBAygWZ0Zs4+eH8uPmfiTPM5Kx
pYnNsX9XxZDzMXKSEBN+b9HhWw28PVOZ4gUfLCgA2ihKHvqHDZX1O8boR2q9/bHXcAUiUfMp23iw
9qd1jh9t8dAj6YedPMLmVfcOA6qIxUWbTLeZiy58NtrEgVrizEXpVL4fTvCmTrP2iVmptzENETso
VXPGYfdfAhKfgSnsyZA+FDlgBohQeB80q7vAOvGlirj0tuTb3N+O9Dgoj+cCC4ffTvxpJMR7JV7F
H/wnaSNCeDHASxOXRoLvuFbL/AeBDr5YKyBiBpEL3iCkVpKUUrQrBUQNG4RZ6N0P2t50JT2dI/KP
bxGvaemBt4WA7xNMgcPiE3f2r+SmJMALCDmFNdZPm84WHhXgJRezU/JYDQ99W2/XICKUtVNF2KZA
xplHnBT8IVJ5k2Gqt0iAUmGSkKcwCMsmVCUNSUN0Mpkk/JyOqYZ3a6E+SSjgAxQYmfQEeXRsxQ4B
jz57nnE8pyEUXfsidUxbIN+J39iuGTXv/KV8bwqGdpgipv4B5CWkry/MeKqKMZ7kG/Kuz5Wr7zYB
t3OwFrwIEEIfO4Skr5zrG73DEwWp33De7vXG1fZx85FCkXfHPTzFKbeBCENPCb+EYHV3lgOgikyz
DT2PHOi2d9aFbM6/7F7vHxT2snNFo5lv5V7DNEjyE1sz8iDcHhPs6hvZ6RG6N1uzgKlHdODeD5zW
+qEUJRtaCNek+trqXxyc6CAxIYCUdqO86sxeEbW8R+D3fTD8C2p5YB6NusrqI+17xqSMKRvakDsK
19+2HtLFbf+sne70SW12TQyr8xhnn0uM5A48Dypq6w0A9IMQG6/c65LHaAesxpOfXtf6wCDww0TK
esh0JUmT+GsFS27I3LDfpGdbbIld7Yd7AeOCbHuNrFOm4lxR+uBRzZeWgo/7E3tuQb/rdjnontYn
4Tn950MS89Wu/3/AijSi0zmrej5hCVDLloRDoLisd2WpxLxmhI2oFBPjVRGTZ7zN0MTHZjXq4NYJ
2wHMeYAAOP1iWZ9CGUf2PN6t/sKwt84yjxl9IjlyFCS7ztEZsCGrfRDPzxA9a2wTt87j1reReKAl
AMJyZ6kwGxC/QNiDTg/Ogyyee0DWuK/Yeu9vf3F5EH9+MTZcNiqD+bhWX2PjEKLi775iOo3QzOaP
HA6nO6GZXLXZmuv0RwDBQtZrWV9AY3qpihlGZzZ2k+FZz9ZtflHag1B4VSlFtGsg5MuaJG5q29a3
71Qgv55gkGZzIJ7L5S15hqw57aoJhUCM1qbRQ3NUp0yMdowwPElBIBsfP4/QZK47Mt/7dcS6cZDI
QL2NCyP+BD22qk+wLihrXbZMHn5vsE2iUadrBYAv6JSLu2cUoHYRbf+uogqjh1AZtfWneucfte5p
tWfzksvWaE0oYNxJUk69MoCpH/9N8XuxGPxYpZ6j3ZosmbYPNb8DbKWIvcmLhnPAN9ZN/d7o4d8n
buQ9GqG+pe7xA0iczosCen0122eJ35vbP8Re4JMyt4emhjB7DnsmgrZIQ1K762RrpRRgHK3AmRzA
oUIfFyBpAq7sMrgT3skVAdrtV86WUzteNhNL34bvw3eONbMQQ8OhN9+M1yhAsUJ/HS1dTOrdeCAY
ZUfrszuieiwhkAckwhUREHZmkPKQ1u5N+YWlikGByUOEN1DNHunBZe6Bcx/6JxLdB6vfYVvlBk/V
hgi0yGlaVBNfx2YJRDB+WHn1YvLO+Sd7DQErMFnF74Bf/Czo8OBID3Fog2wN4DN8bb0KbIS5XOAM
sGcBEhVkSS65EAvnFNmepxGJVfenD0NPJ9hFyLB/HjVX5ZSaVWmJxIYv+jC44LitDKMyQIs/EpkL
taIj9kIbZyhoQEZ5nzbLQEnYXdyTzSbT91NGsE5HTXeOEN9QZSsBx2TMn/AJaGcer1owMqx0/NRR
QBGKKdqS54l6TeoV28yPGPo6zcgmkn9esBldizkU/lccUZuyutWWhfG0DJgGJ9chKLMOqPoLyyLI
nv+9arWKY7aPX8FFGJdmu5rAV5AC5+9hQyvFYReWBhnD9woC7gT9erGAAukdq0mIhK5vyfeRdrlX
dfwUxIYXbdt4p+kvTlRBW8WoN6Wt8hnd8B8vv4p80llcHRW7HNKL+8wCGmkdhcr7v3hfd4IXEKKc
LL1L3lqNgWQbkUDlivI9o/+eLXyXCC3V6Lg7RYMZcXWWbH1a4WacqxILLeFo/rK9cFDNLVFujEA6
s2TAfvqfB21o29bw3JY8SgFVF2wPxpBpmnAcJjL0fwc0aCFm1Tv9eNkB9X6qw6enB3S2GTCgSLwA
G3g06FRHNbKekJYgdrZdN+UAlwXNYTYRsED6lcoMScI07fsRRN0RNwlKpSLT/73fwHTe2npBlKoZ
Q/991Zwt3jIV/GY4DxAXChDCpdbwpkqaq0DefRN7Sj20LrrKcsDGBzfh3BAHylfxNQCfJbnGrKmE
vsuR3R2/fnlHesMe5aE70Fkc41VL3r3R+FpRN4q1g2zl4WKszcZ++nJiFJnQTW7SOoNXbaF5FLQ9
BThU/o8Rs6dw16/KR9hBtKZnZHTy3/OjXibO+BEw/WSJZBMDVLESNkhymhPUxB9TWKLJbifC6qtR
+LlXuCorS9ycMsJvs8OSiKMqy3truc4t1aI3NOxTk9jixl3+XTDcCI6s1MLalPW/CTaWogq+qx/A
jmgE/CB7a4WGQf79KxlwTpkYVlfMUkRfNdXPduhoO/7QEvxQPcDvV1Ggux7Nle5Spm2hYBeiIZuG
H+LQFyrdU2b1W3I4MOVkaekPLLnGw7UKnP6d5R2Fs285Hk2kkD9MKoYCebRo/s5eZHAuYjZ/mjlg
2f+wZJUHgKZZZcBabcOnEabo7sNS8yfRpLBGFEmk4r2tQIS6fTHHTmSbl9RVieEGaseCUaUd6pd1
3qwSYFPg5nzPcXIOBSeEHXvmN8IbB2gAtsXBg/8TnBTrGycxbCGxHo540RWFAfDZ4tlkciKPX+f7
cIPwk2f1f5cxQWPU3IcUylpB3CVrHEz/lokP57UiTma5IrMjdk3fN6jGv9/FSDlQjVDx+AMJF6ZT
Vgta3JXcZm4zS9nIeTmIUu4/oZ3kC9NZndDz5nlk+nIPHUvt4xOR23Z8nRMj/ZLedf/4sfXonCiP
ws4K0juDA7+FCgtTwbd6cq/aKQ2HeLDBHRwIiVn3t10whnH+i14jNb9aRFpfurNhR4q55MkB0m8P
U23h+sY9Cnng6jifhOuA7vRqhODJh86xKxJtbPQYJOu1WS/tlGTRMGS5n2s2B3qFxhuzLBx6orwV
UnrLMeWSAK/2ZLWlAmXo2Wonda3QDSjDLYyNdeKCkQmiMAf4crev3n2iXD6AvIX55xjihPgbjwyj
4OxpBZHfaZAEPO4RqKrCIXJS9M7zGg3jAq4seqCzfPtlTirzv4IKMqncsjfi9E0gQ2UNWt7bjdTD
/UcC5eqgJEMKOGej6wzEkifd1DoNbqXjyUnNp0ESRwT+LTg8pm6NFvorarcKPBY/907O3nu6wQ0Z
K5XCh7wpCla9qW3F2NSJ1jfmY8ln98sHIPrMIlF7SxgqX1lLKsxApkMZTfADh/st3WbOxv9faY0a
d71dCnqpihQhXCtys/FNsANzXx3ZFyX9OMdEJmAUw2+lfnDH55iz5q2m4jFdkgK2JHqcviooERr3
Qv68H4yujbh0/zlNCSnPdb0TmF63ZcIRmCJFuHceA28SNO2LcjGjpNXAREGFGkLbue1NCo0/uud1
dPAL2AUsm/d/8foHqQ44BFpjik+m4riX/6fRbwRY396Jh+9Bn8Qct0l/MJSasbIOh31Yg4r3zvYS
20GcU7QAfQduMz2mQdwSoFW9jZ8S2jVtMIlFYeeW+lX/E/Yhdbqka506a4CA3MPvuVftzFSNMTr/
gzSVNam04emqFPIQM4p9F1Y4awUbibbUAPr8Ca0dVNQagDhDNp/YChKl0eF35lZqVcSILKDLAHCf
/qjG9IoCJAzYEsN9d+2lUGDz31IjZXLqhI6MvzamOmmDwdCDk1NNhkyyGhLrrFE7aw60oYQQa7Ls
bNox3Wgsp6X8hrx1afPqqQVNjjRr4bisnGo+qeGsLuB4o2T4Y+nAztZkC/8lSeRuVviUqV+EYtTS
EX0sMJKEx3gnY12jcvUmXNwM5tGBMGuqx56K9zCrFfh2Dp00pQ5LPn1VRiU6+nW8+oXiTZu894C9
rku5Tq8tQZetuHg50Kees5zMMNfS/fWYP1mPH6RW87plogNt5YWEX4P9HBHMiOmdYpjtMOEBBRJK
TAyh4r2rOGnc8/szqPRt10CdAT0fpUH/Hl4dil9foTKmLfyUt4yGniYW9SaRdXwaX9HF8upnMROQ
QM9MuupyyhkGl4wHBtKDY64PpS0P0NMO4/BCIO5/0B6FwItRgewg+3VdzuRmj67YwWCFK/ErwqWk
SEUWVRjlXxM2SEthMMNJ48VJwz7hH5US33D1XJz/N3I1BC4Dp6OcNyExYIYPwjH9KQRekZtSZjIy
TBpFCVdZ5OaxtkKWEfGRiS0BtUW97LUoNwCsydlnLyK/DAvqyXKws2Im2umEr/kB9jG2BpumGpfp
o6WJfjoMfjbkJA6XRRxRydZTef6r6P97INtrk4CvQ20I5TLtmG1gafmjgkgi2vYWhq1lFoc54RU3
G4fPeSrjoZ3OSDzmPM90e+r3MUUZ5SDs/OlLgxpPDLosd6d/edewMoeDmvrbKsyvr0jKPUWvPoAX
TIZ8j6YfCzSHUEtM7lvUTWqvzn5UlGuRJUOCj2w8jPSrAumUQyB9ONA3vCwQSkSFLRxxfrX8k6Zy
hzt3ZZzdC2dVjGJrpLYIuToSBPA1do8NXHKAuaM2c5J0iS5HHpd6XyCxdbWpFWZb5l0HLBciiP3s
VHhrVpd9GR62CNdgySTGFZDvauMRhGqy4vGXlFW9OQG7XG11wZLLgXnbbYuDNmJdkiQp5hbxg++m
tpj+NBO83SYl/IYHWUftgTF3UGNy4jBI3lgc2ZccHSxLuS2vQa+PxkW96UWux3Wd2qm8es2Oenjm
LeXo68tXXv//wBRZlw3z+yPucT9TO8smbUncmTe8s9KsLcF2HoC2K8nMBCvBbGfZGcDav+mAUjNX
42P9Nln5xivrzAibOg8xL2Nt+LZ7RNxPNt04phFLnq2Caua6bhvI8YeuuHaMrAgf8zmeNtXFgHnu
jRLa3lXDjQyIhMEW21X13iu2XlwPELSl526dw49kCUq/JX6rNTotVdO3EnfGzAyepNolC1RBolcB
1Rjb9GKLGs1lbm3OfjloV/jdq3YUxeA/LVogh4e11M+DutvborFZY2tMPkLdWme1C09kieF6Q+eZ
IClllnlvWaeWFqYQesSQOLmkVVJrhN5pQGsORO/d6fRLZ/Wi3HCO6Q26gb0annBAmUJ0GuW/gJGE
t42joeGQdgGxb5RF5tyggJpsmk6z+2Af9QGbkFrFkZD1HKkFryRXGlKx7uH/T7Gw8kQmUpBB+M1H
L6ki33qwoQ976a49vEFjzYb6p6Ho/3TTL77Dm9bMkfEbVtOvrmsM5//MZ9xe8tRoTDa9k2Fmq8VP
RFQKWJcYVMdGHDc1uyI5mSUQPS9xwVv7iESSUElPkCQS9EcyCmN5z9icVT6pKSAMhiB/wScOP+w+
MlaNToJVh890TXiFMx1VFKtDxSIW+mCOtD9rwpiP4U6dlFK4ZRjjVISj/2omWroszcEMf5c73YvK
tG/wji4onb+EGDgXYcj+OOrwf67PO1jpIJq18iqxM6Hwr9v0C+vOvoxIz23yvg1c7hYHVCGfRlBW
gDU9pZiBOsyb0YnKgP3wr59GMgwfPJNu2qlPwYeQtB4Z2zgd/Bk0G3cygp+aTLupbIZONVrud9D1
rp16qPqftpWnQ9On01QsWemQCF2FbU6ozR3rYhj9QwFHnPp6flGqHmLEUmxv2rSDHuSCHyIzMblB
+mkdIF/mxbEwFm66x15WymwoSAUuZqtSmVyATlAqvAKLRDKucnqqxpqZQ+cC+VLkVI4H7MTVw3ZW
/8l5leDATYVvmV0qEYyP1xwi2648HK2zP5e6UA/9sVUleDA/4LxQ0SWq2zwSSQ22HbJXT8L8T2b0
HShIWqlNEFSR4W2SCEpVy6C28zgQZ+brihxCnZmDIVWo7ritsirLPWR009snVM+rJr0OcjV3/Mn/
COzCmHmvqGl1+2tUIwEEvvnZj8ewQY04zIBHq9Hk4ROPvgsSS+1Mdu/WAXR6ZKT1+Zna4h6Ve2ZA
BcLY4uo2G+07LqB0rco1uBc3uBdaaqBZ1jbJ044yRlaBGgW25DtfWN1kSs28zYOuy2cZjZeL4bRE
zmU7QJvhIsw5stERiHB7Uy7Amb6t+fpvmI8EkOwqNixoomJKnlzn2DesgkBNGockTE9dfgHJUSsr
E398u0nqfmV0X3J6MxxovWCxeCb+Cl+Mqu85+7KcbB8smtEELtrKeeu5TDD716N/Bt7hD2S6W+jH
C7LCsRCoyqxOQDZHFCG8VT/IGWXqtnc7DcabN8nRQPrPG1m0tkJDpZLf/8KbhMkqjN1UFDacublr
/OOwr5tAKOAOacX1TFzDL/9aB8OKFvLUMz1RndnSwjxEAGNcymqGrc99ApM3hnw6qKyQwhy5MDTD
wBx2bskOqWnJ4MXK57sQNaOmBLiE9JYQdkIwu8jCOmgu7QMIew+KikH8Xcs+qArZ3Wa1yBns7WfR
vUvvORDgR5YG2JykGqxgnnSRyBNQrK/y5WVIIPlfjGDxUrXkSmwPKU/w5NIvtWiOkaltfJpKBi4v
+mDSvGilSzV8P25Ol0OYTwguiphT77f0pJadTs3Lw/biHlB689Cm+6yM5rQqFu8YbqbMsG6RsDnL
Ew0jV+x1xzMggBAIueGdaJRJGU5D/PEUaAJ2rnHONBnqgz/QA1RvVKVDlvgtWThUDwvBXnY3JeZM
SzooarnzahaXPdGGErdkL+dxiOCSkHlywgtBXAiCmcGgrJwLDcl1vtdnqL69wSk59mZ5rV04yzqo
IDIN/Us5AGGkekg4JNHGXJc3ZvQJrhy9ijgoSigmb1zlWLG/0ZAWpLjE+ml2NPtWDIByCyV6Jvgm
G5k7RLhMO2gEWnAGgzhsCF/2HEOK9XhKPNG42sU29zYjRnZ2yh1xVZC1t+wuJWkP0qQiGkPLNdj5
WEEZ7j5f73RFdfnrJynjQdB1PbhaeSlmrNipGa1sLIxqg4SgL5sxscisYCd1HWrdyZyeNSIkJLnF
+LSJwF3KRUPD4mZ/nUYQQCK3KN3j+6B7FKb9Bs7Yhi3o0IXnH+OJnWGE+CtU7HUZYPIYqAPXySSU
nRCOQJox08fcZLVFwWGmRb6PGQGesMB53MPLpG49iKLI0lhl8pKGdlhC5XXfdlxPDvpfb7Jw0RyA
Ia3IxiXGZOKwIPyh5vdei6guPTB0nWR83kROSNNyIBEOIgiehfCpAdPfTx5lQwzUY7DrmdOFeI47
QYTsBQMwItKJTYnCmgSTLD5QDLjNLhJdKuoNNrCdeiZLq421XGbCWEkMRZ3FxbNSUgmy9Z8gYYsg
wGlAxZreIGbjqQRIEE3GEDrpMBhXZTa7dhXxHMHAyYa7lbkMjPzaUJkZVmCMTH39r6EAbRwMYMte
VU/0P46Q2gyqi/QeQwGTA/vSr0UcrUFxaVCaiWXKQLSHIU5E8jC/AENpLQZaKjRNqIR3h254PSa1
jY06Xez5n6HrxqRs4F6S0sZZS7a11S95i95fGaFu9bzRdlMO9fZHIT7T2fzPVOzzjLhFWKTw2XD2
bbvkpL/9MgZIX/Q01I+HdelRj/t9nAPiVqOr+V2UDLRnoBLkWThipTCYbK1/GAL9gIOg1QSnnxTg
fnTGZ2Og1k4ZvAbKCusTYlzvEWUx7b4r/pusD66VIFfp0EQuGd3v0jtZSpRZPgpJfvdgUnQFJkjL
GBYDuEt7XlL4sDtgjHT86hjJ9zmmpFMvdlacX1prq2NJzb472NXClWXUJOXi5nZaJSgSVmFxRCbf
fMkf/js/B5wJi/a6iy0qbjUQX/C5VI+qydpd3YhUT/MpTeuGmenax2GF6G25Q7F+e3EARr/fadHz
LhjkwF4pJRouRSOsH0/udt3XyTVolMQ/RhWgyZW/kWCu4WML/mrK+JxGYGQ2NDyhyhZX5lu9WJJD
O/Yo4JxHf1XTNwJBUgGUpYK/9b/FJymqRQ1Fjjl1K2NzmdgjJtwurELIPhOaR8szIyvK6vlRLk5d
VSi6HC11UV4en0wtGBbwlzg70lgn/ZJdCN7s3ae8yLC68FZpYD7254XcQCeg32pSdDs0MFVsLmVx
XAafwUKDnr6SAW4Ldudjb96kMh7tT38aWO1Sr5J5IRulVZGhFHUa3fsgesquG+TQtaDZrxhTSPtE
jbAGtxBqNPp3wBG3BDsMqX2s/trkeszvt7305HnTWCYdCfKH3iZYTMN0JpdpdtzHWL+W3t1CUAu6
9PSvNi4T+L/50vFUweBEA4bIBb46Lp6nMJMt+GQksqcraLeW75LBTUyqj2LAdEVEWRUMSRf3kcYI
eheJiNhHoSnW5NtRArqtc1RbjMBmf1VuvvZL0NHf+orIMjjpU3SJt3YF2Mm2EWotNeNZZR4263dF
gSVJtd+AIldkopJ0EJJJZ02kRwGuaGk+BB3l+Ep9qO9rb0pMzBRklBQMORTYuprTb/KHTGps1ZoB
1TwWaAtmWa6qWOVWFWmerUtVP5nqv56ulIwJFTdoN/wSpo7w8V47owT3SrJETwdYgppel0SrW1Xo
CaZzoU7rt2fzLi50rC4d2i3onHGzg0akm0VvpNa7ZGobulJz8pOL/vpbChXQjk2vx2ZQ5Hc9eg5h
tuJ1IcHaiuHD5F4MVI5gWAs+CVWdbPloh1KOTVQuHZxS+JI20NuymOu3l13tC58Ptn6GyFgyxk5w
0m95ui8jrUC9kRSrAWVDA9eDI0OqVZMAqPjZMCRAUrqFokj8PyxH5QE2EXmdZHyPPzsye3yFt3YO
yUpC0gRuED+cWZybMt+Kxrmjf78dCt6kG1ECQW3WHsRu6WqkyBPJOSCPrDKMjhKiM955i1uR3VBw
W6p7bALn5Ifhb3tcI0L8LY6CyvCvuCHWO3fQZnD+vFiYk52/pRpVbuJBDxk0aAqv81d6Tl9IPRAD
88aSU99l7MJ9U2zDxKXh9yQoAJil681uGHEHgtfbhEKdPWPH3jiYhpotwPCHfOKbYCDCxqCwqRfN
6rSFmNx2zC/yyA6jv4OIuKxlrkFpps0uy19/Z+ZfvWQsLlVbL1WG7MccumYec13BNJ6LoP8s4lVm
BnRMzDABoBD78UpbACwcRFU3CYDAXWCNdxRTAo0OxmrVh2iUxAo6y3stQjh0tw3x42wYk1pmFRUe
iTNlWJZuokbm7+VtT9J713rc7FEZaMXxxNxzh8mGTmOXkKLTGP3vUyralRdAh9Nc7vWRLGqj9BXs
RFFf+rpyzeNDenwDdWnFrR0eSY+jh1SB9w2FU/f9dT7hb6NWSB1Nm28ntfuFUTr4bwUKjgpCjAuQ
mJ7UoflE2iqCsLjaDVsTtKlrsRDZ6X1ZDZtKlgX6x6HyttdLkQW4YFYlgFord3+92ZxL7PP25dnn
gGELP+ZhNvDXWYIUL015gyr9paywwwxxTZ0Cw+cjFo3REwNF9l1+y0VOZp5usbDAh/UzI8P5jVFD
j8jLaeyUhYXbwe6CZ1ei5LG6O0wLf3eTDTf+uTQOIr+pNyuLbI4E1dQCg7WHZFypNb1NPk+gI3dm
XSaAZyzBNW+fA9bejEO4tRguvVDKTcwlFir7P2WzD8K7zJ7mqY/4vO0FVWfnmiogbDdfKQhyM2+b
OfePxsXcoR9h/uE7RPPc6u2vSDNY5/BPJZu48E95f/NA3sN8vuLAEqH4LMakxcY3meSIIdaWVKoD
njgrLy6ULNMG/zOHnt4wyLpV+c/Hp3/C04fmhL32jt4X5BTfnjIDJHIs/gK5mB+wP/EO8Dma5UUA
OMvM2MXaJp0jDMKQj4vIUdO8xOmg7tfQsy0e/TjUijHWCpy6yXVma2E2FEQE/sZIVu7j+z+W7+kp
Wqex3BvW3bSsKh/8WIG9cmoyfM1sYaQjn2m4V3ZGk1he2wz39ghLvqowPha3lf2rmpgym62SLxVF
DlDzz5ItKczs9HwXCf8PQqgz8njLZBRblNLaVqkxcbquaAANhCtJHFvgGVT8K8X0v+3K1s8Tqcvs
CON8xYOt0TWhJPDEMKlu5tJN5Qan9z6i73T+iO3lhmOPNvf3oJzx15ogai9P5ht2bg6HVpORf/w3
haKGZ6YxY9ljQxy62+/7CHiAk1wuhPaynth5La7lK284+MJ4EpxQDElevWRAZfxlZg8siimA4n2l
5i8/nr6xIne4IXEdT/4pbJnzo6gt+11rq5iVHPET3lvvrmky/VBZtbRKH2Qrrw3EDacykzKMgSvA
AHi3zw7ns+j+Om/+wZnC3b9PcQfEjC5vXoktTSdN3Qniy3NCeGW8F+ECdP/puZzgDsAD/YXkRQqi
HrPBpWvL/bWFY5kRxWiwZYm4BprLx2H0IfSOyO77/MTd9pfDNK5+Ba7qqzooiTRK++FrdBMNRWmk
gjxZ/cVKA2DosvfPFSUhlWs5TnYkU4SEXVdyOjGdfezK1Ja0qeNU9W2VNUlhkvQ4rb/FJEwfjnEp
f3+fkQHub7r1eOzMLbEyHkffcfhSz5foqWwFt4zl1uzkiPI4ONMTB7Sn1gBaIefXR9MaqkN3t7dJ
JVj5emjmLzv7zMZXaxJycXKK9Fuqb8YRPDtEH3tk95xY1gx/krlpMjgVA30zckXcF1XC7YNctzpU
0KQ3yPVFi19wHAFerRAi37Lvl37UF30TRI7ZLnrPSiG73v/89o3D5zWkHx1PjA2ZXnASWh9nywfX
t/QkVZj1MESTBCj6IM1Um2eJ12zFLGCSsAL+ZNVDHpnsocZyuWKfUKJBs6maLM964kMcrVhdzz1+
amBoBsptMvdf6/rCuL3Ax0Fw4Ah3TL1lBLxDQ5RgVaUiQbPEqIWg9AZvqNCoL0tWXKwBJJD1VrOc
Ky9pdrBct5KdlZ/QvgjEjKypj1t6GjJC4WHUVqJPngjV3ut2ggcJ5iDDo4/zL+xpTEmyUVUln+Pb
RuLq4GCg8wDN0ViVf3qBX0M0TOqCSIL9isfCvR57G0IKkrghNCGFaPuamoe4RTpbmY692mplcuN+
wRoOXMTN3R0u4bRNclVoT8lOA3H0bxyk3/uUSNSAiBnMQ/hmYCok7aeaHTSjKBiwjMoxlpLB1Exn
hy4fiLpOpG+GX6mPoo4WRktHw40MD26N17ykBdi3wv5to3OzN4OimnN7Np/odt88twXB4Woy49Ju
LKagaR54ASM6Bilm133hE8eFvrwEKx/xzgD0nWPxOCuVK+fsXN89f/dEzAXE+Yz+9YyALyQucmPs
dMOJwLon/hwqGkna1NGa6gAD1Hdv+uVl7mHTcbYQkstXR7k89mxz1GFL77caH/stdMCO8ZAdl5xW
qSCIffj1UV7o8kZ+L59HeOS3zuE0S8EUTYgMrn2t2HzS4muaYUWMvYbksUOjWmvIHqAX2XHlSc8v
JHIgJ89weeANAblvAfR/GKk4lIKWz6KTl3PKAPqEhhvn43ocyo9KtJSy/8tuSidFRzuWdexok+D3
R+m22SWB8bV4s+R41MwF6KeF6PTiKv3MWqCKRHHLzz3DaFEzU+DndCBWcrSLL0YWl8OD9wGlumhS
iYR3woYTg2D9owGS4v7wTRUhZ5qcaWCkBsVMDw/WosgmhltudmJ43xC6te5RxQciacxGIgkPFz0q
GWXGnHhdk/kNpMj5kW2RPeCGR8UCwCS+Z/DfhJ9JRuA5Rq1n4d3NBC968WCxm1jqlUuupWaweD7F
lqREWSf/g6XXIdSlS17y9vCbfFctS7pl6q8iZdY5lyxxiLYMB+vcTArnfxU+oyMHINq54cEw6etm
reDB1sx9WAyDZbOxwl9NCWP9F3DcyLDFuQUc0qvRP4x4Hw7oexfAwAWWJbyPwihs73gmM95HQeMK
7TH8peOwl3+sbn2acJK0u1UuTHwWlnW1P16Nq7Ml0k9pz2H5pCPrn/W5XE6vOBeAi4vTBjQss29j
TQv3fMNWx0bf05w00ZBTIQy2ca1fEb4oP3nBd8WquDoc/FeJrSpSep3NX2ZeBTcli8ar/G+tmK5A
O9mgnUgfRTJqZ75JrEtBrk9F+EYm7g+Mu9XQWNbtixtePdmMiGzgX/u6oeW0is3L2SAEG1GqygNq
ayIm17IXGq8vzgQraYP4dPhGLcnekisuRDFOjDS+lPEZifhb5Noev/0KE9+gExSWFruWm5MaCO9X
sAI/9CvtDJ52lEIrZQOns0oYi9xE6O6OcrWzUov+ONcN+Fe440aveb3GJLk7ZjJU7xCR/IkQkJX6
NNNgd6C3c99PZrLf1zlHw931dhHgRI/R1pyGlwbxyN0kIcOWD9TFv5Dug1svRyOzjuaW2sWbvsxR
IPkXRnGJ6f5T8d4y1nfOc+5LxZfCB0uz49trECKhi8isZ9o9i6lOewMUpCFg0m4hebp8s9SGwn9g
/sXXcBRs0mgFmMdAe5CmbfjjFOx+gnqT/olyeYv6AmSSu/cmiPdz/A7UZIl0MbgrZi35WCV1QN8R
InbuigH3GoDhfhrif4hH2cYRw52NDWL6ww9q5cu7EOy2ig7V/OF+L0BkNxjOVb+E2nx69I5Cl+Ez
re2osMLyzUwyBK2SmKU8DaD0mqLsX/dJYpOpEocxaPD77xFq3ZbTTSdjgiSJCXncVwNcxrdHTK/H
teEZaeKsXrIR2sscVm5xZFBeFLBGHUJdiuYiHMukh9fG/O6hxyQY95UQU0hEjY0sskmnpJCrkjO4
5COike9NWgie08rUvg8k22ILgmXKx21T+XNzUnmfhocPida+l/pI/IADicmDjSYPCLUT3RLtVC49
/GQB+niGu02h9vItqGELXV3J6krEibXnUsuA5KAOWKg/qI8vmB0wIrOa5mb0cocq3BYHUHh12GEe
s370MEY8RkuPFinqyDZIPlzopD3TwuAwQHwT6myHFd0f5SR90r5ahSjp02jsrV9qKDq/GvCvcxEP
LkdH8la7Ez2FJaX7NUwpZJfgjJtme8aT4kHDVEJXwz3TdVsczxyAnp/VDaDWQaMNitsUPkctf2gg
iqG4gMotoGKuAH0wRMD7d2DE9zna7NGqtXJFdof7eBnWp+LvFaKFAYq/oG8TPqXy60AEH0EJCwDr
z/OXaOw107ZQQHoXd3TMEUjHMOKXVSIIAFYBlxUxc14wq3cwEqlGwqJ7NJ7iH5J2x4k0fns6qrAH
c9WttaTa8prff7d6ywvuDzu/HLVDoueMqx+Qd3MV3U0JT4U/s/H6jFD3qg3PzoBzYpeUCmztwKsr
OnbM9VR6Ub+rYxW9hOAO9eGzJQKmtHHkLyaKqVq/KkLCScmHysYHEspiVGjMrNSBJDxt+KAolaMO
ZDEOzSRV8B9/tH76ShWCkMcoMQeybjb11FxruntFBDdFPlRN6SuNaS9vP5zYySiqH6Zoy7M3Pua8
jCxhmE5gcZkUW0bZtKmvghr9z4inNa/PJdLwoshXsQZQMIuztO0fv6jX5mfb/eObAM2ktA4PwX2x
xd/70th6tl8QvNAAFAWvJG0B1usgC0/FIZ/kaPs9/7gVHQoV6aM1oKkJsLhJ68LjskMNYuobNL0s
P4878SRCJ1tERTdT9dib0OUq6+ljykmYbFEX/iOP+EGd/bgTkWbDCn+suWLxBY3Zn4bDCMoq72TS
jsH/6Bl0Z+W4ALWUSfibpMeAZFi7ur1q6nt+P2e8vWdSYFhzzWCyPQKoS4iYzjfvNz0kE78r/c3x
aTHXcj0MnxnWRUzwShC2fTw0eyvY/F1LZvatoWadXXBWYe2JUcd9znVuLlf4yGi/GzTYe2A6dL8p
mj+QUdR+jKj4F+BXW6y0tdv3Y2am0LI90aSG/dQ5jBi5slN/oFnbkmFdAqHdpzGXwbF8Xp5+1Ujl
QGBeXXvgRx7e0Z1fn5FMAi+if5BS2XCLcLXdXRrQV7GMP+LOA2s4oe/m7m07JsvLtjuJA8nqJLVJ
Ebf8KWc4smD6zOqVOCvrz/KL0DNsA+knp4hVX97DT0LejDfBtkjwF26+hH26V8+8h2QiBIudqT/l
dgcJKp8u5LUXtedyKH0SBVIolLG/y/gRk17J+vzv698gMnrzxaaHIRGEA1mIVQkKMAvsUO2T1Uab
CvWmYHilDeccCjTPlScypkgo6uwgP55mzCcREDVe/psBmLvmp+NS04XIqaUeX91Pz3GDccs9SlWs
gJ4vxPZ6hYU0FtIwmqmo+dW4rPGJXtTn0k4bzZ5P9r3ViYtUxhyOub+L9UYGoUF3fC+PJ8Jk9t7x
g0pBcOwnsHhalCVnNZftzugdLhVV9B/EN1SxFllxfpq8z01Imt0o4ps60l3iPu0YpNSjzZ/mVb0k
N8vdQtTnsBEaN1HvJScAZjeHjjrKLG53OMuEl1cjVlmY5OFW9H5VnfQvv8dPmU63VZvn06H5JUR1
6+kwSqAf0QAaEgosrGMS9DZVVvvt5FUVldGTjb39xE/gTqpSAQy6kQQsy1ZhAPCdoCBXCrjPKMrX
ibZJIH2MkqxXAzw7OQQ20tyT653Ot+FDawQv1W/QY0t4JnvdQVvLk+d7dpZBXtyCX1DPtnrEhdIx
H7ouXtEGchSy5d/gLYh0vjaSTDm9zFpe41uZzIldU8UMjJcObxrP9UEE3+p4LzkF84/yEjzrIi5y
PDLbvAfvIdwkLhB3+u3LMJjRV68i5jbnwydetfBaTsRtP1jJSAlfB7hxSFFhkDQ/SkhX+D+Aws8R
sDYpawdEalkiAqkLtPGwvV22JDCKLu1ljP7zHlPj/eBhj3/hItlSDaYf5xHW4BmTDnQqvXZfwwcP
0pkVckVXqkCO9Pr1JIGowuWE6jXNPQ0nw5hyzCOfZovaisofBMdgSRAX8aIzv3JMyvOdnzliFpZ4
a+KPLxHSUO/zAt1zStCpmVrb5yho1sizbFEHx4VGRTYjA32HDzTSjb20ZiNigQZ+5dikILIeU3sc
h8bujz47gEd/QiubcxNVCydJIRkLivpbmB7AV+AuwkwJJHwTuhGS8pQrprK5+zUsbBhoAhw6ICZ0
hHv+nb6qT0Xs3eKaKppAydPZyztp9ejQWwE+m+r3rKAl3iqABNlFKNbHLS0bvOJE8DSK3iXjAQUb
JYuf5HZq2IdznbrK8Yi6aBUKBQQRAF9uUl140JiqGsquXhp0EdBrf3CAh3O76x2h6K/P61IPG/J1
ausiNGRTNDOA0YkGq53pOD3wpVJZoTKOs+IL4MkDml9LJaf4XHkh5vfaX2ZQaRFz7EP7Xpe8QHJB
1ttCMxwn4AZ+j+0jLkFsevoZuWShicni19z+jB9rvQB6lpyvbcD5SiNypjy8K3Ihdh4UdXB4QkrG
s/QztfWFaWFNLpdUVL+xr2JeF5Wy8ZV7vyt9r07O/lIj4E95iLcfoO6MLBHnPqJAtBwesUdSh0J1
xDuLu4Phr4PW37lMmt+z24kAt+VPp0ZZwTdyn0mvUyZWWwrylXYeqaDz3DZCNZXu1DMOU5PTi171
Zhdd9vOm0r7j128ka+Xi0gDqhdwWlgEnl9ozbu/KHZDKKHu8WJmyf8sZ+sM2ZGwoR22yLxrOChRu
RtVTnDshkg90+U3XrNxElRTsyHimvZrAPU5G/KyFjCWTrR+hSbnfZcvhCmtscpeNV+R6IDQ1/n2l
y29i8UORjcSdVq1pZotGP8w3fqEhVQLIk4g1pktm71Q4MRL0uNOViit2zlkWTp7M6Hy98cVe3PqG
oqUwFgnJjP/LkFqUvGM/HD87maIpTkW3jQZZzgoeMa/IkGL+YN8mxV+Y0XTkZJJ1Xr5l02LXwpt5
Ga9JjuE7OhPRqbqmS2JP3wB3y5t8qeocC4XMIPlZ8ISeejYy77HGakJMUG7YZpAXW9aWcdaK5msA
zU5I2ieBndn6vJD12opqA1JCp4wy2G8O/3uBDvMPrUAOkMCNjiMf2XCDu/zY/3pDVHc4gLarGP78
NHwIlf14Eh4DQkc0s14hs9vW04ZdMgxybE2QukttkO3atZHcc2EDgv14B+LCdwbq3OS/wEuOzx/b
9RN2or13K8a3LrqJoWtzmv6l95Ev/2ODop7eSuVIrycTZjA4mvZBbTrbubJ1HFT3bLEK0bXt0drb
TXW5Ytw9vw81m/RNcYr4MCiYWSIUwa3IxEMlBBtVPlKVfd3+QBxdmlS4rbzxMZzaEZTXhYnrcr74
8aFx3pvkdfomKEO9KaAzvlxGyNdtxypOUvWZJXhUwGCCUjw53Za2HsfIyBL6v4eVp5PDQZe78daZ
a5VPpXVS7JZP/FwXt2BR9wVuDofA/XnCmWAUA8Noo0jYAqhjC9Jdijmm2ycsFsOp8UpJEsn9ZnFs
QcXInhfYfTsnWRzN3wMepWTpG57cCDiB1aEGrc/ik08vMhywgRyeBWxnXVBQipUh4CEWHNeXpWHZ
X19YTPf1rsmRTgAaxii0ZOQiTswQCVKrYujS8IDPOSuWA9B7EGZBLAdogc/0FjCHiK5b3NexE16O
e2UWZSjR3Ut4ZZ4+cTnTBFATLIBY0mtxyWDzovlSIU1B5XnUYatOkGJ6AYGRsLVDZGloIo1SnKSg
ELKHj2vWZfsFrfUEA/mRn4sjCUtKgO7peAYoW9mVCzU42PD3Rny6MM7Ec91FOPllkDxFLZsqqBWu
2+WJ48yvWqyBEqryihtJDhqebgw60pciOZWCWlzDo8IgEOPw9kgWQsm+v7m+Ju70U0gK6PalwVvp
al7jk5+esVXOqQrXESCXmC7DXaR8nmacnOMBHTJOAIuWuDej26TUUt4VobsrRyeIwKqGOP//Q2PW
ZmQjSc48FOzd36cKQFBkPxSEp9Ei/liuGgbFWVsS1WIJ9CFn33ZfXZRiR9ej4ftQHpVxVP192TI6
RARNxF4uNWo65Wq6PjINE4Jf1Kd5RXoh6RpHKyN8eXchw+TkLr44yv9/nZT9y1uay+Hme0SojN7Z
bxfVyEXfIRYrDEMJA3S36/xCR9jKX99N6BgWBNQ9r7ngf4RnxZ1Mkq9orqEj6YuOP/5WOZFNXCH1
0bw7+2qJVzCXgESAMZzMaAshdUuB2Yf4fLn3YWy08TCQgCRSjfUD5qASE+OPCogRx/5cs0cODMLP
SZFVH17CZ/kkNtZ0mgI8Qw609xqfSRI5mAJvY8f4yVsMVhqywM+ezpHayO0pa5GKqQHe5NyS/949
/+jKGlA3YwlZEd6Rdj2AeO/1cWb9ycrY4uU5T77ZRcXguArE8MIIL//Ak+HH6icFfMW7iL9k7xRv
ebXjjGAr/rkO5iRm7Nwvf3NZF3uDzk2QKvdK2xqnaF1Si+zFLjhpc+HqsVyBjgCSblS+IaWcLtb/
rUAWKJ7k5iM+PNbfyazvvh7hqFbZe28lZ0ta9+VnKiaYW3wCdaDuv+/G5cFA3P301cjZO4yOwDRm
iz+F0F9K1SLa8mnt0I656OTfGEo0h/dXBx/izMRVmiJ9KJvE4xNKChyToPw7XslUni6fxrste/iW
weW4n/TBVmVImYaJ7j9wen3auFQmOUtSVZQ9Vn9eGcxJKLqS3bPYpiiJLc0x9QDGaWxm5M9vZKFi
oiXrDjMv8J725KBlR1G7uJ7MC8vo/hhouyUGx6FIG6KfGi993sbTyzjTgrF+bGrIk+mflVGrsWrp
NUEDVRvuhUHwMrnXUS9TiHfTF8uRsUqxvgqXisLo+BjUV1RgaCwqIxaHn9QFz8iwqRD8rc7RbMWh
DUHbF85HA9ky0BPU1BINgUguE/tEX1HlvfC4HJkB0DseXHzRMm/LknQfOpB/C9/ym/93JzZdvQaL
O99H+Rn7jF4LpEY+UufL1SjKdGQSCUwR2GhDgDvGgozewtoesPxNJtnca6VMB0mZ6M5yx6/uRWXB
IE9Lwa7UjFk/WFPvXlJHq2xHSqyRxFUKHj7l9zTF+K6TaU3NDvLYfFS7lR28xOS+dF07eo5lQ3HY
Rj+jmxcLXjROq8KgtMVQQxo4cuiJZ0Tdwse99BnPqgsUYpQSKejI7OWF/3Vew2/XA1LZkJS6qlKR
QCdaNmP2oO8y7Echzod4RaR71C3LcCg3TanABMWzDKanbVkRxd49F6hEOKA1umNH2hJ7dHWCbZnr
JVcRdeRuWkFhAXp/Q3h9wt6UQzG3mONoTvqouavW40tvjwXHzQO+jeVugBUouUXCtbYD4MjOMG5v
U772hSodGgUsbVDf62Lw2wKC76/cjHReEE8mZA5HV09THHKLynmIB9kHQBWlHcpKer+EdJWoaWru
V3P2c6URY0Pw11YvzzdZfz8DmjXmVzlGwomajUwN0rUhsTTCdI78HwOJ5sVXMioPogT2cYXezWMY
hvVB8SHhyd3QVP4DOWc8wi+n1aKXcaY1QhF5/8Lfsq4Mi044bczzCLXvOHACGNnavvPN0KbfeqQF
Tr9xSWq7sIGcRHbLvMIJfymFfJxBGwAsImmtyfsxv2l+a5TTYSgLsHWDOcDWCz8Ug8iavC7sdVf5
zfyF2/YtdfQ9+GqiH2CP8Zl5ihwHsvis8ZDJWFgffsdFGzkwYaAO3JAtpfg49KfvUZ9d70hIh89y
8tIlQs7M7toFMX66rp2mhM2SaZ0QZDoj7ePYmg2gs44XY7BJ+9la+ZG4B0W9sZtT+fxQvkX2EBVn
bAoVJ+s2HDzFB56/CgRKR8SFF9yA0NIqGVuLmE3EJiarUxf3J6HVG7t8QN7zZiT8EPhCa+c8zSHn
LjC9yEFRSX8EjAiG3TJnOdkjQzuclLTg0i/OkeVrmBMjWXyLqsMZRDOf1S/sMX7UMy6b34RFJ98y
tkCUsf4KpahERLiKhjvhnSH+gNU6laM0hNubIYWo8Ex8VUJe0OOH21OrQDb+0AdZVKvU/EyNNW1i
ozqhAqa8cAdC4DVHhyPp0Pe3JzG0KYRx1Eo+gRxkGiYP3ItV0qTjLssc8vY1Ws1CFfk5sUMhD7aD
0KvRTMhmEatBAZnFLEDKsvGLgV+KSrxk9LfWV17Au8tD3453pNH2EHaH6J3bHah7FXGRJVABH0Yq
epM/KRy5d0kC6JmLnZ/N6KyylEpZ1F/Ziza86tXyKh41sqwJTc6b4tcNK92haCeaRxwIxCGVQhtO
ZuUcgEg/uxYpAEPRnGwnjbToxCUMIlsGguSNdXPqfCCBjh7uOOmA0em03ZMMGkztr6sqmzswGPHe
QSavf8DNRb58HCN5kMqdJcbWyWD4mD7dSLhSN3n7UQ7CZp+rkwSrA6Rk4bAoiJqG+CMNjTZUxR4Q
aC3mk4xbS1ZnPfo9EisEO4kL7Q6xmDfw8q6Xz9vQmVVifPNBzBBpD00wi6Ttybsgu2TSkYVQIZR4
ve2F8nzdcgaOS/8hKcaR/PE/eODeTKuHbGpDlk7tWQcgzKNVfKoU3VwSZ8AMcQsEKhrvcioCreZc
On1eyvTWXjkbb+0gQjHX/hpu04xxCJ6xjajP5UDq+nVOKT5/ex52o/wyVtXq/ykqzL5k6tetkTh8
W13TSqd3toaDdX1bt4xlu5vwyG5l5FTMVnPPHszKYPe5qjlpVaAoK4mUJOXsEnrsUN1MgcJkYnwf
jQG8mj9CltlnXo2kI4dBxb0z056jOP9FXdSjWtHkLUd2bHAQpPkunQlCOks87BLK2RUVd2uxjFM1
LSAbSeZU0+qh1ZRgv93NeWQytw6euAyd83pae99g+Wh1cx/agaVm6WGhNVfd4212l1GEaO7BLIbO
DerIqv5PGmltLuNoe6L3e8Pkxb6VxjHusFN13PSMjLENyeoBOFsaT29ADx6t5ZwV6jUtsJJMgbvp
apGDFNLgKHZZZ1mHQ+Boc+9WoFas6jd5xiL+HYeTSzcQE4FHL77lBdMKrzhNPgX+lDg3NLuSNijO
VNBWqb0r8yEkfdlLbBue51a25aE6+w4SH3pdRoA4hbicDMnqJ0yq+Tn6sC3IEmTZxlCLM6f1hY9R
YyqaJpMVzuM/EHczB5KGjCmKcRmCYW/4PpuQ+2qs2FCuNlYSXrsPx45m8DMrqFpkDYWPmk7C8ZXZ
3v9+yrR7AtWa1wdsnWm5n6x71niAo4MyVbFGmENbJxGvCc1t0MOQTz8W6+zEVepxgP0H7kcZ6oQ2
AZPsc96dmlxP6+H9wDqDpjzAqx5uviOfNM2W4tY1aIIYmlFy95X/f/1UggRlr/WN6nS34a+ixVkp
iPzaeoNfoBdx9a/wokm82U4o+3wfE2enRqEjd5kzG1Z0lQW6TuNsVwB87W0XzvxsVomjFBCDI/8B
/CsbR56xHyWNa94dJJmjH4BfKKE3j45kthy5NrbUNxv78NYm27OE463MkzSnOGG6a6vGuOi9hTOf
swjdxtnnTWK8FL8jSpYW2SzfjWMQb/bGoFn38llZfHbkMIzXqEYIn07/0sZJd5ZB3jdXEOHwq2mh
0OsygTGlH6lzNOT+SBUQVF1JBphO49HJVeGCK9nzBu9bVkUhRUtASppFw+xU+3Ihb/t713GcH5vq
WT5jlKwOUIKDttbNK9NUgaWjGk8U7KCaeERm/dlaQyM7t9ACrQtIw51fuV9c2Y4HBsiY0lh30ixU
PQ1U2J/simxyGNw5ANYPPgDVNgyjBU1yQmvIUlHA2YNk7hF6uv/B1WEy7WuIKaGY+FWKBlPx3UXa
1Ea/4AxjDzcvyMjR3EHFFkRza29QxPFmGWMXWDkKDcP603okF3REwBsq3HN106fKoMp76p9t3KtF
WT//nSiH5+SPttl++6Y6beQazMuQ1H/UbhfBBjDZ770pcStJTVgbws7dcNBpbcv2TmyVyKKDhgTm
hl9+x32+m66JeF4xRHUbiAeHDkD6kduo35z6GMQKzjiqgsz/ofySDFRf6QfmOJHIosEMQCyN0oEM
4AsEyHURb0OHS9Xi7D/0FiiFU67ItPoutdL2gJWnJF7Sz77CgBtxxWp3EmSOCj2jENTTtP8X1Fut
cXKgM3TEx5qalCOcOXUifIyRHH5e4z7NEJUpwaitEJ8FtcRYqOLA1C2NeFMBYkSZ0ZVCXg67ab0e
YwclNfIkau6+9gwjJimHGQ9KuJesqvsEzwmxzq6esDvNYafurBYNOUtgQO0TLlS3NN9THwW3TyT/
dJ58JdoGtmhAooW1wE5+LbTPKW86xdoAv8PR+MBl11hGWdawzdO4rmTK4WD0uLsE7lx/Htw/meMq
Zj7LXSLyGJvaw5Zy6KDyujpYwYdC7jibkJ6qzz9hpqxl6ya41Ms/DqCid6cbzPUIeTc/MB6F3/e9
3UtZ1VAmwNE9IFHa8HiTUbaLIET+AWTb+hxPkg1ynOa+z89wtFrLKroa8tcLNOS1c+rdcoH2WRUY
xHoHmQKY4wUAz/zmRbL0rA47ZSRf3vSujAU58FtaEzQVd8FY8cILu3pZnrYg1sr2IsYPkcfmq8K4
rwmmJ0FEh5yEdo1/CMR4pwBhQcAcM0r7vQle8HRZHqcv72yUKP6gXfVAlM2XFLw8GF7L+O+HBPKI
P49lnml3M5XglKjIkI35NGS5r2f+TkuLJJ+4TwRqJRWbs4mlYgw4kBTdM7lUdXo8v32ziFzMaByj
Od3MEzXJbGh7p4Br2xSumYujxe3wj1b0aDFWyIg1hWGgXVGhbfsn2upC6hZgRQBfBGOitNB0Pua8
hZNTYsFHK9rxpsUM9pZYL/QTH6s/ONfZSSZ21Bvm+GNUKvwWXdvWmQ3CyqCsNG90cn54cgZGAUFI
u1WnGLNwESkUVizO/6XfsBNk1MvCQXtmYb4n7H0j23oZDMt6lSNDUZdtw6iagiCn1TgFJmrnV/Pe
FPFCyCa327WsdNwl51K6P98qXNfKtFuwIglVpCW5GrewZQagLxNZ6xLFnAw5+mwr/cDwpHu7dXv2
YlYzHRT4S7SnZvdanc/8SFi0yOCA6qWDPIXTAFloKVjhyY2nNOiIuJThBP7yclUhqIpZl2O2dS0d
D3m9j2sMcviINEFYqYGtyfQZgW5sFSDSI/DzMly1C111lAvh6QvNFTWWjK2yQiuDTQXY/s2QNWe1
9K+scWJKjy8RAyZeNR7YklcMHIFT7RHi1ZxD8o6OfZ/GwWm2GYIqfqxx451Sy2gFWHgHmjkXMEen
EIZbUEMFU9XA04uYVXs4MQV5itetcpHZbEXrVybq+3wqThqVMmy3by4jeuR8uaP9Oqrc+pYP05Ij
ADtBQ8xBhBLA4j3FSYybeRzvSN4Pxj8ViURXraqajfwJvP4sGEChkkJnTiu+Jv5OGU59DWh30180
kH6KZ2vRY/TvGeS+S5QSIY9hCgsK0/cmzBzYgxRyCLLg6uXYTkQyoqL7JhdSSL5L0CvqtBU3V+Lz
FqlXt773fbdWo3JOccKmt4AszQWFVZC6jzCJ8fdUtE0NIzFfQl3KTyg1i+7+8pTN1hZE3X3fgS+2
aJoMLSrnjc4NXpuZXe2+Nv8Y4FdKly+W9nbGFt+FouxVDrZV2MEkzqWe6fhvX9UbEmc45RdB+ykA
9+HR4w+diPeTCX+Fgkv46zxnM31uyXNhZ3crEImrAzYGuSnB1R9JSYFL+AHG//fy1D5mBQ5v2TO9
2uA1Mn1heGmGuG2JNZwdxYuR9tHzM7ugovbqAcGmxVtQdBnpgTHfyl70LwN1QZDxcQ0vlsZJRVoo
7ZoZRTal7keKx4uVSn4DeF7S5NU91A6VwFyABDq68f1roDCSMu2pdnVLeAXecPXaW5V5bdFYQ9bV
W7eku/D7cOIUjYV17a6x1s5i++ER1ChSMdq/jtioxjHw5oCtJt0ooQGZHN1OMSlg9k5x12iBZWNp
GqolX39ZYQ8eChKEsznOIrt6mJcTREXmEYkTEFhUFq0eKzlNfErTav6W0frfQ3BHxS/szetoxP1g
FLVrvJVzUfWqZSGClsb7z4tXayTmbpy/2hNa0hP3pqDbswfvq5s0nTYTfHMZeuqQ2qOLJuW1DKFK
ETCqPsTBJC6IySP50ExwT4lAJquz9WlQtK6yzRKqePpNoMhBBdbEKf5bmROb8C83V637VcEjQ2vY
z4BfMBHkjtia3TesTyZQwccFi0ik1pnndmd0JSQ/yczPD7M+OSsPFKuMgyWVyTMmpleLhLMtJAV/
1NY4GEcsrDGZktAY29MbqMcfg9QBMvMa0eqht+YKzSrv4DWLcMgV9gXdXN9j29+dOAgwSQn4TNix
6CnznNRXP8c7/0V7VitkWXMjKAKZdQbunSwt9ex3oT0NVE9Ton1KVe5Gcbca3DjOwhOqYnShaCNS
O3uX746IE8cbzUtQcWkIFBXzsHwj6BZeWlIuSS2QcRAZmBOYcY2QNDUg3i2tT1BCWwwx+1mlOiyk
w858FRMFXcnyRzwx4v+YHVdFZVyxneRdVawGBXAFPHUlARu+TvqWd7LSVyYTBEmVdxfnC8J08+u8
PxqoszxAOJ2k9m1aTmP/HeZQYSNcKNKbm3/gwiqG/PG7A5WSV5TifO5H5YIUJyBeyAz9Dc7iK1qf
sqQb+1p0NLnh+ctSJDph1/ST4FRSb/iwjVvnm2kVELpe8AZi5DmejlzGHKAkN0604a2qHq/lPa6Z
XNHNNf9LWddO06ZRbua3LfC/BjsYw05o+Q3a9oFpjB88IH3/nIjkPmhHn5hxHdypmuWjh6AN58X8
ScKc+gZWhJeYkaKcfGW6xgAxCYOiyQwNqkffzeYdkJfFPOH+hg1plNqik05Jxyb5SNuez8TgfVv1
334lcDzhNFl28tszUQUg11Ifg76oK4pygh88xZvbbJqVTK+lM3fVxNDYvDuP8rXSNpdizSgDXX7I
vNCVxSRYl58tCWiKpZpqEqk/LUNHyjCgBj4JYEcODdRHZqtp4EzPPW5fSpmW6AXEb9Q7mbClCShE
4Br6p5R403irwcaWnOunHOCYPYj19hkAGU+zXpyIBCCbGKoRaki1dKfDKqzJpbmnm/9W4kMqlwKx
ef6nKmUMsuy942HxIHKh4LjsLYnuC/oHDb+idB4xR6SLJTiuppYX6qv00t1fMkQcgKuJYK1nThRv
2Lvn/ZMexcNicfNPDKwiaHRHAvasJcLb1XzKslEd3nVGgvnF42EiMQsmwm0ICKC/t/8HNoPxo7VY
aqzM0fqcZUnDun6n/bkCWe5iHwLEPFwkhHfro33COuSDybuiS7H8H5jb5Pzjvs/kDPDjlDMmJcb7
8c1ScKO1Cv1Jlv10yVXzh9Khi5VFwJF5xQL9yWjdNBozrbq4EOIBDdauVgS+gKz12sbH0nJDzjbN
cbmXNu2l2TWafEBXsrUnMuVNcLM0m7FkN9nvPGC1vfbsekHzsVAQM1IFQk+FEWT/oNGMLGqFQ15Z
Up/SHFsE0QAk9zyODaF76JLWKHFwpGNHJZwy4CMixqk/edz8x2ioicGJLderbc6kXDrfBvFMac6X
inJW8ZZ6JxQD7YIqmv5oB0VAJm2ArxqhWXbf47qZZtrDzmtcWZijc3AbdtJvckxH6etHirADJr+s
Nn8R+WWUhr2J/0n5AzNBzKQzqsOmL2hfi77/TK0HhhaQngAG/YlfE4lJX3uErzKg2nvMmjrORYUx
6wq40O8IGN+bH/wyNNQ4EI9DcxpjyMmJZmIFclm2UfWZNWVK/cB2KTxt79eF9FqXAfTfrZndiret
AlyXSksR0ZvVPFkaSpHsADj2gKAI7+v/Vg0JK9L+YbGyQU0/q1RPl6qnDZO5rFMQb/md6MgMbP93
FOej53P2XcPrJGOeyM10AjU23vqbznoB+PDY3ZuYVpDtOw1RmS283x8If/e3B+Xf46OSjcwXcR4U
D4BzcvVcGCxRG+oC0yYGI0a+Tl5ieACiqU4fxP9roB0ow5+LEOrlMm4NJEf89OzR+zsBzUtlNAG3
GosGP+3M1RsPd8V8ENKVYQGjP4r/bSvNTbxP0KBfbmGrNh28hMQRDEZLIwrqzUNsnmVDAb35oGZB
rOMyTX203rPKqS4xYvqH5cr/reyr2UEgCYs3WsdZeYc0dlUHCyYERXnm82vIP3ZnsO6sOgpmAtOn
BC+vPfzjPFzgbsOohq64yxMi+jbMEOoSCEuIrM+SLWg6JKGoEMVvhHcHVLhNV+ojEfPQ8O40PFXV
xBS3dVr4GEIP4qm+Tnq3EbaIFJwZlQKUOOit9ruFkynYyfHuMFU/4wp1Vp1SgB7CxSenhaZdIX3m
VVpbGNrNb3EPjtwkBwuElQ6KqFlVX1HS+PgTfq7CVZkw9lGkGKZmEXckW0qb7ShuZPeMSbVCpon2
2mQ8MgSCTBw+36bE4CZLd3ylM2Ii15jOjE3LsBH6LUpwp9j1MKp4+7+Zv5KiETu+DrjLXfkEzrXF
nRcG7t5Ivct05xUwQNSsSvGQPd+aCfoMrz8LBrLw/kBLn9jpT22G+iGeuO7ibfwOl2iIDNWM9iY/
JmAMxvXhYZfZuCwtEAN4qDUm1XQ9bSxMLbAF9e228waFShm//4jZm76cWGRRr5kOgrvo9SJ0Gs0n
1TDljNm0TqMadNFle9IaSltb/ETcgWI2yyGSeNZICMIvDhy0j//v4cvUGPg9pMEkUMLShH2o2Mmd
biW8vAQWSKv3NOEVkHHpI5hNkR5+wEzbpFXirKx2vtBK655Mgi100MjOVKWJQL8Qby9pqEp1eYdU
OlG+hX4LbXkivJbZ000t4A6GHsYvUh72tJKBMBjVgJ4zvVI1q4BMyWqCpoa9yUB7Pyn4zY3rIyel
Bw9VgmpFKd6SvpOOnhpIVAD7bVgPNuAETHlc8Qw96rv7cShLFCKzsWSiCg+Ov7aVtIrxwRpyhvCu
oSe2Kedd/IjWtgH11VELhLdnAaijrRhG66eY6VG3RdEW79zCBMPXi1KJeE3BdI03kkqL6S8iMmir
FUJAK6+omFh3cmudV3r+A48bkRBLC1GfG6QcBalC0drZ+7QVwE3s1qElCdDA0UlvCWl9OKOuWkCk
iMDMWT0V5hkhQGL3P77zSX29TeH2rC6M72+ZlICaV7PkybThx1YLFz2drL12TbuErZSx6jMqzYFn
IaB9Fwn4gHtHhtbYaD+oCJiuBqVb0PLDnqplO0b38q0QZVN3ih3/tKPmflSOXaD+k1Iwtg7K806a
WJOKdPcDUwwdMRwMvH8kx6uSHZWstKE/K3LHZpG8I1YEqoK69wunmx0nEoGJuANbnYCtNWckILT8
xFp412ySJSoFER+RDGAYzWKAsfvnrxcSzwnlNr1rYtYXKFiThDR3plO7+F26IUsylNehELLUj3YP
DcCIqsTU2xkfBFivWrYSpVQCzpbjwM69Yy0CSVoH/hmAjsFTr9fzKwXx9REX8jC7Q3DRmS55YAvz
GWF+dVR5CDSOw+GECuuzDFlbMbIM5XAQeeXKBGiMYJzORtz/KLUfHON35P/ni9nyhRiU3WU83NsK
rQnaBL4z4wAuyL1P6083xhPnPjnkXpQofRqqHZ1a86jyLukYce+zOgGCQKx3I/V2yOaschnZnzLR
CGImcX9XuiZPZI9rx6FBQcwa1CDvs50xMOs+Wvg2NY0M2dKjUyi+5CP57H2pIazsivfLq1t/qEnd
hgVpedAE2kqYSNar+FnceFrjgoGl/FI/t2GXHrUqQ2phs9c1sb6o/di0xxnhOP1BI5SqAJhOPFCd
6W6G+W6NN0fklGsl1CB2AJ9ocyeL3LNpSm94nLLwRuSwqfEhQyzpMy3mLjclXrHChYt+8LtrVdZb
rjowe7se2/YBmar4g/izmCbQ87tOSsDPQ8XS3iIKBWEnm5KkkqzzZFKBON7SrLsCbDw0t1ID6FBB
vYfUxEvM8BUN/twZlgO1ZwDAf1Q3mQ1pCugi0h6GfxVmftlM0chDTjbh8+q3zH2/s7d2DwKVkuAJ
QKor94pJdX0xwb2tTyhgIYMmIsZeWEGFt8g7HH64HcihLU70fChztpDV3ozU07NOsuM3azb+wRB4
3qdP9Sdg6i53Ky3wdOfjC15yAcoHkbpBKxXXO6eaLfK2eqN0eLTOIj6UpPhueFsKDs14NfltNhVE
Du0uE0SPPQSVi3CSkNdkOxRllS3+iqZqy2GqD7ec5zxJfl2CboxflZwIPUtBS9VEL565NCPwJAH4
3VI5gtZdWSvMIU38fu5DCMsiLRDLGCAHpZq8FSmcid94q63upoW9iMjndHOU/PAMWO3/D621XVe6
uftjMKKv2/3jaQ4l7778F8k65fPMnuqLHT8PIESpztWK+JDKfPg928cF4YpMsEX4UVFcnqLprdsg
jteeQz0fe/57lyCNumQr8DLhM1cfGiXGtk+5grmp+KcGvFA6TRCm8/rIqs0nEDZC0MU43mcQH7O6
NYmBNj04YM58RBG3ki4bEkVkCxYNgL2li6a7bPVmPg9m17YKyqN9OXNn/dvq+F/wAmziRCc/1YcR
MAYaLbknb9aj/fB7gJ6Efp9MZjtKctMim2J8MgE2D9pij4Grk1ECCK3IilzHOs7SDQ+9yMeHvEwk
8VW/E+5frMSVwzvEiNxblQDG9mCfUQbNCIdUI9c5h+05FmXhfhOQxcnE0O5oPKkWpCzFUg+Sq+qY
QRDv4Pq87Tj9jkRPQexprOo9lVRf4I+EZpGnX0R937GVr90uHS7kTiY4+HHxTdPfNYJtYH73+gjk
DI8djCMT9co7cu1ZqvtDbCj/b0arON+LioqKJNg+lvs8QFNxj0kwH3kq+0UthO7jDag7SNtTC10g
lwheeltmpiYdvjZkAWsfHq1ZVJLhmQFYE5sUPQROIlHeSKNjDVnhBbdv/lDK86t7FkeHgFQ/ZXNh
+OLgOWK0CrJXpoACGvkY4c47+h9PPnsSqG1ESukub/DFQ0Kk0BZ3AVGFXzxcpyIowE6pme9BUzhy
CmVKTZryCA2PwY+JnHeaSMFESJLp8MME0dkacBK1g132S4sXsvMjMpoPZXkSO10kUgqRQFYxC7Qf
2ekRuQLNeF4MycLIDZKx3vncZ2oMNs5jkO+mlOzLxWHz8ffZQ0IXFZz6Svqa7avs26pe7BlVAduq
4Jdq2eEENRh4up9fvMs4UqpS5/G5t5uNgrkLhCaJwe8idPeJ20HjNFVe0E1fxQ/VT6hoHyUL0VkX
iukLN+XoM5VFQP15DDJfCddLmpdUqSFyMrPE73/92jzUdrm4SxcO0j7uqz+4F1VlcWKTCecRh3eA
ZLuUPzhywk+NZiVaTMSt7CNmyhu8smabMa/VFAbdPtpHRCP7PyZB1N6RaQQxOC0mZvaTQP8Rpru9
dUSvNSmcYB3UfYuhhlrsLfxr6I+cCBAB58VBcUdpgXnyDqpaIh2Ujeqwu5pKFi37wIixvp0SoPEx
07G+sQKmQYtyLEoSFO9gqJygsBbe64JJeBx4rJS9jYFuITYj+BjsTpHuoQ+jYnu98v7dYSQGxkwP
T1mLOm5sNEvwca5gSFC7NNRaJwo1QVICeS93j3ASw/UXkrKd1o3TIVAEI4njlwbfUkLQWuqSY49j
eHO4bmyw53PRk5wbKid8lI8DEk4C7PzmvXQOECZ+48zH4dAAXQJGBEta0lvAvz8b94Be/lWD7mxx
4rpblhd9DT0RFsyAu3wanqEuWFyTL0EwOrYaUw9eaJq4Mlwa8Ijb0yW2aIxBCxoHN3USvRvqof6A
MffNBoBhJmBFKfC9Bu4oI9ESEA95V5oo4OBiVya+iTJHcUjW50Jk9z4GUzkgtTKjWwBdv/vBQhhI
aPkCGfUUaRGM2U/7pIj493ak7R1eh7CULJx/1OgYaJREV+3w6JaP5Kl5t+pkUzonzpSdxdrtyfxV
UgOCXG/cDwyjUBkF2XgchYRKpvNmnZzblw5Cwbzc27Mq5qh2RYQAEHu6VjrQkC8e25ZTUrs4VJiW
IwL4yglQAviDZgHWjZfKOv78xbWsugA/urwoTr7VJLRwZiR0bNFGuIMtujcOthSu67vCI649KRha
MvAp86tMDNz/Zwi1k/tCEDhimR3tYFxlPmpHgV+v4f1oHKWwnCaWPBsGB55vzrb/aVWtdNt4U8md
ikOHy2SJFE99zu9yqyX7WLRYolvNXYThOJnZkWHzSCpjsDlA9gLAHT7P+LJwd68jLHj1MQ7Wr31h
yQkuNo0cbveqaOgwl7FJoapVzc3+MlukbLp/kB9nD7OFkROQ5mzumVr77MRikYqQUB++Hva7T8HS
KH3J8+w0kLP2rue5Jbzs8EYUODtvx37VczjI1kuvkMvuMpZ0/6yFr3q2SXikeO0dz/cQ46KeYBBA
SnSv16U8tzJsvEJ8JJnNQlEI2NVGAXqQjxsfYd53YehkTjhAOfobtGpJUKMvs1d9/FCsf0Z8mrRL
CTind8CW2WQXP87q5b8koG/lbWbwmqEq3WgV8gCnVKcNSq29cuKZ3hp3UPqM7vwhVT1GMOc9GjXD
jfEgmpxZxLmn9jc/HazXRcbh4BTb5/qJWHjl6oSemZM0fOamYsM7Fa0nTuamUEAbZi3fl/2PEwZ3
4BDuBJfrpPr9t5r0AZKEg4EiiLIHLY/oiG3lShNiPfdtJez+WOCQ8d3aLcvnSpR9IgdDQLYKPjMT
pY8unuSpkBD5fkvYo7MWf4z/tt/BwyS26eTGmLCSGweFalpnVvQeaT7DcfeTJLwuq2eb7DQjePYc
5SObTePXUSEccJ6W5oF27wShJBB/GQrI7sDg+ANzhjClRGABQs4awId2GM74lSVXmix5kL+3oVIA
ABVaFDZCXQDyHNcDM+G06TiUnIvnHE/xH8smiHT3dQb6g80XvzGqaCBevOPwnnaOi/N4fqOjUjiv
gBwzQI93p0v7piM0o7RAQ1J1siv/Two5v1P7Fp+YiT4iKINNkL7d1fAprTLH+0yBYIeeArtYDXNU
MSbQXIE294tHp8zvei0m0Q6gO2MPe+oLMnaptVlsljFwM+rbzyhJzunSvmQa2tkq1PGMZHa0qDUf
CsmrCoSnXMN/GRG4BAludTkJsS2zjdFo4Ho/TlbFrnqV+lSz96VKq6dhd472eDtTE7UWT6ht4j0s
eB3K6SpWcQe74xFezqAnqEQQLfUZa4oEtwZqcP3NxcKwfw30Ue4mPpsP/JwNyNbxLVPJZxw68U0u
qkEUyWKUKtbEqu7xXlZJczhvajh8YzxY//dqgkGxfx1i1IN+hdtGblQgjVdvsSFfOHGvNRMxNc+j
CYk8fnd24E907rwiReZjOZ5x0HXy+K3bLX3XHSIYj2WUTlhLc6aT5h7FfAXMLS0YKC6sPy3omQ5C
FgQ8cqr2fQvtmOStEQTsCa4LwShWAzDBMORSv7349EN1+ZZg3TgY4CSlcrnBo0LuttpgnjRN+tbD
LfG9Q9yUWvE3OigAqXSGP2o96Ure2mXTe5sMSjWc5/P4BH3z0R8sCkO4PyYIuswujESIF1x6O5Zn
tig8NW1VG5wnpEj5ak+vdErimUQfukXqR4r4NJKcVYjiRln56w0gWzTR0RPNzI9/fkXWGMWz5tvr
J+p+hWZx7LMexRiwaKQHiQgbCpbckWIC+PWFDerhqKX+EueUn0wv2Pm38R5VLxEzJ5upTUOKai5A
0Zk/hwlD70mZj7RhDUhvBNIIPEDAwaTvWLv7UoJhdfIKC+dtANsi3R1hW/ZrpCGjrvVGl83jEY9v
XuiNC/kE6y4OlbZsgNwcr2+wGCtyFh1cdF1BqCjhQpzys3JoGhC3qF2kCN+yC8bDgROl79+VZy6J
TolmlW5xIzDQDivUjAKIXyGl6Lsdh2qK7/1wr9tKBM5nLLQaEzFfooN2uPC86pvnwF6qTcd/lRSj
4R76iEmJB89z3dUCokK03HamYTQmkIloPRRCl+KMzAyRw1x8XeL9EyJdEyc7D53Re9WdrRMMAh5m
Ua8pgc/TNk+IeqdvcvkpTWF/+RaP3VmwO6NQbo+GjjMxhM79HYJyW5eV0lHc8wFc/G7EnpJ9hTwU
XJLGyy5kzGrjmUo3MyqaKyRSAIzbe6VeOqMnG5NtqP9KMeXQuaa9gsLxXnaKk9OwCGy6InsaREUF
ocZb7wFg6MIbV9pIAe+6pg0KVCoJcUQiVemC1hdkCoCiWzV54Ohlz7NQ6xRVHByvXJET821eOW39
ycSXdQuNRdyt2JwxtTQo2yZDT5Ru6PA8dnMAkkvJidU37wdho3y4uQIaGdHEt/eW+dESFfu6eaAV
HRgLRBTMOLwV31iU0bkGxRIdtnn85NBaskYN/NXHTzUHmBoXvPLM06r2J4NVG9w0l5gfikI6RgmJ
+Vf/mRf8FJOnyjFr1DisogFrObdZlyljUiXNX7Fx572uKaJfRmUkXsZvi5HmdM7Utd1dwXh10UJ4
mhfyeF9v1kkfE00Gt0PLj6nRJUl099HVWU5EHGG31Cj/FEbwFcRMtzJqVVd+ObEybtMfDzI6zNOW
/IIW2uwLCQwbJHXHuFriQhaAGElL7a852ujEHoOIMbOAdBN54MgPNovmPEFgREZMlrNQq3U8dElC
roY0Y0a3K9TvRjVAZTfC8y8EbTc05U2xmXEUHSKRCMkMSCoSpTyqqmY+sTR8lOf9BtrMhvmWQ89M
4FVppGvHE7d9Z29ls500SrQt834OvYQzBSblbeR42rCMQRM0hQ52iItP0ul0s+VtY9EDQo9IOWMX
r/QYcPFROGEyZB+SV0mK+5Diy7B/YUCPPfkGuKmZW/wGmkeJX3DVjgfl4fMJ43/7M7piZ5agMp8P
CqRGbP35A5U4pKrr3e83VjMKCeNpYj/2hgneHmSW7B8sSgJvAgrn9xzMDYk2vlDTRJ0an46DyqUN
35lSNqbgwLqHGVPLspQs1qYaq6E7Hj6qnIVN0p5CkSaI+n7nRa74F9BeNeuuWMh6VLmMwD60FfEi
gSlZdtcDh6+4XUbqwxzbvC/xzY6ewMFWHNY+P8cgU5+K7VpAQGShL+NL5JKxOxkDtLFAyo0RlHH6
HRPHLQclD2gJ25nRhn69y1hNo9pRFd1zROIzxD3oQ87vgZLyGGpFwm6OL0nupAA7OAGncK4kxXiv
GD33sVZpFGv3kEycD8n2qmNEux2GMP6Eu4W19knEjg6xQXf213NlQOKsl2ItTF9pg6HZgnf8bz/+
Lq/SuaCFNyD+YqyGTtvYrBw62+h8dEhPooL62w4raxEVL1mSprrHAP7/OEaqPLR5gFy7tR2mOejo
D340ci+0AwaUajH9/8DcXjzkEhWtvgqJPPVXnEg+zMATlQgEGHc6OlHs/+oP6Oo87tUiDl24CJNB
L0s9bkK8beqvkPYwn32hOnFAD0E14br4RClcMtTcG5hYQS2HgpBQkmbSy8kwT5zlbQNrRqObiil8
sQY7/M8z+ep3vPunDlD624HebrafljCCsSSqGGk1EnqJlwq3GZAKaUDp3Kqbpk94B7I3wm3Uwda9
/EpJwLFTWOG1nBWcAxKPdCzYtr0VnG2T8dAXyuuUPFHsjbJffG2wzgFnBXaPAC5Rpa2iDVBfFN5/
TDoARB1gLMXNF3OR9yq7Z95+p4YsyqzLu5mugxlNhGp3hugVkQNiigX4D6Shysgc28O0392psPY2
P1Cw8sMao+3c4FrD15HahQN6ftvAx7c2+S6gdRFaC/3QXiVBmvV0ATu+tQTAjKAUCj+g0g4Y6wJ9
Rsu9lxkrnOy0GW6N3y5ujD3qs7k467WB3dzk158vSkP5k9v9jNMfuQtJf31r7rRTl2ebK76xN4B+
7fvRGQjQlpXXaZZ9eciFeD6qcYTfg4umrtGKtvnUiuqLixiVWE6/FAPdXTVCoZW6/D5CyI+IP7mi
758mPOhifQfEo8ShwMqKpevylyfZ42B3Nal2SYJCtOyO6uP3sO0DV57r8KvW4TJYQtX3YRK8ZwS3
xjwap409pQlS1+yCdOWoDCcHxrhkOsD7d+zJXPTtbz3t/NFEUb8rVBmXqiT9kOILdl/qqGqxK/ER
q0A7R4V7BPfDQDtxSp3lWobrmwP5WOOQCZRpLC1johvOUXe8yLw3JOrzcyjxMg/tzhP4W/QS1Dst
VkADmUW+57JmxLQ5Vgh6K3tjssFkg3EoNl1dgw4qmxANLrhwGF0lPWyQWsCoGJr7yjeEJLq3l7oi
U/rr3Yg0tRHAKyoHdl1FXB9nXOwh98AKd3oYoPwM2L37VhebBxemL9eR25r7adEhADcm3rG9oi4M
i8XCup8VxQUzxDJtHeIwRxtfXZmT+x6xFcsf/HhjxjpW92VEvaifTiIfsx2EjQc+y/7xfmoy0ydG
KwFMze0fU4KDaBUrLDJ3DyFjaP/lUvUfDHxnLDFsa6V5m1dh5rMI7+5B+2Xo9xgKxicGASMKxKgL
DXftQPRh3YZ0Fla523gGLyeIl8pR6v+BF0HMWG9CwW+GgtK9FiFXNlHO0ODy46sbe+PSRiUCOBNX
8TBOvo6IAEqT114e4aEJBcYDPJ2m/+6IOn24hg4HcotSugKf/FyLIi1wVxNlT3F5M5qrWbk05XEF
w/uzdr3sR0xhAArTLnerCC0D443xRXl3jFqlhJYof83WAk7JEKPgmeMW0bx+mBB7zkFs/IJp6cgb
D63SvMLFWR1fwjZyXWY3E2+fs1gf7/0WdzZVNAgObkFEiLt8vteLO0WxuVjOWAxz7xsA9gIobwOB
VieoB1snwHK/+1BsnsKkLOtKTp2tM/gEW4LMBFSE8IIt87LRUGL1o0PQ5P7kkwjKzpMDZPUu2fKs
6XUsGzQpx91nldCw+ChiZvXbRNVPvOjhu/BbOsK5knO67ljUNaJkRZW3HFcvXd5yv1tveuTOf9Q4
Pg1B3NFjopPwZQOi/7vjNcbisoxYPLvwHhScZhDewI7xSAQyaiNsEUHJisTwKm9EbPyR+zQUKzzM
XA5hIISVxB7PR8dxmWfMeMhiTuGtBnS1WPywXs1mbNBhf5rPNMUoBAgyZsSmzUlkj6fxva/V32Ha
CnVoQ7PvWUJKgOAoFMaJfmy3+QHQJrvKv6on+QwKj2oeD3AlhIBhxuSx4KrHdCXBoLtBT6/CM0WU
f4T3z+T2ki/XV5x/kAl9SjZ5VZp3K/z/Z+7tjXpJtoFWcldRjgYspiQv6Dk+uMT196OwAsWRj7BX
Am3RiDCgLB9TVXgnNzftMSqVP7H0zgxwB8aY1VGqhx1liKZgo5KF3j3L6rfDbMP4fAF3rTD+B623
5GQRuZ8pGFuaKhYaatLVCRo7fMOlIMWmVXQKNoC/a/7drbJexJhI7ejmfZKkWKYfTt5Nr/80VDal
5lcZhNttKAfVS03jQSIpXwwooUXlAU5QzHymvFAfgZLbGixPBSGhX2DVOtaWwy/4xqSIcxVxwK8F
mYjIPKdlw+ngtGoqvxg42AY2lMdEoTha1KDP7gCfOb/aZYHMovMKXh9zhJIeeJ7AB5y5gS4NraYA
lGWfKY1W3OlhbYVCJpaVbkAJJXFFiZVZU/gCWFkTiM4ONr5qgMPpdJHqW574xRW9FJZbUd6j9Tfr
a/3z1368dHWyiNGr3vG+s9uG6BRt94OlqwNDXnQzrv/J92EbzglBn+wDnyc37hwIKg0jxaoz053l
ir58IEel3Vrosvh2ZaCapAgjRuSIcqxvWTzm+7DzQppbWYe/GD68OdhF/DFzwZujd60Pcrxy+UMn
hpDIzOHPgTTu/Jj3//sUoAjAziF3Uvkq6ofZKE/VTZ517uS/ey0uZ8oZthsfyKUhEove4h7+ogMO
AnZLNc+HefDHVRfcXs/tnYxuiZinkft7/1L46WbVJFF9JbTVLtLD7p2cHDbN3XOXwsZDCHN5NSGW
JgUp3rVuViBcGTm132MjaoH+32KsurKMKg4NjieVU75hgdp11oAiT8+kvq11iOOCKG+qEIJu3Bpj
PeUcfuiQRyFF9r9b6HRlNo1eD74aQ6Dd9viwrp5chAaPW1ogGgXQAw+zeHheFhKOlVu6d8OtsqG/
GHZBxDX6XJauo6+9ZsY/tyud4zpx5s78IvTXub39lr8DYDyKgZNbPAkEgu5vHI/VqT89+o+31IsE
vAba6Tx7gN9Sm3pWgjsBIvy5RFkqeT7gULFvDkqA+5484O7ECdvdWdxj6UNGSKgMKNboDDnZEW/r
t33B+l2cEybsrobNuK0eEL+WGUl9g8p40F3d4uPNTYDaI0nPG11bySkuUismIyFvj3pG1+0IE5I8
DrMAu2Jc8fIMpeoGYxJjo5UVsJpj+wBMb3uzXycdqrpHV7mwCQL8i1i1pyrdIjzpbvR/FRsTqkkH
HbkKPL0dJ48c2gz04P+ImttHFqs1TOp+i470eIdRmvEYd3kz/Rd2Hy53Rlg/zxgsddpQ8cYY3smG
aXqHEsSfqvIyTLYclYZd/OiZfL97MzwQrJM8rp+j5FxJFjZUIHNzd+u1NRfyQcsqijDycdqQCJDi
MKGYt6ZFZy8h/uqKwqFHB4IVCYT5ksAx5fOi16fqXY5vi4sGh0BcBoisIncdrDe+Vpe37nf9T5zt
2Xq6lhPGmh2RlPujdbRTtaiuyyb/821EamIFFxJBB6LP3gODoy9Tw7fseTUe0mor+ey29d9X3D8V
6E61fHhQPEJ2n5GAjqpBngvNLRAxFDQqQ2BHfyjxJR08WhEX3prfx4+8kpfoJA4zp1pj45ebcGsu
vqO20vGC47aAIhlL12A7s7y9QNRZ6y4ORPuiSkSEPGwEjwo30rsIKcDJGTyD+6hpDSnZGAoajQm+
/tUhAJzKTEFESRNdwBX/Xg9M+qfzyucNLEpY3bnp1jl9oJW4dB4JNmw6aLaQbKb849Yo/YFAXWO7
KHOPqFel9F2xKoZlNjr/AKpoVg2ORauYHZ6ihw/0MxeBacQm0fsNp2OjZjz5ImROSExm/Y02uqvw
l52Z0s7G/Xlz/uTSIMyXEhFISvkYD+iQyabXOtfOtmXwPC2TREvDA6KaQKqnnsogKPLzwdcgkCrD
yJrnSI1nTmIhAIj1Nhi0PKz4YiRqjzdEmGXov+lWKrv2cWOvsB47CkHi3ROUH+8CVSqa7kqvZeZj
RWHNUuyMyTq815uMSkh6M3dhyp7wWwgXIzvOplObIcRM2G0O2oDeBp8Ab27TtgT0W/R2LuMBF3PJ
i0kAk+R8Ve+RXYzYirjOyyyNKHEijqr9ISSWoXgcan+x/bEXqBBBOM87jC2XVSMlq1CzkrMHiuLw
vT7b86Qzb1B2rrIH66MORzQJTmn6ukzZeQEubclvQfKppPvf0n03b7AkEn5Ix9aKaH2jTsr0K+ap
ge9VsLAx4mZ2k8HyjXOYM+HO5wQOpToT9rAsRUkxjXP/j1zIVTY0iZ/eBSd95CcvmW45/OFiFR2R
6A3dXzQ9YxId4DC+KTur8ji9XEg1rALLhP/dIpYG9BcN4YIfFSov8bQGQBzPS49WUZ+dIZOHy+tq
FHfhbfUB9B8L5HHl4gw5j7GI55yufk3jGLeeYD4yjhTrNXD0t5USWSl9PqvYmcSdT8S0rJFidulA
uVgV5CWl7BTy7zO0Su8aM6pczgIoSwoneyWpw/MoC7kZMXdFY12rYIKOIDdAYi38REzD6PSB6vy7
XRHrft5jn9iT+JiodKORsYdvqaRzRAzfPIVi2iX2+iyjHNe9c7tT9Gu5rbpCg25/aAwoW+NSgOw4
/d8KzMV16+NyQ7H37RFGDqP3//IBnhgpWgTqwHw9FMG9T0OdkNqiphVBngyhU7FT6c6E015bXIBr
5rVIUeR/9LLiZxOAVSn2YrrP1xR2rdD6Rs+4xUvLpAFw6LoOJT2LgCE571A250ee8jebnhpzfjTH
kEagzg6NNuMYHrQR4RPzM5Q4kxIE1xou1cle2vGbBOmJ4aSBSvvv5nzJYlRllvxtMB75sOaJQPGx
9xK6eDFo/ltFJBbDCGeJoh+juHPytZRHuJoMZ13kd7EZiqDH1ZnaC8U4PJeKJjWqxCsDpzsMUrGB
5XIm8ILTC67AE0XCGlfIks6GqIOY2+i3fxeHfnZnAAYhWJ8WN+M0JarN9z893tLHKQdVbHULpyoT
yqy+nYfUWNY3hF9PxZKL3s9KbeTr2OiSqvJMAq2CYpQG60zawwKVC1QFWgvJFLlERug90V4BCejb
/odt8ozXtXEtWDJF8O/Yv4B6ueGHj9sCZiN2TzJPbfQBcX/W8lR5YBep+c++2QDMtjUp6oO6p7+Q
XxCmPFxi7oJTCS0JqHdlrNkBP5MAPd5QSrJ5guUF30eG4ZULs7T0tb0OCXYug0aX9UZw2PcfOsm5
86H4U45kG3XxH+C4/S1Fqnsk56GvAUYLueATNnm05zR2mwA+IuWbPS55rAWgcrgYH29Mfa7dOvJC
+QTWzOyMTqSismftJimlb5fO5PastpPykP2jqZSHMWGnggtGns6pcRyyI3KGW+A0Xi9fINd3IbVq
qylqcH//aQipUKvHXmyFqt9jlBA8NJRcsT5XMYduHciwtyp8bkCh0pBRko8CqQRGaoO3tZNptHsH
O/fAbW8nHYUyEk+RyPTG/nv75D5mvbGxRKW8ry4JlW91QbA5QU+RIfQZvITLoVq84/0Opdby4bNM
zHxclwEIGxbHg4m5l/q7mo6an/cXTRPcLsqn0mpNXdxLXLBu8RS8AZ4MJJ0LhiPtV/oCAcG4Pa0c
8ozcjJj9cXzdIDsKqe9gmFITLV3l5O4UgG388K6Kb/BewGif0HHO4mzQmNwLYQXoM0HbDXLtsKsT
qS0DARIps+foa3il3luvayg0uPt/rsqrw0hC0gOXapqD1kACVoA6g/OZiDnpLgquyT/VDzV2PozE
YUAdMX7yjNmeai4RUNGEthLYO+Gn6gpP5tDwbT7nolDWUzhHyuApG9Yximk3MR86DPAlmdTZktor
GlKT0LBbCyfvdoUQA4K+1E+bQgXw0QKu/+9POOurVPs2uwjXv2fhgs91NIX9bXdrXKvHrws6qXDu
V9PvzbaTm5nAcAgw0WbYCH7EkBWD7KIGAQ/Rpqk5VF8LiVsA70y1Xjuyf+1co70V2adArZyM60V0
HNYNUVQeJTU23iERyNGBkTlWUgworevPqdniEo42UWqrjHcULBdkE1agQ86Spv9CwY2kp9Q4auMk
7pezXH3w6rRa6WK9qFOm+P2lhSCaF5gEXAFMtTYubnd852j4CUavKWPmRN9JOXHnvozDKFO6bc0V
10tBZV0GDtUXZsI3Kto6QlmatPakMCHZhEHpFEnnT+uxPPw/f8t/jF3CrVwkKNincgh6s5u/e45b
v6CrRtgS4/VotN30pkzgixeOHDa7/z5/BpBzp0lAloZITtRH6NnioF/quGIvLAUgsbP+6PmPfiAX
bXwDfhYya21ZxV1F/QI8kSQWLYe4X2fsN6OLRB8qlv+h6NIDbGUReEACekcT81COYEjN48q6sFaz
rQXSW4YSYLRlzDPi3Qgm/FyohYVdDLbCfQDXKemCQWRjx9oZPViWi8ctTck6EGATdLKIGXm6Q6gO
7f9zG7wpT3vpvwqFBlFXyvWRePRABCRBNc+vjdFATjvQYCYLVX5c7WfRgUo72LrBKohk7NrxJQjc
c5AUV85kAVKrLe6wbW6wNbgIJYNyDdVUf7NQzt1+DSLicGN026V5Ze87TnpgvnC1utbljo4RtHl7
E06DcbfXdf9EvaFnGDUoSmj87C7G3VE+plxbPULM18IA+oMFB4bkCaz90QToY9BwcCW/uIwdMj7P
jlfj/bjWXIcGVsHtQ5/fD7da/343ThMylppwKKGY2WIpLt09l2vqwE9faQFWeTFrv5bFVK3dwP5e
A/ZbCrZ/y52k+UYPicnPqdhI+gBzX+Xfvk1d2RHNma5R2ZJudIR2eW0UYIQzGHsn997KO3ob1WBT
xpm/lsxllFzxQId2b+ZeUD9i5elopSczCj+0pVyPyBzYyhCrNbVDpoQYpdO71trAPyWW6h4JOqM6
vdaD5/SGnbsxHeyKHnYqbfP9/6iPicUi5EmeUg2d780Wk5KzD1+v3ppYctCaWzgTRgXoROt1vzBd
W2rawwEYQ0+8h7n/PzqPxbG3ltvexVHRL+yACz32y+lBAQQv92rPSNjcwGRdaHByv1b/HFLGh2gV
+Km885mSSsZPyyIaS6fyKBKYUzrbRqzFLNlYWzQwDpaqGHznx/7NYmgL/kcnzVQ5MTp81EDJy4Q0
+Mu4BIVzAN8CAmHL1EwVm1vbfJYoERvej9ACT0/oqVhMnW+ZcgiM+1eRnHXk2Sa0/UONNIAYbcYT
/T0Nk1bbXT4QxLEFxlQD2FYWpnURu89v/oVGBWAUxtM7lXwO6FDF6Mz0iGwdeSKa74MFfAInM2h0
OqvivlPvbl2JO/T324qt1w4kcs5WXv24mzPCDUdvFHT7tfl3k8/00gKvN3AYiSPxg9nNnkqlroox
zan+61z9L/RLbCkF6dJ6JhcFQOFBVvl8I4rd2BgsZNKLFVyqqh6syaljl/h4AoPLuftwuHLZTnsd
vkw7vDXTLV82VHPUDP3Dugg3ob3YudWy2z8iPpnnLKLMSi2dz+bIUPotqSnMNDykdMeumq0AlAyi
PSBbaShGAHKk2G3F809MdpQXS8O6JycU8LfSzknEWBEi34Qb4hFn3X7MvKrpxGZIGFgMp82m7aG4
9Gn78wJ/dhJHLRc6e99ybzgX91ZQ/7JiCJ2RiY0KfCHpIFrucZV2SC41PbP5hHfQUH83yBqPi6zL
WhddlzrsPLljSIplocA+boS9/oAvvAu3c4RCohirWVwu3TtWc1vKdzdCB9VLHaEBDHmX5rnQ0m5/
9XxTaPSzMqSTHsGm93lD82dw3w0qvu9AZG+x9CWEIJdXVRs+bUbrPGHGJZLoqesOZAviOD9dABgk
TMYpwYK9UXIHWTnD8B85uZTweFUrf5SFmnfMg21utOsJEvgG4oKp+2LKx4mfLpGicCzPybS9Lz4j
E9VBEQEjlvolr2qs41sPT3JU/dAhyqMyqdxqlvppZ8V3c7uGD6/0IUtkEKLx/B0iLjQahWZn5c1s
9V3O9yeOjNfy6SM2K55sGxBSTrw7Xe00/9/j1rswtqlBQab8E6Ih1pxf6G9Vpxz+HM4LLlqSSiqY
8FLzqkqrAzsbN0eD1WBdgz0ebNzw0fs7XGX9CdIvHKGgcGSz5pjb+aSuKlVZ8lJOz0TKEvzQhElO
dvsMRpERGOq63lqz9167VBkqElOHm147S4sm3mjdvd70AAz/ntKuhmrAyLHS2pxuZ/WpPc9x9eeo
cD7YCxywGmB3VKgLpcADHqSeJzkq7worw64NVs7PPHeJqCOSq5fce3l6/vdl+yjmmHmKNznYlBZd
NmRjm6Z1ocMkQCtaBFZBMoUx+j5YhUGyLi/4Q2CiWYqJJVJygCYToKKC57egUIdU+MaY4VPRPLcz
j60tcOrqEUpOZFB03Yay/zeleMKmyp9ufqBHMFgZKyiRLw3wm+wU1RnQJime6tGAqE/Htt1EuLLy
o9M0k0+ewXOY5T67Vd6Xrc/HPDgiLEs2Q303aQosMOZvOaN9NHcTIU1ac2pmHjxpG45EG/29tgjf
EenM8gHmU0cnypOBb0TmsHZPbv7ut7vzOUtvI1Nx7DjehNB2s/0ivADajvZeefOzAAHatf6QBcF7
5nqsdNd41ZJE6fVdEghV4rCgPKy57/dJT5uAvPTqJtuAiv0/KrkQg0HvhE0tl//G4hAx+5kvmxM/
tJs5LgeYZRrzdVF3AqL4f6nhz52hERoyu5kGc8MvHWYPJf/hNchkNBYMKENXE11Pl+nBQUeoyxB8
iD4BheseN82Lr9WUGaO3SajI9+xHYxi5a/kF3XYY3UuGlihvKmjSXcTGCzYVkB7jEH3ih7N1gmRj
YIXRmgVa3yhQh6T667ubWsmbXEs4Nbln6oAaqbOCaanEixANiovYMLPia9OFDaScJfRsCdlPBXUL
gO3OyGnneMwSb0Mj+2+pCrkyvT7LH7p6W5rTE0ZA4uruPxu5bdLBzcUxLdT/Cd8Ofw8DW6fVCm9z
3zDk0/hlTQ1Eh5M+ru0TIV5Y9rjWJBpQGMM4G8+1lGiwfAx2MXWJ3oUURHFHwefFcoIa9RXuGkng
ki+eOWruZtJWZiZJqCLNoUDLdXuIp/iffJBkDHJlt2COsdTeAkf+8md3SiIbho5pcjnkzgJkdQ0O
6MK93vVhu3q41GG8CweMioXlfHgoGS3qFAgZQOnRQ2c0tLoAKAtyO/F6+eTZCcuJk7UKLWK2fo/T
q0IvLwU2mBUk6xJQ0dCsNKzjxPCb8ous0IfIahu/Jzi0ezyFEZYQP7qsLSlatcaDdn16j9CBg5Lp
MUByIrolux05mOpyQCJeV17HnRs+jpY1IiE76u+ffIpebWb4PDrKfbi32N3RT1O3MQWQECwTjwkK
vynsnFumhqEs0s+UW/UwTrxVEaSCfQoKHFCNPaFJj32VIvb7G8LoivrvYb8GYccVc2QXSn2U80wO
K629Y4zSGxQOFICPRcfzoWdkBqHSVFJLeqS+Kwwc3xECoYkafAkL553kjKeyI6hnDeAaYcBC6TDG
eGzIY8L2Zs7CAN1pXlrwdrDSdScsvvIAwMfiOZVtj+a3bSaY9aone7k0mdMij2dLVilsT/Hpt34l
wM7MYFkbYqsUm4XnJnFd9WJK7AF4Vq5oqEQwz/8OoCGdi5qparFPcPkrxMiR7OG9jJXJocYd0NnJ
1u9AZfTeky8cOfaZJx87Ur6teX/ZfLRg4xekNWxNAOHcNV8TBgC3x/Qgboxb4y/znB5FTwYDtBsT
C+ODSX8obRYRx8Sq6Gfn4sbv1fQexg8idWdcC+pjeApojWQADYr/bN4Q46BOFnzq2Rl+EnI0c7rU
8kakU1mxVtP1L1KhOFE9wGtS5Izm9BkbuXGeIrJznV/BSJvARPYoW//8S/Ej+5mVANp3AOJYh0OH
oaGKbCk2G8MRxkc3M3WOcVlUWJpz05Cm4ztzk13We2X8N+uVAJeVZaIgLGsOd5xYHk9JfKYqQViF
ng4ZIxdxOsFsIO3g7/nW0pHYqflhMRSthPVw4e4k1PmIKnsrY8r7xCx9vsCJo7hy2b+3LIMffyYG
UlG2V1yZsgHd1HUp603uEUSqHbZUioDZJlWDb4c8VoHX78s92UkWjIbBuJBN1zAeth0jtqFkL0uO
q9LoiSbK6cdpxdPk3QST/cco4lrKzVdOvuc8evmMFgp03sXCF2Im9gtjUCIbHCFvog/hMztdQ3jU
7tnKyVdSUPHnvL1LrJ8yu4SOOz/fH46LfjoYrUJnRQTo12HLfBfrzH6MxnuvFnRTdBuH5KL3nqzs
nnBqrmAx9gx3FV1Sx8iGLFCG4QgAOKs3X9nXD7pVZr8qRBYAMf6tXGI6vaiu5ZZGA+b+zr/h21vE
saHZZ+Dtyx4yLxjMKHxkGPZz03tX5dPyaNf9i/LjqiIlfA9jOuuxSULW9JhoucBuQdD1MwfRXEgH
Pmtk0Bwoz/+1CletQardffmuKp2GsRimOT6atmKWPO0sAcm3O4CnB+WXpS5dqyMxAKke5tovHw6S
SEv7yvF3WQnfQIrRG4GTA49hFkP4q0riE8N59Lm5WFIWjPS4f9GSqw9PBBsSYS00uOXKIm1DFp32
lUv+CSFwoUJ6oFNc63nTl9o7LydZ2aZtXkV6z6JUsgiYIgXL046lgtq02qyraBjWuU7nC/9yQ3js
jWC4A5EKIcD8j0YJumQ6Ks3tBnFPQC+hZYSwOooo2g5G2v1FJOxYhSe2AVeMaHDoUpIs98q0uuSN
Gw/AwqdqGVdyJ8CZwcvxeLIqGjLh/njT3Y9IKL8ewRcd9OdQOuRVjR6bo8yFqcx4H6eqUcHBiBZQ
Pa6xxYMl1vtbpSGn8EPbu/PZDwGdzx+RSfWpflfcs4cRTWcXoyL0oeaxK0aSFn2yQATNejuv//w7
D0sAp9IqnG0HpLb18zaTDT36aOgstaS8GPfUGh9XgE5SJlsumEjDRzLmZcN72gpHkhdPw0jgjnyE
9NpexbUIm02jjyUaOYbBWzYkezp1fSzDb7y3aYRHw3myOz1OkR91oxwsQt3uSKCxqanvNjaPGIny
3JqPBmsns26+U6p8b60HBweLNjDHJXNNIBXLWt0B5rV20ZaQKGm8ROdpJUzcvrFW5mXVGz6iCawG
9VatbNcfon2nU0jYv2uVZX4M4iQO4jq3xrySgzxIhFdt0FYyyDxrx9u/9kulUe9jmab7Ek08z1oT
KxxIl4pyCUKjPvdLeCoa8ZZJplB8glQtXnzuM69D+lE9n2vyeDgx+cX6z1f/Uz/lk1Ue7dxtPe03
kqGnXPEAB/FaxW5XJqEHHhUm9v/eb8ciDqjF9o0Fas8XVLF/7sc9Wk1pd6ngSIUwCNpi4RwF3/86
hdm0ZujwnEmrb/A6gt0Up9GdbOU9xZNf4SaZtg3CVeUbHOt8nZupWY/dIpuNizzxc2jAUb35+hPc
Mi1XStx4C4agJlLKzntNloBcO8Vfi2oYeib1biM9BmKJSrhIl+Wn1UE3IKDBKkxTQ4s0ZDdRoCYT
qcg+9zVTqcrnnPctFBXCWI4SiWQ+X/g+vFqYCtKG0Idlm3gS4CMsHXpwzO+8nE4tzVkierOROv65
j5ZEDBuqDpK6qZeI/oECzvstAJ3KalaB+OazS02M/z6b3QyWRetpbGYFbcNHhdnM2VY54M/Ab10w
554uefASia+jRqZ2g6jc++FxHDr5roDXBR85AhLqCSwtqBCa3ZzbazflFbM5vM6CzvcwPJ1ZoClD
H6EyhEEWx6ZAS84/dk3IIT6JCtrH+xumlAbD7Ix/mCF1IpyZBIXE5jFmgpgc15mf0bhWRhYh1WAx
Y3Vnt7b/uGX2hydy4toaV7npSgXXFZcnSal5udXwmiFVyix69P9iYgyL5Pd9m9Y7zs9xwEObfF/m
riEhPFyO92NXt+uOHWGQdS5msQlXCIElW0KfOfFufn3VwDo1vZ1LnrXvXaFmdkQ0bpSbR+MRCw4O
4hTRR9NC8LQjCzCNkiCxdmHxmYHuJ5k5DSzsQyB/6byJqw5/z6U6yRSynS+EljkjQrVJbDzk78jL
LGiILCTVBd+VZ4PEO6xphx4GWkiVFn8uxbK855YY4WDcs1FYab1zF9ksonIDEc3j4IRCg2Ncdew4
peU+1XcFPKJWvS/R0IPhwoxd1wsCOieghQmhrQSSx1Z0giRTIWU8W7Q1yrXJJpimDYw7XnToZAHD
/p124UwYkfyLg1nTzMdYqhbtPLyyHTBTOnDB4oIt+F2raD3FdBEa9+iGgbu5yTKGIhmfqtyQjY/f
6QAMtuZGtTCWSb23t4eK3Ke0R0TZ/+vfsMGhGV/cQAcmnljF5sYFHNGbGoBjISZMib2PDfYMVp5q
LIbLPihy1pN+imrFXH5gTqvtXAjKYwai4jBYyqp0Yyv6TZjyFXIeBhwQdojJ5OFSC++r9u0HPVyZ
rggUC0Le6pDAHGsWC0cA77r2pi/hqY3DInJJIgMPia+dKPEIMAa4s/oljtBs9lu6pSUau1E0VFAo
wiC6X5sdDDz2Do417w4BmV9CS/wwGbyT17diL7ab1PnUQ//LpYjKTfhdOOu0onpHlihhwQc61jiO
ixtAmYNYZ35wWVDKVXONRUpu2lVqH17og8f0K4n9Rgn4nfTmEUGKntP6krKz7LrolHke5dKmKvnT
UKnhuevXwS+18hy8vV42Fjc24tWyEqH/Wap6yhbRHvLyQ8Er+Ng92AAlsvm62arg6PCpFNmCI1DX
nje61O4hJoCMfIwum0zhA1RHvscIKpFNeKtHphuAZCglcM/Lf7FpmibfQmF1YZSplDMXFKHARwdw
LJAvw3KNzX0KvnLYUpoydaARI0xmHCtpiFRsLtL1znNkwxruk7Xj857W7Vz4EzPggiudvIHcxFIR
fOJDuvQZQRudcNsaPsGMw8GFRWtPnZxO3y/lFsZZ7uxmcnSs8zam1et7zy19TjLMCws5AmBV1we0
r4KWr3/vksKP8uNI4Dt3GgvAFk8HXqfF8VKdGoJXbvfJ2dx5GvlPjYgWe0XYvycwHHfnUd7h+WIm
o4TpQqr/rfRD5Mozed0SPlenPFC+iPjz6f1PWy4K7bwQlAL2S5hch4xM1lnZOi0FebR75q4x5cpL
mV+tPmluTMNyOP9bWOwpI+Eo9iLI9P9vpocF5k+pLQAF2DjHobvNkOxCSkW3MU+U5s/EmhUWHBEH
srPDC7NXsF0o3J+N+XF9/5fN8DGI1fDMgrwUzvJ5Dlbz0q6mUtEuGCHeShgAfu8jMrxxnOMBu83j
AMrMHxULR4V9FpQyTJwJ6fNDevHS0XiFpYVzbJ+K6t8pyTlFFFC4nz+ORmMp66A6WzKAAx4ZHVTy
4jvDc8fq8n4GovEO0Q8xSdtCT+F9SegnqP11kFlV985JNbRL/gA9axKOxxX8zBCpn/Kg4WTUMFW7
QfP4Ya2M6zwKIM7+9EazqSkCGhwihuuOUwd74usekSUhCDdpl1rITG36t6ucCb3ZoAUDluJ0G5X7
xoWhlrzePShZcmaWqUbgqIF7wMqh1LaUFoBHRArKFtsGm3Ne2Bgc7/gU2KD9ieR1+j1ztOCXfn96
LilZihDud4RMipxLlRO3cDSXIL9e2V5Fl0foo8zC/grEvJ8Va4WJKudx/ngwDwyJJ+96oru1HsVX
FOid4660RjNVRNnPB3qUYeIbCgDGhHGbnkz3x6/r4Vn9eWLTTWf+znQB/vMu3TzMKnqH6hOzxGHq
nX5OXblBJg18rfKThbr1Uveb/nh/+CkrAJBoUzBwnGvqH+KMLhIqfRqq8OK8J2Zg+uENi3QvHKnu
vGo0Sg6jl/hX82J1dAakDKtx3J1XjSn5WWKX2G67BKhoyz1NaLjui4lfRVOsxLTklubBPx78Mr1W
Ap0PLKN3TBvCNH64YQvgbVY9t9W6Q7xXdmL7SK/6EIIVpV4CPuUOvkgHpwhD7/DDUQEqA8vL8J5B
nfdkaPsdAXOFHw+IqCCCGKbWc+nUS3LGf+CkrWCOYJRZ1OGMgZpn7TFTo09jT60DoKvljf0myTFO
tDyr+MD40m1evAfDuGOtRt91pCwefej7wjEWBNkyqmkh0bHqv8+hQoTgE/vmlw3JNjxNbtbOWRJr
b8uVcsYq1dgoWEr7GtwjhVYIHeyqSkI6d6Jv5w0wo2sc6qWhnWuUT4Pu7mN3gEfYs4PbuBI2tiT0
8uHnYVICyC1Um578oF2li/fO3v+uBYMZ7TJOxhhtILAGyBwsA9fQTLgxFwND1zE2nVLqZRndU6IQ
QrzJ/43fFw4C1WlzD2now+oGggk1LBmiLh1g15dKpeTX0A9azgMIzWgh6iIIbHOv/j+RYhy5t7Wi
dxTgwb9ruOWI4qXj8HvIiP3vrBP3R3+7C0iNrzdxYrQySk1FG1ZbVqEZdH7qN3G/meMreEAZj/z3
ItHU+RDVhBuF2ooczR5Cpqxqy7mm3AiD/Tqha1pAGOK9pCuTPY/62AfobO0p9m8giHRflhhnMyIu
vC09+XVzsL+abQYH73VSqyIWsUX8SXtz7FpdsWVV5iiv8vqzhrUju50vWyttOKyK5XtuuXy74P+a
tdSPWAtkg139LZSo1XSBn5jICx2HmcfPZMZVcyL1YPW5rDQ8wD6mBQAwiyq5/vO6Fm0orSAlqtJ0
ortmzAHsz+4QEQPI+WB9qQLmgUIKvfwXqcv+ENHxOdjVCUBa28eVzzLnsVB17ak0FlG/d11wzuJb
ZBu3RhMLNzZBtNPY/S3rjO0lW4XisRgEDGYiha+gZRbdgq9C7YQhEL9JBDN5q85M0A34OM8Q5Nfh
w87wbXHHIssxeq7jik2f3QLDtR4btX/9T7Uo76a7ohrUyHQpMgJSgb1/0ffV+tYQElMbFIi28ENB
+pENvOBMx9B/eQBKAvjrxte4fK9IXEgxDSzfK7RnhXfptQ/FCFEOu9Gq8H9Rli2rZhhPVC94YOBK
u3vGfibKAF2PibwYcGxNRpW8k9S9wTfBQmIg5vf+wpfrHG7GJebJVe7SWz+dz6Do4ahZfUDhgMEK
If+ZxZX+Ne3iYqyTCHWRCwPaykBlSYoj7GK6jVLwoYCs8Sp9o0C1bYEuS7aSLpH9mxWv6VFO4tTY
GFMb8q+IyYM0zXU00T74SgQha3ksepw3Tn/EzEmmQtJYw+o1TBAqfHXRsR0lOhR3sMJ+KHB1h2CI
dQdw0apximiwYBmGqOvJTAvZ+M3r0C9rpZi071e6kMvaQNzlt1ExxVwLMG/1lTYBm1EVRb+8FpUo
q1RGYOy/DEQrVzkNSaWclCv6TTuPvZIhUjf4DZdIrX8MniMy77Ylxh7aYOtCC7fRUU9XHSXTzdMN
JCs1wgy0zyuXJb987v8ffoP7ZM/CjTeUHZvg52tWT+DYz5Fsu4lhcjFyVv9yukMle7VS8WzccYfk
DzuXmDcKtbWWUCLhiAdME6yhjQ5bHqef+lJG5GvDkYRZrWFC2ILdTlFXkRfSCNerKWbm2++KGMTJ
n+6Vj9Dnt0R8DrfN0390g7MOHfatPC5Ge5HJc8xtWS2UDLHMCg/gfmJyUtB1NzunEhCemulnXqt6
2gw002l1dyxIY2KACAowBe83ch9D7S33DasXu+xFosdAfe5SpQFO8bV4KI0rFWOoZI5Dbn8bxRrr
3o/XAqD11H0avd1U8qHW0B7n9t5Y1RIvohAKqTRZF/ioVZHgINADkewUuvEh8/bslwqXZxKgHhID
Y0+jB09+cWXRyPo5Do772/4j14hwY31RMcJmgBbLOASF0hOK5/U1Or8CM4dndWkIsbEqPyLemAea
UGZJxXf90dswpSIfRpwh3UgOepoQpkGPC5NlODFVvIHfEpHFAb5LCnlmJ8fBRPsz0ynTxd++Fonh
7z+jeLO8KcmG4E7yiZEz1n7cWDxDaegAqnMyV9TAe8OKyICrrfPHML2Lyx13KRNYZRWUcnqIiSmC
xCWGzItx24b8zvsHhy68cXQccaR4X8xJgAJkQ8BKXqhaMARJtCARoWMGi/l6EmZLSPUd5BAYNWel
LWVg54Zo+VIUSgWVH4iORhLMMhpR2owpNWGqYPdc1ir+QgdHDLpzq8pbhXTcLPzkDS0ACxPMhFqF
r8IcDdFH1AuEnO8atFthvYrULxyG+d4JxTDATHA8XIiiWcjlSqZlL1yoU8kLYa/ULEMqKW7tIQLu
nxYBJXfgHr2KRyntJK6NNseX+1Rtn9KyY0V9MUCBbeZaOxPUFJ5SMo0qgt6uOSXKlZVOsceo20/2
+MDhOz83JMCF57r0ii58NGjqufS8TM5t1go3Jk6zi3hb8p210P4S2EbOOp1rKVSWGge+OwUxeJu0
3WYiktV8HNwVDMcZG9jpxo9K+2P/JOyhErnBqk42fIh99SDhv/Ae3QjFanbOh1I7lDgUVR4Z9Kni
otzq/7ZjqHkYy3OHGURu4XWUkUypkScayZhKCZm+nWY/JLk5xagO3LFbvbhX2cbU6L6l7yvaUtaJ
JRHVZaoBnrQy4FeynbhAAGqzcpzaf/BhbCEjv75nEloLaIEnTetJmXnVtHFzijPYz6RSX6n3B1ZG
RkhzWw+3puu/mqu80CU3Rc1aJZvw7NjmWjJZdqvKY0A52n2hNeWJKMmCfF2B9ZnhDTSSibkia50m
IO8DqbPMZNIBLmI1OQFKfA0KZWTPPvKIIIJ6moM1oxlW4TqUa2rkdIcifESQT9BB/anlmB+oQO9c
gSwEVvPhOMrFnWWM9eyCn4Jo7t0SHGiDKxAYvS9UpJBEn6jhBrn9Tlf0aqiTDc2QE5HKMRtNZUXE
oCYkfw3GxzCa1RUTbDrXgggaXOPhwpnqsIxZgqp5T0SBt5iRLnroI+ZHthmwc0l/2eh6cPjsrw7B
F3aQZYFOhUQ0Me8Imb5viBP3S8qGLHv2bosD6A15bQKFELbqF/F+TvBSKBXiZkoNXBavxktN1llN
7BjSJtYkF/h32rLGZgSny/eJ6IJRPnXz+32+J8tlD4Y3SgenAcs+4VD4HzRax9Fifbc64DpxoPaM
iS3bOMZxHpLuclnQI1oIPe29tBMn6cr+DUvXrIgjHAp2r5O1fEsY3Fn8nxRkZ/JklziC3tjqI++6
9u5gFkPrcPrnSMTuUkjoK0fNk0yvlMFkCnD6ECZZG7CSyMyIlihwZBSLAzE6SBsVPGnFRtZu5mDO
i2utvJUykK57Mw9xIrgoaUd8Dg7sHfMqxxmAHvpPZZ2ZnwkpJtolodCX4/cxkOp8ZejOxy3Bj+fZ
qEA5ghnJuzqp78fj9Z52tcC5w3RU1Yb3Gry1o5w1mZR//MyikjL7b/5d4K8s6RAKJnwBJprv2cMb
PvB4z7nEixqUm0GpAQG5oip4CfiavQgYcLqifl48brtW8CVUUpoqRYqj81NX9hDDZZVjQ+tfF7bL
gxS8XugdT4fJyzVKwsNsUxicEpXuKjWD5HQXh0qM1oS3jQ8ePKZL9oTUZpY8cAarAfPCmGoIxzUx
6B/k6fW+zNq2gyuykjn8ldGvrZm75N377dSWia9BgZHIB5NyEeGvdMuyyEyOBbfvf5GQ9NFReYR6
7y2V2Rc4xPb4uOtGa02IN3igSUhpI8DD3sTJtLsrXIfWI0hsff0coA8lHSi8FR4VkDlxgKJWEm5c
vpHTRV0IiKLvrAo3xcTgPYRZWUSXPfweTmj2KGY7rJGLRiTtsPNQfw883MUcKAp60BC8eZxSfBrZ
pqQ4v7FxfbHB2u3Ko/wzCdtHUZIrtLExzYtoOkvhs2FdF6HZQJwIvKxSo5ggaHmZflUVE5co8uVu
dpRMhepO8KJr2HS5CLzP5akEzUy2jNHv7HxXejopgR+u2Rhzgb3odFCiaiIRrkHn1F+knwdtGMA3
rG6HcPSELOusxJS2aIW5Ai2jmDumWXkJbEz6/rZ0oFJExR+Opfbt3MBUfJPHzzvVE4C4rwpvU9lx
AgNDnefyVKX1cwoR4qF7FUc5v8QNL/+vkHZnWQCVlLRB78GzM83t6nDfRqzys4ZgZJmZaB0Jkkgd
7DYI6d+kqBeFTnDY9+4+14/vksIQPmkdSr23f2pywUJDcjKt09mj5bIpId5o+iT9R1lrFJl6e/Rt
P9pBL/pDKFL/pqqoHP0nvxQcluC8rDrwoPN5V1WqM7EeabHwTsKMX9bgVHd0YCNFo3BNSGT8tbed
231ivyI2AZm2pb4O38Lnk7LZugz4WbJedvh09r+LhJu9CNMVk7e5WogQEflNQ62LlBk+NFuOBYtR
gSzrKcGzTyh41egr4VKbNQRHgctmBF/SX0u1YifKBB8/UJ5aQPcbTe6XF+opz2thqKURhO70Bbhb
E5w3q3rClvP8tEWgYdyJuMZcEG5t6u/qh2fso5HnvDrTeHsWMc0hyJEY8G5wo/E9ZtQwT38NzAQn
4mR4kzQoO52SyPTUpclw8CCrlXhouCgVaQTjUO5JdfyjNW9r2fBkFtkhKA0O9XIqCrzWnKaCFhI+
AwBsvv22pf+uhLHWpZscHdBGcEdwGHCaAGsbp9sW9F/606fDtDNqiLtcPTFZU4aOGQuioNR1a6gl
3fTTqXgThP1+468Tl6IxEyVi8DmWaBTwPwy3dOTrkxMVQu1XDWq8N/DJ+mDUROriTQ/RO8R/yBFW
4NgGnBQRXWa5+gxw/BPfda/Wstw/Sqtdompsz0a/u7ZKl3sc7UfGidZAD7cQv1isp2Ge5Ehw8lRj
ZUQzKjNq4eR1f58zRTLiwnauT9JF+QeckSvNtHKO6gUH15zZCllsPHA81VAVGgv2Oq+sHoBI/8H+
zaWpYiEiwERXDmc8h5/KvOLNjkBtI3J9Yx2Iyu304cj+Cqd0AmTyR8/+YJA/3R1WkdTrGbmCTMda
g3ymlAP0Oqza0MFwzgp/E77sM+7VCej/fjDSlaFzH0y5uJmsr1ijam1zkdFTvP/swHenTXIKtxwS
O+tYHcBECZRLZjYMCi1Fy+IQjAh49GHA1PQhfbVVyVvLs0VzF3PvZK4916ApvzmvvCsZbOr+Nfnd
UqNH8/RDertvA8VQ6Idva9/l/kxOpS+H5FnVxciQqQHSHj9Kax/cj7PhuzZQsme7o9/0HzWLcs/C
DP4WHh0EVi8tdctMKDSyYG+duoVq5F8TN8tBIEaUdl9ZEbWLWZuWeruEd8+7rHF+CKJ6712xfGfk
HskiVv8ZlbaDJJt6zsnP0aBSEKsDDQoH77Ew4RqJgx9tWrGRptqcanUlHR+Vvfx8s6IIS+cxw5vR
2ZbOgqydMlNakBsWUjKpnLmVo3WKrTqyWvUzTyAxt3yOlKf+Egk8jlWg00fkQEFP7QqE5TfX9mrL
d5FVvWJ9gVJ19LaYhyb6g3CAuGllkjoc3QQQVGgUAhF9i1qQQ3vmhtP2Dv72bNxBWeZNzq6yA6zh
sCVkabXw5221SIhZ0aSGJ7bN8/C4D0waHp0MAt5ZFfaS/LeZJYheGndGq0rFTxn+6xCNAQbzCwRE
8EVJXRaS7cnR4qwbDMXcWRXRErvEgHWUa5YzgX3UB1Dbo6xraFnu0C2nAPR4r1vNoUJvjzD7HzAG
FTT2MgJWAJ98FNEFP4xJtVzOr0LrW/iBQYOzqlLySgD5X8RupuTdfiXTTMsk6hjMnFjGIky9skCH
lcHEeKSviltJ9kaxiB/2NQjsmQotvYuqMSJ7MCkXHCBanyJh9qLZfvslLeM9BdgMCmV6Gz4XFzHh
ljJA5WXn8hOAvEsvQAk8t+3ClA34DlrJS3uKL7t4vOEZe0XJ1wUe4gvCGnKooaT//mIoZu6T6490
17RUcitFoUxZuYIJtT7qgRMqHF6+qabcI/ynw1dLgDGl81btNuBgCmhSzNebBBy+FfdGcJCJlcld
QqnuAr4Pe2VfFLN1zqblHLUNlorfMSCG96owkztLU0sL5nVWNhOipxpPH+eqtQyAHu8sbGB0eH92
NJji4EjLgobY9Tmqxpnh29rSGewSK2/OPbBO/NQ4PmRpzolc02feRxT/rhUwILypWyO3/ku4/z8Z
DfnbJnpUFQ9kzrGWQCqmRknMvff3iQKGPau5dfWHugTxfUULb0ecH7pWaRYxyv/DE7YYbdPj3WW/
3+ED7LfoMWU9tlIimvhuxsM9SVq70s4cym+d+F03My9eV9CYxMfP8TIzuZGZUryxQeaBPuh7sLvP
v3bmFswYLUimz6NijM6Pll3jjvMNAE/0tnXfEJQNuUrN+/EYYQi8S1fe0fx3xKPeLt+Yec445Gf2
oA7NPLNyyn0sewRYpZPI6Ke3Rkuj8oxmeNJ6uUWIy/sHTopGnsHAHeB7feChojg++PweCxgtmL6j
4R6RDYW1Gv03nujtH57xjOWo8zAYOn1sgNwLSCvkxMa4wxMWl5sf9f0D6kiuq6vVSMJ2unB/Na8A
wGPDrvMFbGMCTybTIlwxTiipQ1gBP/VCI2jbK4e7rIFWCNxvC19AV/M9PCWs3Bu2Nmchsni7yPTS
Mwq6WJTYNFPBi/vmwkAMCi5ZYrIG//BhkWU3vYYb+WMckTI8S6p/QUZp0RhLsHtSeu7FemWIlh0l
mFPuiQL19npVVJQ+IUhYIG8GKtim90WDhnpjuE63j7Hs0QZMmAOse0mXbVIfzVIC/ErUyYtpfgy0
4XJZRVdiLGaO/T91HNf6TjtLMNrjqrgAL00I7n6Ab0Jt4B7dDVRhselIYVcYGiREvFUzCgU7oANm
WHNNaXka4em/z+3miwajOUlpHC8dPc/pJilik6g+sfUpCGveYH6nkKqJYbM+KlUk+m9m0eemUbcX
9NH2B1H/mzGJkvuU1Wmv8KtzHGicgtDlCbS5iobFP0muF/lL2GyapdCdRdmykgayM7m79tOmZFwa
c1LCU7oXFBJ4SNG6S/d4lIc1rjg/khF97dSatpcXexIjbxj58acMiJXiVLJW8ZS8ofpelSTZuIIe
qv07kHXt6JEDJaJwgzvsfBeNitDc+P3kONZrQJgsTUEM7Z8cjU8okHgQLvFYLE+7R14uebA9qWPZ
uLzgWR77Tg8NCMj5iEuktPTTkNKnBXpoLdqcgvYlozdF9eBXmmP7++2BrJEs6movH/+O04ySrUOb
7J66Q5yguD8tVRImOFR9W9gMHGg0KadGUXEa2hhUib23Fpe4FX23RnxgHT2lHBqxV2eqTdKazBKB
eeoHTT7gw2u0Ov+rr+PLrA2hik82FdgJcJl6xGAHwnZe5smcs/gDnGj9U/8zxgzeUCsTPM841fsC
Pu3QN+Alr3FPkcfks17HbfYnL4Yc433cUFaFg6dWgiXJHktnfN2wg+GA4Bvq65SufSc/jQUkzwJ6
zw1CwtnFKvrGQmebRbUUsMRcxfG/b0iqmWL6AMjGhZY8moEB835k12ft/LLMB5aHVjNloQVxEm+J
guLNqfuEHJoVq91oNBVRG38BsEa75P+j38JTebvKpp+gRf7dKPu1e0oRXWFNIp6m6e3gSfkM7KFC
0xltIyHIPgDpU3jtNl7JCC00+XeyhIDToEJnjgklN1cSmMOP7UHnHyIrXCoOmOI8KhbPmf44CuEG
5iczyuKegIu4D1QctpxIBAEquDHT12gO+Yn2o5idoKGtgI5elLqEFMsE4z6NS0sU7xx1LFdripeK
lazqKsw2qrbsSnmVhfKGeg+A9KDXRQ8D+bw1joy8JsH8Sn/OM3SvW4htAnAuDAx7A41l1YLDWjfD
TpiqQel4p5gsyrjWnOQiuhlJLvo9hOnz322zpBDvDBQX7Z1igHjXBMlSSI9phw6RgybttkOlMT73
wRO0EQyqZ/m7OXqaKeTEWXymaaUU26xe0bYdXxMO6KZsmbu/DFL+t4XFeyp282cnXvJdkniDRQLR
Vq4H95QRMAmyl9P7wsuf4Nio5MAixY3zIsRQ12jmlPLJoYngvyhRyXhJBjgsLS3muo/MNZhuwJ8+
z6fOE4wKqgCihEyFEN4onrqfsYaQM6dQiOPof+9K13M/hJkQCCAycbX2jm92li91OGNgOnZ8sELF
3DDhrQ2GRpzkclEAnSDl6xrseKXfBwXZEL6K3+VR7jXseDo+2md8ywPb56JNkZByZjIre9XNMkY/
bBFxtt/+tRwZWAOGnrySyQVHPxqxGGanbuf3MvLB+zkQd7/mQLySW3HbzGu+x1v1W9wYVtWdi0Lt
dM3aa92e7xX30yt+LInb8G2w6yhI/VG4IxmVn6IQsPIFmZuBtnFOeIXv3Nd16qJhte92DpR/OLYB
Djd8SooBEKnDvIAkJYqNXMNg22C7Of9aIjf5bONQ7u1K3GvRUcApqdg3MyryWIjk8rCQnUWNmSMs
1+wLca+wL9MES/t+Cnvqcz6hVaANOAnBv5mlatjsdW2XqF59hv/hF3bXjbsWepDMUG8M/yWP6udm
RDSD4+qYpS+nvcHoZL95Z6xMrl95h1IwgKUctgUlhSOxih5GcgfEOuMzPARC8pNlUhGUosr+Om7R
sti21nm1MbjevnBsGgkeFQKU9zp3GDhromgnv0p7WBWyWexv48/rvZMfruY/WwrJCPDJ85uS7Qi7
FEv3LJg27gP9jEurt5C6AjyBWEMFdIxU5mjdiyUiXeWZoj+n7Lhb6rakB5mRRSMgmlSDnTpQLZ/N
lzPlGyeyEmuAE6hbZ2neJGJe7TYQYoHj1i7dYFJ4AvEaXXx3b3/RvGClfD6QJpXh9z1uhORkMwfA
V7VJnrVsyHlQVAYan4FA+BXOT2Di+FfmXMiDmJjgKZZVzr3Bl/NyS3+Gg4nf54RvHADOYlF3xQgQ
Cnrikl4Ww5bw6cd4zy75ze/1yMZtc28vxB3aTwYeZFFhgE2ofT2rC2lYCIVkHNZp3b0a2NDjKKOU
Sr9erNOnNpYo5roPoo3QNd5J83MwFgYALPBvP0M2g0uujNpzHn0zDS167dCRwN0C/n2L00l2l74Y
2825wEzIeSi18y1n1qInalDFLp05EIC6vcXwZibXXS3+v4v8Ee3ihXtSTeeRaJfAZ8gNOoBQy/Zf
IucwMpMxn0DQwgSWpXe2d+HTjOOJ4iEwuVKCVW2AzKqzMh4WutZrlEK6xsvid8KvzIG5wUiptdy4
rWUdwmnGaRQnviAODvqEa+XUzH3V3zQQEgvlzsFQNC1VyRPp1UkSQG08qD+a5SSSPKKfofIsonmb
emMtZDepHFdXST8zuMTlU1gJqNB5/eACU2dIcYoRmmkOq37fPNe3baVKmu6DvhXyfuZylkDXdVIJ
qwRnF7/2xiYs1rvHGPGUCIc+ut5dYYFq8gJz+ftrvREXBUt3jvHQVvHvsi9D1gFKwBCX79twXnNT
6P19D5/+9n7Dmmj9OGwgathdwIB4AfMZjqVH4KV+oQCU3hWr19cfaIcodyr2zPhTvSV5O+HBdKke
QI6xIVWj+sD8MXra/CGr0PzYgFBiSGHzm6Ig4+KgeL1QMFS2++Fb8iOCcXOML2eLMjqaOlEDZOTr
7QDg+T8kFOivLb/Mu/N2YZ7g4kSCYH41MdExdJuJQAzlroUitHB7v57Zj5FeFeG79Ed2ofcykDQ+
VpOa6DmP1ticgSVGPZENnmoWRQI6FZDmp4BSZyUAmho3GYy+3SMU2owdIxWKJldHRlURwO2vI9vQ
XJ9yaT6sJiwe8514Ls+00cHNr7o77h6idzbJeOrtIg9vdl4XoEv5gdZhABt4OXrVAkB6Vge7ZzD7
g0mI6WdjSvw3SnslAlJzXJoYpZcHaiGKLVvfgSUsjqn//YshN4pMorVYA/sSfnEiERORZ2QTp7XR
0D+pHKTMIe2ydeNhSKjyiQvCf2LVrFAeCodsX7Sq42zkIOhZI/sKeVcX0pU0szR6mB8zsIwyaX6F
xXWxMibsc1Av7Z1riOF+0TT/Mwc2Jc6YNFoiXh8AwwE1QFhjPvsfK3rZEEOKCJ4au3zy6NNLthBK
iiCR9MrQw02GjH1zJ/be4+xfffMiMlFM4yWSAiAxL8lCTWGyBTxJyUiaUTjwlhXoYPPmH74A/Fpa
vH3jrFF9Nah6+wMq8KbAt7etjkEjqmSa1/7Z3S1hlsbLDGXRujZt9j4uxG8VJ0BifpMgMprAuDCM
aNQLaa/95vF699XWMhQr9LX5qGvqDO+d6wlm/5j4Q1kVrHt39+o1xgDt8Zjd6Z5U7xDQgmPN+/Tr
1UrMFA/fnQlGsV77qC5W3wpc8vUz99u88Dj4FTLNcu4uE6eF9l7IZtqRxR+ha6ByqQcc4XhiwT1W
aiwtmGTaBaEI8UD5AqrWuHEz1qFV7lMDt+G2+vwciAq093G1h6jcubdEAlR2pchUSVJ4puFRaomn
p7ahGkADs348y6sPfqyiNFUjvdd7ldc7Xi501xJli3YTFyQATo3xL+y2oavTxXN3/uuBoWjDN2+C
5kZB5lDFEOr9oZjbRMGE+dbmvfoOYqfD7PKzSv+nZkr0xIKvtZi98CZ3HzHnyz21g/IQwOW5cdWq
RnMmq3X5gRZk9kdTs4nYHm8oyBm9aWiXvkWl8EeZ36Yxi/A39c1EbgBsJna2p1eamG49cumHxlyi
e3Axhv706NqH+E3/jQqbakCfH7x4MLRsGVjH8uC+PhtTJipCRtOdjepmiwLNMx4ChsEcAdtbORme
xmacbVUL/oUScklMDFrA29SwQt5IP9E49TTggaZlt7fN0ael6k+oLzh0Z5ZuqdEN4r9HaLyg+95a
KxDWnuDNx66sEplI+G+/rhUL1FcwxQ+9HM33oxJAVUoPq/zdjbr6jFiKByK1OaMr6Csh5CWG0Eb/
doWFOC8pfmmq21Mlf3mvsulFLQTCtpvNFbVbuPo2O7ubHrapTzupYN1KCNz4J7jMqzAUaO716Clo
zR3QMg5H9XwrMG5U7dqr2er8p0xQJ8rVk/df98ZjrBRa9M3SJw7anB6L+C+QWIJiU0uv53mwo0w5
mQZqReFPJyAURTWHUTkuIBRbCbuwOihwDGAuzxt2V634K6Sci1WAD4ROfC+WAz39a2NG21adSb4O
gDf1io74WVqMX9r+ohhTURfQf8HiHs2VoRs3PZNJezpPtm5aOj5fLww/hgoEsTG4BDLeDOa+V8Xc
O8hA4nRCTHXMjSqdKeqkvJNZoDNrQUrwa9/ZJIuYJP2UBrKFzEeFFNqDvKqJg2vMrPfaBSViNyak
uKiwBJgLXNtZvq77QkSD9sZUD8fbgLAW19dmnHWb9WmLcRMUV00r1YpLmlNBb1Lagz61hiGgto+w
yjMrbsIQEs7XeqQ8geVW22FRJywWqvPBSyjouyqIFx64S6gwqdStVrNM/eYNFGqTg/BmZeZxKVx4
6mmInW5MAyVLTVnnaUb+AHHMCQfyVs9SEgudTXYtU50PPhgGhyho9qODHu4LAyOb1W0Evecl1rxV
6htGH9Cd9WPPCXDGG3POLzfk4Z5YWOqAI6cPArAJYRpHLbnsv+SuRshPk+u3mg1hRLDf+gaSIILJ
mwTadKxMoYpk7xuDGKt7moLcz6XoTHfnO7ZhnfzWOjsJZyF5f2+25vT8GAE8eIb3yDMHsz87Q6O2
Qj2pu5zG+Igpq2BunsV8r0+oMXrK4BZETyYDq1zRtfrh7ra1UpvixSCCW4WJgSUrpalGdIIf+pFp
IZGxyj7PzNHTRZTprgTKCnom7YP5vMlLeM4Zip/Fby5PdciJMgjnLXCiHxc7jGTnkPpz1VpcpSre
t6Q8TkWCP3ZsYdRWyS9akjIP6LUeaYUnO4i6r1Kp+AWLMT8RU2ksLo7bgvJS4iSpH8eqSUIqu6CX
SMDS1kl8cgmZ0h6NajhPP7uM2UR+NjYzdSXmm2WX5MQQ5OwproF1fMCohY0fcx50hKgA5363K3Zg
QWXMdTTtRUJ8WcsjtB+vok1OBjpzOLL1mvXxB5T5NHqBFD5uIK1rgGvs1iN5QivobwH3DKMgCUmX
tQ3RLODtf1QaYYKhYWjJxNC4yIn5StodPphr5ZLXrA6j62ZWbuq1NNxOp3J6fPg2jqmAcs2Hc2Gf
9aGroVNtPe0l8sD25wxpnDL2I0yWZoWS3F1uKNuMpsEKgYVWVkJEfhpdWVy0/FiHFh2SY7+5b4Y3
igLuXYTe2AuIEpWRTRWYdqfvB5ZsQEhblYT32NUU5xuJ/ovXU43/wKfHAVmQ1CwB/DlhL6KlxARR
8zVHqGkalBGhX1o4G/EJVHx99509J92SKQsMacoiKUFVxpBtJsL1ptU3+e/jQMKOPhm3a2z3OWMQ
Sm5xFl1Aw/xUTnBLnR06fqOO0Os78rlTRON6jh7LCzQD7BFG0+odXRLDEQaNRkt9Kb3231EiTQJI
hNNJ/2Jb8PBlklfno9winu2ZvbBd2ta+nokMBxogfXdlpIIRZRkFjSrwDdoLumzH1Nb12Y6BKSiR
onexmfZvcXkeisVR6PXYNkh7uQs7swtbBnNPoloDRGR3Ver/4Fe3GfNCuR+bvQiU1BtzinKw6Ten
QFQf7zpKmbQTh1Y3b3H/1ZKalJSZ3OA2cCGxBiu3zP9TW2fKFJbdPfTwcUBk9mTigl1YmrM0YfnP
dwsaFosd56wEby4ia9dC0Bx9P2wQsdhCOSfxIjjSEylSSmd+8E8ceaLlo+RljELf0NObiv6EymJ2
6BKo/dSr2zUTaseslsAJe9W/aWgFHQrFVTkbZZmtox5syXM+PaY/7UmQFnq98AcZPRBQ9I5ZdsEb
UTvMH5Tuwx38X9NA521FpgJsEp4fmYMlZqAf2iO2kTTu2/z/8TUAo0zur+X2F8vD5B8J4ExVK+Di
deFV4gDBdgJBCfyAOhbeeY/Enq7MJyL0esXbAfxeEj+AoMnO/L3U3eWnO2V9DtA8AcPq4Jqjzgk9
hsuNHuXX8WX0FueG2Yt5p0PW8DrCD8hYSOQTaMs4Xl5DaG8mRtez0fnTmkbZhYikMA9lABn72CzA
BwxRX8h+l8wbMSA1YcgbemBxL4pXrkkPzyRNkIqt2/Z0OhTe5WUZ0WUKAfz4fOwnx3qE9KXbbqyk
8DyGoZLKcFbgds2KrLvHz92KzvcTt54bHbZz31djR4m0CsHI3LaMu4m5ujyPCv1CqRQbDLyVP5tY
FGyqafIRVSGw44ykI4nt8ocaSK5rq2Lryi6g56q04M8TVeUvi7NKUSYJOXrKBtoLFiCOTvAv2/Pv
REmyv6qrCxHqXoZN/fopWsDW5yEnJ++WrkkwbzcJ3ZtlJ+e3XmnPveXEoP/NLLuzoNRBCqsM5mSg
pbLgesDRs/j4fLdE3CAv35dHe4oNsvuPzVaqCFFq6E8sxdsV+zapR0Do82f1MZ62P30Py3dSdWgQ
Ut8HMQcP1b77Q7Lx/c53ELUiIyLOTe1X0YpVMFofmVUCWHg1RYq5iZUKH4/fH1uaED98X7pbD/Vj
fn4A/XJ4EWh7w+oa92CGwbFClwS0c3TRRIX+r3PmuPg+e/lfIudGKa4hYTBCK0iehsEIwTOCABbJ
OlSIdugvExBtfwZk9mPio7zMdpN4G6ae7beDvMAUWrUG1mePW6MgSOW/3j16AVpOSxcK6ueP3n7W
oyppHU1wOpiFAp2I0/iyFGQNzpBMLI71tjuRq2eShRzyyqTWD2egCSNa+k1fhY3wG3sQqOukk1Xs
jpU5a8vfX99mGiW5PPXDTlR4OHFSrzxAcvCl5lDx/msV6zNBxyA/QLDRgxQ3YUelLK7f+PcKxiW2
gctm8pm6e3pRugA+yLqv+Up+w3eoxY6K/1Et/CvAT+uD8t0bwTaA0/NKj/uRnro62hKan8lrIDdp
YeNDf2LkZqjaVkW+znxSFf+1IAkSGTIXKA+IxW57pkqTo+/yy8kGHIzaxA3cGeeLyeVcN/G7Owh9
XUqp4OZHRrFnNpqlGnThNqwdWCr+7hRUaaEL0N9Ys9UMCFzHedF1nWTN/n0HElq92/AJRK+OQMwj
7F4My1P+L3MolEesfjONQ8df4BHErYocaKWvhxF7Ary7rNS9buhh0u8cxjvJyVQMWFnKftBqr6bf
VAkiFir1kxG9MDWXJroDKMuVvbi1huEy39Qe6kj3usK2W6/BIzvy3kUc8NyJW+0lv2I1mXZvb2wY
VmZTkFM4YfLRuG96lZn5x+wtOWA/wdFIBgjudKnGiyjM8kkAbTE2s2DCCdp/upbgSK0KURh6dfQP
bVce+RQAN1C9CwseuItOtUAfqOvRMJC7NMeG5FXzFEY35glut+I/ZnDKTUAJ4rGCg2X+feQQsqiR
ZS0xkaFaIYMHMdOsROaGoxvIliQv/sIrcP46Mq4IwiPJyaOiWUYKPFp0xS+SpMGYg9YvfZPvaGV8
z2pqnxQWcGkVxRdKp2iLAYeBD0bIYkqpKTHToOX6wkNOFqNuskXts9CEiTNYSWOfrJwhnt54hpP5
f9SVE12nhanQ83dYIieHCfrPk5TIcCFb7aqkb7ZZpLP3wBdr9Ud8Pfa+/tdMkSRKWmAq5XDqccJm
+9jm5tOEQ97riP1/jf1u/EOgpX7c689hRLzmaJezDR/Kxd8L5NK6iEExxFhkXW/BNsq9HqVsy251
D81GYvKS+yDfebpqyXdC8fmDcxnuA18vLFUJII3umJSvXNa46U3dsDFo+DVJ1Pm2ClNt1niS685q
gHflQpw5zC8/JhknJhZczo1dZf1wcPq3Jfa+63ZYc9SDYNsU8h6nWOa18beK0RSfjj1gd4J95uH+
BTKf/1JJsLW2Dkp1SzORZhggU5/E9dVZuUIGKFGfq0CzsPpcaSwsmMDrWfOKWgmy86kSacpaboSb
NtSlaZfeAWimnRtLD9Eezx6yZd8Lf7wwg6YHLvoD1Y6ITCb7FvLyRq6A3IW5YjCuruDgIrHhbxi4
vM2DRm39+NU6FAGWqfce7ZehIOIZgKdTApCMpPUkEoJWfmzO+jQpoAGRSurqpWthA71klgAXXG0a
N86+ssUSLrDe1Ui8UCbsacJVJVXCyxm9j7Dq3WKWCUX7WtEEc1cdIi0v3fTPWwBb4tz1mGhnOMNl
uTv9rcPngcoOznKN9KqsN32sAByzppB7l5urit+HtkV0Kw6OWPt9uP1IdPjxDk6mjiPq5LDzf3Mj
xk7P/5RrJsipmqKU/XlaMhjvpPQgrWZFJ6GZhpySHVVDNyFCCfAn4bXmVBT1DFR1ljIGaakTpCdO
t+Fb0TwKAJoroRG74+xmzkd9+gWxxX33usy8/Q84rzgztMQ80rSz0TxSmvM96QRkA/yI60HA6pCZ
GizqE5zYaBVoZovneywP/ZIf70/iWe3bv7Xu3VDwFONCN4GGoXEMhl4jXSY92Xb4G5GqWXaXmEUX
i+W2ct8UGkvLugAB6qaZ7vyIfat95eXvI0cTzcD95RycQxmA8K7MbkxaUPXV2iLyfZyS34E1o3WE
pHquAJc3vdoRLjdVINuPvZL98cuoo2XXmedy4ow3g2qvBeMvXF9kWhdOTSiPCQvVJu9DumJdsBQq
6z5sxNLu4rWDL771kvMWHgtDs+XX0A7jp+JT3XMYDVg586kxt9qbtP8xOtgplyCEvP3JMUvbj4vi
JQZbjah3py8UZnB5ItXPHkADuG3CN865VX5V7z1oy6GYzCoWPs2nBJvWbaVlDVoEYXteSrgeNtPX
Wk2p8ydErX+ziuTnIuAnw+dc5MY4vPeDCxO55DVCL5Q09K3V3HoCDi6Gk3hXmqWt15yX2SZHD5VB
nvaxA/2B2j+vFHKmgEWZAmoLMiKWKU3A3TDMqoXwVIjwkQWQX0Xiv098E6RHc3k1dQd2e756OTPY
PsVbmUkUl+B3J+OwvZ+wWOGbYu1OATYA+jiET/z5QyQZtVzQyR3CriZqXB90F+EMADrbf5EiMhM3
PyYYmUcnlbVwY5q/5SLri2lW1f49PWjIYzG/8OWzGowoW9gEMrM5zp7gOcJVDAg9fB2wvND6E52Y
JJ/EUkeFHIZ/ym8Xk2cI/rWYkvlMel3Q6WhMvTZz073UE4Rtc+NfttfVAdfIWQiaXdpsJGJ8zpY4
Mdj1KuW5dzsKYrE3X33SOQ+oAL3ll6I3XQb7Seb28NXDIc9ag51BkcLWD0b1aVqEwSAP4SH5qt3/
R2iDodL1wG8GLtybJ+d5YnSDkDP++3FYQajSHCOmjt2kufx+MAC+5muSpIzC6yf8x8TZeRT8q2ZN
UVx1CgRl/Qe7/Gj4rzIaVLdsSYwIqGpFv34SjDkiUQ0j8WyOQDadJ+n694tkfQYXOChKdtiM6xJs
TAlffqt7rqtKTKE6HQQq7euUSfMOsJo9RZEFUOBn2+GFC4Vh1HmUMnKdC3xotFLIqKtzdVgChRBe
4GrI9cTgufmtxAhTi/JJqgmvT1iDmMRQOmPI7jpqS8Ft/OL4sEpDHWR7lRpOsbSzY+E9bXnA97iN
vUjLjVKq6HKVde/+aHkFyJua6Rra8icSrnsHN0ucUqbTl7lxsEA3vo31eo2o3j+wQp2aPen7sMwK
qzCja6ix0Z7k19EeifSoJgAUVNvLEdz0v1IRkyTDFfIagTrtaWjcjSkyZXkWEndFV7jjHBVVUwr5
XAzVQwS1JNx6Np9RBiYuHFi/KRw7zTnaIN2kVbDoqWqYB3dB/6rt7+Y8AcifAuo8k/d1n+993GVF
p+Dg6u4CrG2UbbwrkeqqTnpGYpaCGIe/qryToiQd0bW5100GInvtjTt550byXPs3ecvd7+3WDhgE
jceJRTPKAYsm2vxurn1eq6ZeuP85cAuCUxvUMwiWVJAC1PDaQOBNuSG/ZX7tw8H5UOB79vYuE/qi
m75nSNOPbvov2F/THDUraJKtGZel1XajcxGHYqmv1tZ5gtFLBvek8FSXnkiWkDSn0h4d6RO6SpVt
qv6fXNQxQhoPkQKbWCzZu1unk9GBJ8Z8DCx8Bppi+rwc4gLGOU0TCk3q7AjEP9Llp6Qi7GegNPCI
xHo+w5CsFwkj/EixKNsJLQPIhPbAHx7Bf/H8icP0jyON0T/VFp8c8+1HJEjMO7njrcG852RfNKK/
P/pb57QK7Wt33PskLGmj5l524A2jWR5FgQN2opF85szentYTUvDVUedMt++C81haXP3BYr0FYxdj
UkNd//F1P76nDHGG48AY2FE1qH8eUdnP/8avYoHEiG1d9nrLWYl3Pk21Xqvf3vqfJp6qXjW/vOH9
deQrVwUNL+6ELUNmlynd1/elcME9piumZV8ntCW74hHtWZGasRziMGv7Mlaui6r5cQh3tlPRec/t
oADN5i/suYKTrkKC4CcCVZv5c8g4FEfIyvwUgKq40pTUil+D6HqkGRUy0W/ajmG0TswcOippnpjF
QGxE4uGAQ6x8yO3P7R2W+vIcm1uqe04YY7vLznlETz3nBRBkl7W6DXROJvgUBd+Biteep/QTpei2
5eMn+74xu88ojpX2mVSFC9fSBId0VLo6xPSgl6CdeAgdeygONt40/coRSLXNBYAgg9W8pZdGIf+9
ng9q8NHU0VBs3Ld5SBaS2cPgy40GyeIP3OOsXIG8AXju7O/oFf/rOJaxBw3zE/cGNGjLTahqmBJW
QEvp2L02CtiIvy/xrc1lRMO8Ac87vyTxO+9PY+8nnL1Kp40D1ibnIu1CwXXj+PieNwzREhbay/eu
LHApJ/qTYjfimeorJBGCTVB/UwIX/fckP4oxMMiZTVFiywr1j++Bo/KVTqbtGOfBj8spvQwhwx9r
3vqvWvG2glzoOM3+nj1l9y35wiMImiMh5bqcOh8I4fKk8cmlRGpp6yy4tCFAwzbLjJOVAgmsUxhM
kr6G8ppTa6VM4nECQnCl80pcngwtC25XU4HIOA8Ty0Ec5zEVLwwoFJ2Hfs0HAGx07NApIUI4Hmxs
htnsi/MO8gznP+N07kMg5YYMhI3u1Y+1FIT72UMojh02zqn7CQLBssoSBkYxambQ+7AaujloQWH7
Gb/bOXyVQdeRSmRgyyAHFxKr+RXSSKzUq7d4KZdAALDjqSJphMB81kA1Aw1ssf9J70hUoP75cSDm
h2g3KU7Wb0DBiHGLBswe071rcbQdDpYmsx8XOmXDfTZPHDFDqFfD7KDgg3nUYbWBQufCMKhTJgA5
qOziyxWWT1SsKfnXCOZ4bQL1cU63k/+5/uWqskcwreL7AtKKEAFOTp91DvjtllCMebY74+iku16r
Gm3c3rCbNcvtGO+ojG4bf4A9eruL3vwgQQa647QXL/8D3lEEhHRadEv9PAvD2HWow2B3ITH1fSD7
Yg0nhNkLwREt/YTPCsMXHRswT7uMNlnnwDz9vYuzSpmmryN8FbV7/UzsQ58XE8mPq6483jdxUQOB
jfPe/6VdTyBCtXPWOu06LyVi3RCaI2RpBNSAazZ+kkERYmC0KiwO7l9CRlaMaLwGFXLHqA9//3Id
CIuP9wzet6MgBXEhka1QWm8MTHC28tI5wJbPuZn/iTeQUydNl2cMFhWPrI1UOiZqL1XoDrcGWE4O
FTqzdAB9bPikdLr80MOaejoKZ3vPABSPhPxWqr/5bndvd+HclZ3EdqFG1PcwBS+FtikHw9q+5Ofl
i1P4f4x+ZMLZek62TnsZR5VWyopOvocSq5vIza3GswhnJ75yLVuK9bOwHSjy95m481UFvcjCN+1p
0poalY9VAIEgvNINJPifWoxu5KVL35qLxRyZnI99d4afwGyp0GWdU3py9hgb5rGzq+2h1jJvewRs
Hr1ZQmxExRWxLRBlTNLMKW9gHyVHhtdRr8JCwSDMW9piC/5og8XupnIoYy7Vv2QvFqVZdqPemeID
tj/j9mmSOluqbIIMv/pBAqIbYAE00cxrja07mV0SmJwbRo0fYZ1Rw/5bQ20f3gjixepPTESezuZ6
swX1aukzmxR+G2Yw8s6heMbkrNPrf2oFScZYxEIomZq3pJIw08vjMNW15ElE0FATTvKIXnkIwkYu
1Q2zo8afrPkQD28QTkpETo8q9z+H4wn4i0Qf+7Ni342iy8DCNeC4H1W2J6+JEvmbR9XUKj84rHkr
d6dxu0n6+iLKMybBxq1FlEC+Bb8iwwwdePjvFIv588R3shRev6VuwUM6j4PwtIO64bS9P4LrS2ND
eCvClAm4HTFIMD+eaAi9I7X6ezSwgy2Shuos6IUW+7WN3BV+RH8IW19BodxLEXf+hMyaESSN/I5s
axEiX/hgauTlOtetzE1Ls0kvmPwYHNaSBcFQATPtBXqvxF8Zshz8OQfHein4RHCeh/mRkmfpR0J6
6+aA/027AnrCqGN3ROajmjaybXE6jCx46ckBtKHNMjQIJ2xnFzn1xezYN8GgGCdOG1VL/oTsr33J
papeLFzBTsJoIHmjuG3gkvMkYZ4ItjFEtInu22eJy6o7fNyzkGvrBOflEkxHuoi7Yr4RfY1wusOS
yaYsLOUScp6VeNJtpuJzHlFGujdJp0X4vDfvYx2ym2lzWWfsLyzHL+hPg8xN7j5wAjVoGIsX5WHE
0zMWksOvba8W3c9JuP/4q2oJObHbrf0MSZA+Dbley3wizVmSPIlMSjZ3M53EGPL216HNy+T/QGTi
xSBWUQiL2OfY7gNBhD2lTjN2GZrdJnV9WQbrAjnkiO4mdga1OgLh3Um8QNgOhe3ulg4ctjzKL8Ij
LdMef4LL7/Q8KtsUeiXridXMHBPynMdcFCXpS3BOhCwBCQSfMm9Ru4gkdtstP4BvEaSqj8tLrE/j
x7jbf/1Jp75MsIfxRFaIcA6idE47Ng+QX/Aq1tzccAnOtfZibGoYG669Jvlt+d4xI7uVXO5p+YoY
Tjgcl3OC/ONHm4ibgJX+rlz81HZIky/QeA+3554QeHUzToqJoGk70gMinyMhBhLreKRQAOn5gpRv
PYgNTxIv3ntvyGVZEQGIY/FFJIokPLL7sm54w9u3w8Pvl2NJ6BC4uNcQ2RZnsUowxBLuXX07ClvH
seZPfArJwPy9pIm5qgw6xZQDvRHINNL4YXtUunRkevwD0tHHnLwPH7hQLBwjNtWYBOAgexdiNCcf
7bI2raiMsjiCHD4KoSODovVqruBF3FP/kwABWsX/DfFpowt9ILW3wXbV7n8BC6RH8liPNvn9RkdX
nAayAukKil+eby/deBru+MaDY1tsBRWXkwYq2sfXIvvn2kQ3GT7x3HrgdC+6mV5fx23UJKSQpkQE
hGK+3n5ItngiBkaDuzZgXVTlbL9IALW/mxg2mjiUnpRLLaD8xRvYcJBmoZ20MBKSOGiE0TwbpQKQ
vBKOTpDX9PAH+KnsG6BDx0EH311d/T2rs71SZhVbHj1drvHfmOcrfAgOMSeKlvBKchcNnsWzM5xj
c+IYU57aKzfrKTRcSsJM2cx+I2wijEkX8P1oRr3hkme8FNOu+Ko3/2mrv35rhJbtrZmPhQ2bFw4e
auBPPOmrSLQA0sef/BP6tG7Z9oNDpR0DSjvBTk0IwM6Xn7Vki976AFP+i+6xhz4QgORMMv2yNCMb
Lkc/zoViAdZG1aqc9oWpOZzLNyCIUj8WfnrwvI6jeXicWl1O6yEm+VTfBp79SV3qYTfF2mdB56gk
MbIszyTvK95Uze6U/aTCkAfoIWkKBQ9FSeRhgG8WIHqKnyxIasBFAY3PKBEkCL2S0tEiv3GGqbGV
9Z03RK+Oxx4ck/JeSWGWT1nf7nR7+K9nfC84hFEHP9qUgi5yeQ9CWNgxbw8McQa3Cu6jeMbU+1xl
7rKT/VGrCK2unlElY/0x+zWpI2WGxuq4LCsuZNNKfAZkgquiwL9knk4FIgLoIoGVkN3+0xpSjWIW
tLcBvXjZbbY+l1aaYqYUQpoI/5oZuE3SbLtXhZjdIe+EcPvZ4aFD6t7BL5PRDoaD/nzqHCPfoKOC
bGrxKpf2laTATXkmciSrapoP/3jN989lJw9jIXmbpW/fhUo7T4MpZ9yzD9jl2OJbapi8016IzDnT
/J2LKqcKFo77spEYX1Y58RBtdy94Q3XqscJlWHny3DaU8Ws5stwKIjCED0bj0fsQZWuxTcl2VR6w
0wWwQbrfnqAohqCairUrg+FvY9IGiQHJn4qF/PWYZrZ6EV+/jYXpkF9/Ph+8sHdWmBhWt6PRPtIf
YkVqfz2720kt3CXk2WSBDyZCil6TYH11sGJnSlJQkt8ot7Q9niXJYmE0GBfwHEHp1+ZZ/FxLUbUG
J87ohkQ5Q+lbBWYLsEmFecOVrVKahk+0CSIL3pa2uUmqEGC/gF7eXevJQ7henuJjyTtgWSxKLhOj
9nTfF5knHK37rWP5ESQ1mKzzjhFlOU80euF3AdwZ0OlB/sFF87jeMwp50ShXMfjAQP86x0BogicO
hc7icRXzVhFPAFWFGf9aEgcBjpEKjKmaD6Ko+c/A/1w5ZwUipZLB5o8BYfwpfSzpy65JxpHrRzIH
5gJdgl7PGeDt5N8d1Hu5QGbueoyZYiGDDDw+T6y03IOVgouEw+nWptVX67nR4q1L6nujBeCsL3lA
2DQilSIlY4hrCkVqaZJnjaPWrPoEtG6MC9LPjxIb/iQapkuPSD4NEfzR2KEnpTpb8huWtzxBsWWg
PH2N95Yq2jrMsbe0g1arpggniJkITKVhqhxUanc9B34IiuoQhZP/BXOGGHkhGBNnPWbwNTOYJFvy
XiTLQ8bXCE0BKUoBz1Xytyehz45dTiIzAMs3+EmCkhNv7mhY2HaRy4zeR8qgRAjpw45Lyx0rOZyc
mBrwt+8j5TLaAm/n7da8O0PzMWeNn9TpuT1r27fy88Yh/eUOlJHyaqwFB5zpuF3+ENyASUeJWFSd
SiYFEw3W91ycrGHR8MsHzZcN8gq6Itq6WAz/Cp+ALhO1QEkVwaWkHdffjy1zQcwCzQECIvGc7k4m
Q/au3sn1dpgKhvzNP3Pynzb35W/vZCZ51CpR2r8vmza2W5o3FOYCnbvogwCViRodnid07ss4Kkxn
OX4OhUsrbBcdcm8SiQzbkSXJBi7+H7BmJRDXoMiByptJEsUGXQxtGvc2dXKOWPG6U+nudOjS5Dbd
RIUzKIS7zlirNbzVmuM/yEFRz92bVtgJuImL/Y2gQEcxrdQ1CnEp57NrJRFYRtwKMo4UjWR56eX+
M4XPhrfDwajwKyKl0RYyeCl5K2eSjQWl47bAISxpx54rbLAt33aUK9Fwq2Q07OklxN2UaLCq90XJ
M0yfDFlB2pgGs31yAOpXHV+JlN/oMNqXnsXnXAUVCZ5vD8f1l8VGg55Uy5JQGlgSLHVd0ehpj2W7
C824XzYb9VEdB5s8bctX7TIJXi3OfTaWi4NeKaHT05Y5+gdJ3ibzGkz6yXm2gW7oYc0stJN7Cuyj
OC/BAmBpS+5qTyMUWOU/2/pvL6Uihp2Gx6NuFb2I8nBFX5uz9hcVgQAmo0XAThnTcKzNrEh3p1lO
2mLS+Tmi0zUTQ4eFmVXWrHuUn8HumbCjidIcX7Q50vMtbm9hR3zA/sWyGX3o5eRxCFksiO5zx8XB
GLkp22giiqVeOuObz7mPJPdyxB8jbiAQlsdNLuN1PyIJgZJy/gSNBROaamkWdJZak5XkVrrUB4xx
URRk2ZUykxDatDBsyLpY6KeYTmFkkZ+kqAjNdNcD5AFxes2m98gaC+7zx8p+VlU41m+bErh0iUTt
4JoR4akZQCs26pD6idOSQQwIdGjZPiaEkOAAWcr0ZP0b5mP7s+xn+ZMLxXNql8i/oz1TKGAKCr0P
+dIdTOKHOQBWT0+NMLlUN6+o+XUv/bAaeXkAqUZnW97/c2Sw213RWzSwS5iR9iAxY1wPluDJaryA
Qkb2j6JfzwBnFKia3VAGBOsF+v2HKWIDigtvY4lG3JpeMLQ4oW19jUoAOnhGFbdFh1BMM2gdLdy/
4wbrYmuktCAqeiyBkdVeK7iRmKPD+kPS8ED4/Gx3aSssl0qcHeNcXNm5FjtU92OhspGmI201lcba
pnGMJNJjUcoYPdNZDd6158GjTxQYpS24Lgk37jZouZkkJQI2gtWSUlU9RsP6H3znMA7wZRWiTlPt
W19gcTpCVTXR6f/WENJORufs/GqsZVvrE+YpD+4ja04gFXw4akmpi4opRnvg+ry7aF9yCNS2B+KM
AThSYqI8a4N7qP6C1VqNhUrrdOTN1GU7Iy7cX786TShP4d9E0WmySfF/oU93GbFIGN5YHcp1lEN2
ldhIFvVOjOvTLnmoFM4BQwE55YZ1cf48xgkVgg/9mNOOvufky8wyN5IGAdK3Us0RWyZhVuEpHRdw
w0Xm8eHcNL6RECyw6SNcmM/RpdCLXL11oAvykEndYz9mMuH5GGHO0E48hQnu1VcNm5OhHvPRbkIg
HHydsxBWFrI5NCcCXPaNoFrWalkH40scUM52uoUs96BuU2Y8nb3A2EkwI/P08zlZMCEzkPToUiDL
P+dMeNgaXJGSEBcfN9ly4waNA09JpKMP/gi/EAWM9CeOMXaWKufKcU/UK5rAXY4bPjU19pqgvOmq
045QgsJTw7DfUZyhtoQAjysds4coSR0ngd3g/ZLeivLORYhK6TshteSIqai+cp+sfdqYNUF3/J6Z
AmzZpl1zQ69TZGa23vnv0jSvEF8D8nLiEo5Kcek9VV/8fCUtqhR3QzmF2RcMyGcn9/h43p56KKhN
QjhX0kXaO2vBDDX+Yosy4rVKFa48exOmSSPmRDtG0GVI3oOlFQIQjkflS5y+fTYUK2Xdl8Xk0aiQ
Y8e7Tes5taoYYU+vKGJU0atfiB90QA44G7kofNJ8Cvnf2mHBkcR9AJWKiw9x4oeTaMC/dvfKZVcn
559ONEOJzwDVOipes3BOXg+ZaIXBjzadtaJ3mu86obFLnG2FWbnQk/vjJes3FRjPrqKZzWwRc3G9
BcJ6l9FyFG2GA3KMKIK/utWf8Sxv8UHF+cUgDymu5S21ROBi4iudmkhQsdqgEkUwi186g90Rpx4S
95gsHDg+TddLIJWdtCxy3CBfBk5qjJcMnZRHByfXNNPel3hONZ649xTxrqCgJ1hs5mYOfBuTrRTt
cJJf5ie5XnHIki11bzCRYsN1AlEDo3LajvAC8keqbcpg1ZRnEOKSdnUo1dyNxhDY6B8xep9ZnTz0
R+3UrVHH8WcpcsCbBjzVzse9YjLT6MjvreFWUHaLGCth9YidTCzCuZMVHSSSJfZCVLy93qcsMGxk
FsQNRmrOhtrKfyj0ZpuUMErOWmPxtuejEi1f0F2H9eVXL9UAmP19izMqs8YFwZYQBE23adIll0Fe
ai2t5J4ALSVMIsr516skX2/9RJ77cndTH5UMHqnBkWAcKIePWKjL8u13EkYf47D3OIImAH2Cwd3H
uK2WCZj0Gae2y2G0KM9rWAvreAffWFDh3zi9HtkM6A4v2ODxgBuFxmAUbs93F9aI2PxrdV7INViR
D5QMdpiKkMAUZ9bjSJ9I949GO51jUA+bIqof0zSIfx3/mJKmwUOO3bIwsVkkdYrWsOhmkEUmvPV6
/krSvCo/BSRXpYuga3lTgXJRFR4sWfAxsgyGlE5OwnekJJMQwyJzxXMeGqeH9go+x171z6gqLn2M
DleVufjq9AWUWhpkhMAbtazt4M+r4SXd/FP1qvGBwMutaKBaECM4EOXtEoAVYL+/E3LESkCofczu
VXGVvLswVd1RFBlR63IgORKu/yXxQjb64eI9ykpWkUMYVuqm4Ya1WL7UYJIlUndjn6ITifFMfJkX
ducdMCatDoNHgW/ZKx018W3JVm0Z/JcX9c/nqNT35LSJRQVVx9qUF76rx5ODRi1/HUa0oL+ufmg1
AeSOnxkoruiQ7OUuLAL40AFRWBmcIGJvun0h0YigfTguKNxe6TOwskNydhXUQueCHBulMV1OPD0h
eiyJbPb2DOKkIjryQi4AZ9rn2s59hmiQIey43Hzb9kG9R4suA0BT2LeiW3gfdFI/oR0m2QMey4cS
g4k+RsQxCbcW7ncsAGgefi1kvbAsFQxVXlk48sE4P7flqDgF1C4xWduQSEFr3A3t7Ao16TqREO3Q
wjLjkfANjrQBLhSDbKCCdunICP35NAhPGTkpvTbSqu0bkSkYqeHUeReRBNATxD/zusDVJNTUmea6
xf+z/VD5pGWvs2+6ZoNg7BdbcNzj3aBz6F/Uxea9Y0lHoudsNzLsnCHuZOoxm2WuaQ8j6wqmC1N+
dqpw7zV3bhZWDEDVdA7xURDlTKsix3VQMO4FKUIo6mstmDHppaYkXu6jaW+ePWfryqjoo4GsAfRf
yt4UQHnewb0DFM2CL8CAhkjBu0EWyIuJJNUge+rtsc8sLk6kPUVlhZQLl9nT+TNaGpjFF4IiWD7L
WyNH7sgNVJ3NQexGli2ioiuQju/X46YdSvna6EzmuRbOVcoXNzyVLs2yKbB7GsNBf5jAaisbkTyN
ljUJEGiAWQ//gdqR1vE16FWXQRmGrfJiZ3+e3AzM2OyjkPvh1+1eEj/XgtBxQ0Xm7Rb6K1xZNTbJ
QnlniAXHnrRURVeksXLJHH4kgBOCc8uJS1riAVK7WcTs0BzoSBHSnNvDlOIXmCmRVSQKp2vYdRFi
q0EWLk4fz+BJ/kI/Zhjot9jNwfJWtz6DlNm86BkriKmt0E/KgnextjgYMMYDQbR0vP73EuvGaYNF
iWcRU2/6PBcJPXnS4JbKqE8Nyh7rBLP0RqWXK+zeFocYP0EyVXJA2R7HoDIbsQQc6KcTGdLMqwCB
13g4lYxCe6Aawfo2+ExuHm6E7AYcUpu6Mzo5qLFVSuvWHOB18AGdiTx+1IwPWa8cuR3P3hShj94A
uyJxQJNPGL7C54ke1326M26D3ecZuUG8R0SKHQevmynZBRxgmmOnzR4suwHu01n/IjXEsfmAxfWn
9UDNEqAO0hRtW+tBnoSJb7O5FwtfIJH8cxRPAKN772loewyVdE2xChw7/CeeK++Ls3Hpgbcpfm+t
XecEOm+b+R49DsF1fL1m7Exze1bDCiGwX+Px8bm4XcENDAuVAHeq+8bzqOBFIaWgXjuZ9cx1Zq5b
yiNSMg73wCpDS+TG9kZLTESvCPw9VxTzTKyUwcxNs8dW/Ze0F9U3dswRx7JFZvFBmcvtAvQxjE3K
rhBhWnOHLhfroKIS0g7bhdcj2wYG2WyfyG42dBABepO6d7TVCyzxxEhmacDsAINz7q/uzgGntbEI
ExxtSJieqmRHu/LYX7Pz04zWcNwpGoYjLIlrBfDE8zFb3uNKCoJbEKtdqD9VN/UNkLu3Yww+8lqh
uXbqjJXRq6K+NhkCEWTMAdAF4N4aucI55KefJIa+1thXmdOS01m1A65+MrTo2DPEFHt2rgyLDSK1
9vu+BHOEMnOF8Vn0rmWwcARwDsrK/GpU2xY2rP0bC/yAQb3fQSJysdsR+a42mX2HzU1GKgvpvU+O
0XyavwkkC9I3xy0arvpCDWaXjCmjNe/iKGcyjF/qOjyn4yWJvWzz+mgystNfng/8vfWstftGq6WP
HaqvPUXle9UhMWO1Zx06VqmMdvQPSrvnH71c99/MziGKIFvy6NYDCoh32u2ztSyKjI98MTFAJSBr
JY3Ule6HvvpqThTtm57aPf8mbBxvCQL0RO+7PyYROXfVdyiHfcHIR54XgxSOS5G1t/nHFYsYLWpX
O+4CoLPoC7MTVY8GlPPZRxJQzYWBz2FsxeankgyMOzG+Fry3IsM99SjSc9mfm052jX4tBlDl20DR
uC0Z1/Zj5b6fBhTxpGm1vIm0hHRBzrSsUHB7U7NexVYVnpg9/OLFFCkF1AO9XPhmWlq+qRJSCP/2
MmSt4iYXFGKDc78EwEbPI99ynPxc0QpCGp22Yczm7A/h2mGBstf30RjpLKz7uEuiamAcavwm7v3V
7cWY+9UFu/V5kb/gA4ot/MdZiMfj6TSgGP2IJF0QfGnzmKEeGSZoo+NBzNG+sGySXXTXwgMUsiXv
8YHk+ckmOmUSjRiqBoxJZdkmh62qsijwqE5/7A7MfnK9nAY0MMl5T05RLfC87wauIrTyM6KqbvT8
7utNwGYzVcczjxky2GFTiBuORAJ7eXuHU+91/qn6FCPbRyziX6jtyJiBM8ULA+JtH2j5zsp38ZBG
kGbDYU/eUtEIkTqiBR2mMWSaNuAsRgUCERnN8s8NdNKw2cOmCFiwdeFSGWrSj7l1t6mCkP+qIaWc
10zIgzNpE6+8W4xk2k0t5qiHYFyNXTE2m3gwz9wUu1Jck7F8qHQL0g82U7u0ZAQ37B5Ln11NNKae
+vF8exa4vx1bmrxwGNpoW/jFJY5yVeke3dFpts8R66bJcrsFgltLLzpWcWTkTjxl0EFMw61CO3YS
4vPNWWyOXbXm4dBZ6OLge8tjkDPjqQfwbcUY3sSNrDbRlwUka+ImTOriwr/RGrSafd0vzhA4ro3E
FhbMFWa26c7toIyyxEc/vzb226NEz6M3XseePIr/5E/VR4QkMbKyTIbKWFV1L0MPXMtJaBdPNEKW
ZrE7B9pfLX38HhM2Mp5YhVj1V/x/GqKCXKCEwKCp2O6vzttuR7OPSy3gC8gn8tHdy8N+Bu/e1vtN
RwyDMswLeg5tM0QrFdougMhmgck61xo14TTXF+DRRs+zL6hwu5BE4rJ5ElHBu3pgVtOT5VUjS1Kt
gsjvg5wrKpgDwD4lGhy7Mk+90EleD+ff4Cjp84s5tsl/IZK2qcHGETlAs6ipSzHps++DNZW7IHGJ
GuArNz/lfiQpbOkKezhYlGek6t9fC4gEiEGwrqLwvWFxjnj0qnIH2Yj4hmgNiLD7WUfK2hss258X
i2vbljdnLBhfq6WVpsMg9aQ41Pkfz30KKNjaRa4il8C/cKbj1NSFL4xiCENSrn80T3JrWlytdr+5
jcg09VjKBLOh66i8vRIzgN9fXRgmCEEG1aum+4ZDyss3Ht3c+NxxyvZ3b99tq7H7/1ioyObm5fHK
IIq39R2sqcpQTSU6bvVEQQgm0/jqVVTrWCncxcVs+kvlpcXni1z/aE5IMPqxGT7eDcFTExBkk+7Z
IVN998HOJMn92e90kKDmBB7sTGljjalbv9buRtdS/RpBekGQi81dJnoX4xTOClQKmPy2MgHzzXgl
bNq/gEfDwwHqUptikF0VVwoyChWSNQHrZ9Sf6gw9zZd36MqBMy5VyuVteh8Rm7TnOSJEVTVFYaWl
vbxafa/liG8fQ1TNBkdU1BIO7B9/l2Gc9ddFDTAFsVj9s6DpQLIYdJ1EnQxscoKehQVS5Rvf7hHv
klZe7SRbmEHy9pVuRL3Wcqws9N+nK6l7QeZIvNQfa5lpQ0VzwZRR75kKp4oWAnpwoHGUzLQ9bj94
5ZylL5s6IJff2NDQsmXUn4zNH6fFzuMhCgEuT35si+dzYlR9IiKYyUSBztSQ42rnCXicnuIIHBri
pSsqMCNTjvyjxMjOZsEuVz8dDoIqhFwvJBc4iYE22hoZurR92CcYrhJTOi8T7wpKpEsOPYscFcsp
LbHSXxxcFT5g4+C691JHalNc7cF/V5roOyACyf1tzyLjYlYimeo1+ZZJKf6YGeBEPbAjurAlrkKc
RjNRvF50uEc675AFd0SXiLfkM9SWp0kWpUhYqc9q1FRi/40Y4RyY0O69sw1ZS59nz2tRcBG0I42F
9e4ZlCiFbA5fLsLuErcCYvfaenRZmywI0GHpmznc7d0XUGft160riRj+AKDOXiz5YmD3fon8nwfO
eLI5IQoiM+kiQPvzeW20P23mkra2jnQyfYBT5BubQt4CRhTfg5rAYchE0Xq1tZ6RRVH1LTYsdkR/
o1r5/v+dI5sFBDcXChSxNxnpJCb3G2+2o46e9TiKC5kLTDB5afjF10XFgP6NjtK+YKeXfgvbebuz
dbJCJYEi7JhkjLcqCHFtNQhQX9yOpVE2lSouAa5FESMFTY1kZgPapeujlnDtF2sfh9YOsqY4KRv5
ZSYlr6Fr1diinwISXZ3ulZl6GbVrdx4OO0ONeqlgOKQx7wBgAjMu6urRi40z3VksuG6n2nHz2GPs
rNpOmFsP9kXJaS+X1YK0YlAxQ1z3V0YA6ChSSiyBYjjbm3/efNlQERgkj0dQaJFBcTdLfyBFUcad
udhtitMFYLgrO8mwDn/RADZIMyP7rk0p1aqTfa5rKeGdl+RcUck/m1G2a1ONZUS+aN6Ew5YXIBBp
JqUC2hRjWe5TIoIwmubWGvGAaxwo/Z354QBc0Rm7Z2SPnEixPUhG30A55WguiPlPeX7ZPYYnMWO0
+97frvQwazYoQ65Tk2xZOAl3N/BgK07+3cYVZjo8jaOSYQlkWvHtKsn8ftzpM6Lc21emBVvSOgWP
fPQdSZ52qRLtS9U9Xx7GwjH+zih1j9jC92BbfQw/82Ym1c+8Jf9tvvB7lxJ2rBa0tLbUd3xhUiCh
H4bnUS+OnS+rnidigW1ijTCKne8ezBELClGd9rH24enHfiwPic/2D423qI3mQGKqIGcTC5BtIdVz
iXtQH0wVA9RqHBXIqEmV8GIoLTqKLKISW81+ptmH0yasCR1p70XfDzfw6/CQNM4JIKfKzTg6JqZ5
D+9gxfGgKoUHXW0+LUZJ7dBKJYcUa6gHrEO0QBzMcTh4dmUjnakYjFJ/u/dZrUjwGfhEs2cLMLcY
vp+bbXdWqOm3AmpSd49O4MgyoMeFkGI0Wxdbkt1G6fiPyFKnKBZEAqwnYoKCF/3IwMpjXzKuqZCr
kYTaaj0ctx29N7rB3/y7tkB1OU0QpD7lmCOz5UDZxvgxmzLIFSLpiCGTI0qNlTQF5AuuB4b70kLc
VzXs1hCAGEHTIzOwqVSE5+HnlHN313XfVp7YRAn9RgW4+5b1FxJpdsH/mzGY2lzMLE0sDKjUo0yA
tV9XsTm28ncBaAPdFp6Z7WCUUqUGzxFS16p4DHt74MALeRsai72Boh+VgMMrV4R+EPxhaN0JKDFT
LwdPvBdEHSkSHo7rntTN0v7GcHrLRUPLUbr5xgpi+UQiuySKYUXnlDYH/+bDv5YFrVx4PbBWTcu0
4hiaTETpNQ9H3Rh4ryz3Kq8wO1xiGnbxm1Zmbxf+lqgs/ns2CyVUB3AzWkYd8BR+hjTD6JsEdTUv
SYVBnJhjrFxQuPq6RmrOvp9Q9eKnBtFR3o4rQZPhB90bhM0s3DJS5ani1u6ynB1/Fun+LIGUNQJp
rNPP1sBW+xVU73lKZ/iwZvjnUcjMIss8xgP7FaT9Vkysx92mRAnh0bl2b9J9vKjl10ygpafDzFji
OIqio65jBuDrgEGCwLmRWhmywSHe21Mhya3/ha7NIrLwBoh47sGUXM6sSjNNzJb9teLcZM49pfO/
TLOfHRei1Mj44v6ubPyOfauRecNYxFo6sL3Ts0NtyRhdAMw0OPc1g8DdopsY/7tVAsY1ZYWGW6+N
7w0y2ya926shNsjT2ptKBCOWPwNGEAnAIN8jH3LaAH5sNG69w6zyc5lUGFguvBxJzM/DhyhCrtsQ
uFcb1ZDu4cLDYop8hoZf/V9vSzIw0i3S5/G6BRYzSumXqN5rVkChrcIWXcc4xv7EVnSI/75IyehR
hwgWycuWEIHU1PhvsXkmReRNSLNpCgxncqlCWnd69aqGDy1WT9OZICWdgAFU/NaRckPk/uk8VViy
p4dBHZS+ztMI5xtbQ5L/1Qb8HDHT/0E5SL1N4d8QCwq9XnTN5bCy4WLtangfndjlkVI+T2OtTxE3
B0UMc5/AJX1wS3vLgRq6bg2bIzHPqhHxGw4WFzuAy6hFA6U0PEzyL8/NyZx06SEJgOUFrO/MI/U2
J/g1beK0e4N6zG/6TlLoVv4azUau9mV38aYuLcSxzJfz0jaVz7eXnKe8uF+0Pfm7FuRR39uZwXrM
IIB1FKY5EFAiJWqgaoYv5GAxcccqEaLGM05FqZcd5xleLirsBwDAwhQiksMlH6bKd9Nt6qcSJMe5
xLBakdw36nVYfc/ZGMXilzG9DF86x7HSuOSfLG3gUPZrPfHR9axGfPvWmbz2WojxMi0ts5i1O7lp
uVJJqEq1V0X7EhV6LKgrkJGacCHDioxtokEx3miMK0RhNeoRoEcyPD1iZ4uhyPgglSEvpBmitR3y
I1FaT4lv6BWkyhf6Nx/tXDvcVielAMryFtu5Q55VmE14V+FB8n07Q8Nx9Yi2XfG0KJGoTgGmb99y
cGr3wEYqtpLRxsCUFuwW8m5N9ShWgl36Na42nPpvwm+pEmb0wkw4bF2/lvU/z8SE4cbuUVEpFewy
/YeJm63kESgSBeraHbu4csaWkmo0JGX1Sm5jvFMXJ6i3E/kJqozj8WjPaBYW8YI6gqUMZgW48ETW
UbmPenDyztU8wzZewT74A5ht2eGu2vtwZQm0WOebUPzYnV0K5tF+mYVDlNfVatqQGWEGKiSHq4GH
8gmnm+oDRkUIkp06b2xjSjhR0tRDM3i96FNGLsJlnuXR9zebaHJdO4A6lF2bh45pgRMJTOMKRkWT
/A1LCB6OiVwRQ/oUd9uttxyRuuzaoYpE1RB1Uw+kyqw1AF+d0HLQ4LbUOCFCdx4QA0/P8+FJMWCJ
SdHQvx7j9pUdecCaYGtsN5wjY0Eoodadlylk+htKipuOa87Z/rwGeSUfIFVdl8Z+z23ltkUEitPy
tELksYP8BFsrrzql3sWnPX1crHJEbWc9VhW1wRfcqr4h26Omg0nSB5VeWiuABw0P/nV/60oepkfI
zgRRTlw+exPZ5E0C62PvSkoC8ugo2JgHWDw/dYa7nZxP4H7EkhaGwqakF4S5qOR/UzIeSTw4zbIh
AIickJoKd4RpyZ8zs2W8uz493mZeLaHJq04SxKudxxYtoNaWQxZUeRojkbFI/zpH9eCclXlDsYcB
6wsjgmtbh/gU9o7ZWbIF2cdYEZEjfbljvXasTHidE33dy8YND7hwRJHtae7FELOL0Yu9O4xtEcLp
Lxm8v9xB6+VsQ9eZ58oHD3HVZDoNhMpoNmDMQX6YCWAquKyIsBSd7UeRo+aJmEHKvn0TWnQVHqlx
7o0q45YT3znM+34e4EXPTUdG/6OOvjMuT6z6zuTXCjaUnVs8IXZ8gvF9WAKvFApkyzwXpbHv/C1g
nIa8Q2ZAOqO+qVCN+aycfCqbtn3YXu1o3rYHtU5jX3pWCbMSPMx4z4EUmNkpLWbA9PV47V2Q9Xge
yaBOqc28V30KUGjCy8C642sAMuAwbiFf+rQtkj3/14aDueDZ+2wRwGG533zhLLO57uog2LyT+jSJ
KrQYNh/QbBUklMkhC8WdpMdO3PRYRPe6rL8LsYW+HenGQpvmTIkoRRTvgVJYvsjJp00D+RtS+yZA
z6LDwYn4jDbluB/3Rhrr8VbF+h996n81z3RmNFNtkCMd+APlUndMK1G+zDNHTjeZTJQ+f840iCmM
Ste+DeV4+tjql5RC4JRCNc6ZT8g73asFmOxYTiUrh7FCnVuYJoqOGWQZau6MlqFfGIq/yFgdAWWo
u1M7W0kbK/b5oVAFZ1Pp4RWkET1UcuIqTcjckNaHnpuCXAiSl0P2OshuqIXiViYupeTAW1t7lwY8
Ajx37mIeiE4v9pEDTXquJyDWS5vsSIaDcxmrvEBS43AA5Hz+2OgETeeM71Uj6uPGUiHu+C8ZQcJ/
xeLXiDNAI/srgUpykXta1Mc2VCkxf8dANWxxn7k4Wvpj0ihe7h8ir+/53K7NUypr10W17u6v18sY
4Jss/vkajcrmQjnzpXJnrJSUM8EXFrSNmtJfskHEt7hta+Y080E7hRXygqLbD35bNNwZ6dDbYc8W
nbPjcnmahOgsRV+lEMmDI+jRQ5p/cplEVTSOgCkwMmRc+VDlQJktU7viTk4PzQCXPrglk8gQ80DB
p+sDEUtWmDhqG724pYzalaEK/V8FOW7ms0ENQ2baRvvi6+XFVriWSVAGUdNlQ1WkQzrH9IK3RPqu
RtQkuSJMnKo38yx/lYu5wUdyG+2oKE1sYeUFi1sgniiysRL3wnInbb+02HZwZ/moEoHBrwhWSGtj
Cc50MnypKd2O/DW+/wxqNmJYRjLPjXiPBk/Yf4IhjCOLjkah0nzWl0rHjhVhD0Cl8zknF7agpHjy
XUx1lohG5IgZS6veNORZ1pFE4xU16uyw+6toeZ55nzVfNb0sxi1KtyUoHFDIqIFrqIQ1a2l8UZo6
UNUP31weXRAenvByFMird0EvTyGUSKH1Uax0x4sCOHMmSwQQzDhI4jR7UAi3UQJD9uj+uTT+eJ3P
pA6BR6DMx7VvgaKcUxj1gRGnrFpQSzzpc005ACJzO/MQB4FQIEP2YbJxde1PiYFUSWyWTTG1o2Ne
QvTMOSyhY2D1mkzN8OAgAyQNzefery+r5melEl9ZUXS+zFU1kN94LoxONnFO+wyT3vg/9wuedgIb
gh1zneP97bvKvU8qCWNtkUJCyShTSq/YmfNKggfCGgqPXWPp+KIE9Nvvzf2BU5vVOzbzVfw2L3Ql
icOFRV0TnDz1DGYOMIUrIzjvQXlw0mT47UM5hJdNPULyqFe38BeWVbKcErxr2q3F8AVY7dF3d6ME
V2pKVjccUchYJsYrmWQkBRwKIHuC3bcxL8ZRYUIvbIMdRo2i1LbqxxNuGPCLFeurbnxoiLgGIXiP
v2hCeA2/7sYtmGvZNvMKww5YPpH54PJ/NQJDBFCUaxJXLVuBwkSGvEZMLxBSTWKvN7/efpHzyx+d
xe9twhkmBuFWcNE+QFpdBUDAVaEO7eP1wEtDMS9IXMdB4oBAVmJwV+tWLnvNJCiulSLtK81YZHIp
XQOiGR9iv2BAGxG1VJ2D37gXmE0kYVjrx2W7Zxr3V50V+VcQZ96gDNFO1K6cAw3J/wws8lUhf+I8
O5D2+ylckdTVtU70aAo+YpR8m8LrZNSg0tcP5mGQAQ2DN0WOLyya5XD7pwDCUVyXkDmdKGcKyezS
gg4NBSiJDW4BJNgC7NY/hXWUDWOB+UYHEzwrj2I3Y0WzrxJIdJy/KC32kfq8SwNsAgc86t2AZmJR
7mhKpu/rzRR8QZjlJaCK42tuuVP+ifqHCpye4l4caxxZaBJvdAlwStFbe5r0YHQra/5Pihw2ZXo7
87JU+1NgI4ne9aKFArfpOixJ/tyNNytdvaZ1ptm+gYTKwFEXVahKRYXv1urPxd6X/KAF4NF6cmC8
aBrxd03uzzdwXEZSWov+zT6pSTigbbzUsIT7ykmBC/F8Di1srOgrLfPHjpJhdbzayb9MNmoJDhBG
PJ88kUmXgBF+zEOdl+xTCNOEatnzJU2caByovX/SK8hXd+RVqAfyNffuuSsRy2jqfNKh6ookMg/0
ZJ1zeuTcLDgbth2TKdgrBeZSDa9+OSOH8GwYsQ7I0Q9CiGjzk6rpSYSH3YPSuqiMTib++1pd6p9T
b6QEdNYxsV7N9XPFfsXksNroGokAstQr2FC29sLo7mnSmNjPKaV6Qt7unIam5p6iqgkcIjpKLskM
o0M3oFTRtWPziEZxciQsmST4U8mqdJr9KsbNoeLgIT2ONqZ4YJiNQ4/2RCH2jZ5l7nvLxFUZ7yly
nfQSsridvnEq2S/FxF0g2jjzx/bTgtZB9K2AxDo4s3oLKBBu3qPzzxiAdZB0k2ndtkHFeyKPKAoV
Nj47O7wC63pmYWqY8zu+1eE/JWlP7m9c8rPmLGDxHZdivSC9g+ugKOWU2drtnytGkPzdR3AGTQW7
1ucMdAtJk6Qj4CzZVgW19EDqnFnZ6JxBn7xNXWBOMVJ31XaTu9ZZ1nvWuYPiFBmIVVB1lbDy5vqO
+EH2RSmN+yIaGIpT5uZcpiMk7508gXhuQTWevU+VuEgR3JpcnNZFfO0xQ/2bSZoyF9JNT5fLfO07
ZfQaUeVjsJIrd3kvznk2MbLh6x7opteThhkbX8tqOqUirD6N7jT4tnYipNaKcGodSstckVDqjxMR
fFiDQPj3sckkYpPigQsL+A2KoOlEZUmlL9qDNBw+hbZJKIZfZhZCbQm/qHKI1GCEjjmBwWVbDS0R
/9g4CwYUllutrpnkV8mVB8dWb3PozMguHO1Z6YIlLqK3p1y7YYI+NWMe4EFlKMGddnyWG4MeQANz
pwqf3CrwdC1mZlsic5s2U6x+hWOFOgGRuCWhzRKY8i2/YTNyX3rHtTzTHTGWZNgUQoBf9neWBw/X
hpTU1tnVpZcboh2u+YqQe9LD0GeWdYpkGvVkgw72+WN9fRlDVxhKvKtoC61gffqDVvKP7LkDPnSe
JCDAoSRIv6xXcJ609Ce/8tHRS1MsC7uCM8TdO/+Pl2UGql0xXjra7hpIpkCegLuMPlPWa8ZJc2VG
58VtBH4iEiFwIwL+H4YsEjrjwULyDWaLso/Z/+Rv4OOlCj2gKulJhXP2hwM43qr1m/ZBjn2dUgN7
uKPhAVWF5eB9P5SV1+ZEw7d7HdsVIUBHltE7pm6eAKEWFhuz6tuZBrfsITJMvnptFVKihtMFFe0E
m7JF6jQb2uxldyqmUFwLYjLw+wme+xNPnCqxwA4IjByK/GGe5C6P/bpudw1HEjJOM3RlgCVWyrJb
gFnw0GeAwWSLVo+zTJK6nX6qc8pT6YXMmFv3crYXWMKt5VnTRUGqKgbv3Sb6qh0HWj9es9Sy4W+1
VKyARZ7+KvNbzz4mY3egLnO/YzAEHdoq6J5xezo2yFkZwD5RB+RLlosaEyU5I/6qI5dcsN8lTREX
iPL+L3f3akq6ZtZRY3sNUO4V26eA2sBBL+I1m5b4LJaBsNZQFDYbOPFo4yPaIBDgHBwqURa88vGW
dgfn6YPyuMs4hwc4Cd5GvnMWmmU1NkenST5B1YiCua2jf1+z4q5qc4MaD/+bqjCcCS0oPjZzPTbk
AiMMFPsQRTXOmQ+iTAsFl6n7YitI0uyE6mmgJruC+X5Ayy9yLBd3okxt5qSUH+hD04/vlnZlo++P
yGPgzjzDdYNU9GiA6cWUYLWf46p09ZqWAms1pV16pYRUFPXOHzYd/wbeg7QA29HkPdSC2B0M++bQ
QBNYUJn5xIJKfv0uUARjVFfGF+wtl9Qt+ws4MD3cpjLWKzkm4p87+UBb263uS97KgoCjR1wf+1Jr
V7y7UnDR5z2JrDdO6xg5igzSesMe2rrWIOlmX5nk6XhF1Y6dt1DC+n80m6EY7dAsHqjbCVZu4uqj
zys7M0sRY9RF/3Rr2dd48ATURsMzbx+bK6Gy2rJHiZV4uq5dG08SAbfU0RdxlaLZ0qMuJFntNBk5
L5VNnz1a6zuim8ZikkEKGbPNFlO/tZXLjlPh/2crFsYu2c3UjV9Z5YSJduZFzvEsQO9IAKxHJiJF
O6U4NdpzfDUdtpKIWzYwkmiuxuDQ1/QkOu2qepnOWmnFDScvbsg1nGRhVIlqR10ZxMDT6NmZRtMn
bwsdx+TAiSSh0i3Xqjj3k6LCmjzvYe7QnMGrpyx5wMxn+VY9x88T2yHy15DT7EJx3FCeeMPAZoMC
2Oj1uHtxDrGj0uwPjLJyGKdUlu2wwej/QMntP4a8jfeSvWrihcpaV3wDJYrJ3lOY0z+r6a3SJ0kB
UY9GVJiPWH8pYtjUttKTLqg1EAqDZTvdkuVOWQfAE0/QUYLclG1H0jCW3VWjEg9NyEoUOe66h/0C
n5YRJjkJdLUVdA2AkaX8OWh/9SItgnN96O4sr0c+ReowjVIXrGX3L0GT2S4rzee9srrhHAfGh7RI
lGEnmn/PqaH9RkjSNY5UkaKjEeBUMYUsc1Mr0yVwmMqz7bm6QUKTUxh2OCwjRcZI634vdMeqV8E2
n0TgRKxglqmf1XKHE1F1MVuOmVKfrQXzgBvkF5p9PYoZsDva4+9a7u3VqW6fqiseK/8nMDPtjT3c
DD8CViPhM9RXE30N2ZU31UgZTzKyZL7CaBY7SqBYUEpRTTO8OXx0voNDYFOVWKN+nSHD+eUNm3ch
0yM3y1huzHnv8mwKrwRJVOoDoEJTGiK10VMdG7gwWR1y7bbWSPCD1F4sUhEN1Ts5uD5JLbroYyuc
uvOtKKaoCdkIkq/DJvpm4LYL/ijioiw0vvl4CR1n1nP4it438PTPKXkoVmXVnyrir+3XCVmYuCzd
noAFgnHjvVevriSfekcMIXGE+ZlpXyhYxt7CllucpCSN2GB1Axvyp73qeQr9VS+DKSqrL9zAeQv/
eOKIxPMH0SOyhWLTsGIyW+V4WIG0Ed/M95lbXb++6mUBJTgKbsXtSB+1SpxOEcVi6jO16e3MSiLc
vaAvioLbZfyvWKdacjic+9bovs8yeoc0ZfcXZ2GyY+fkMlZpjnfiYlCs5CsztQBGvczdnorJ2jwd
SU0qPNhXGZEXQrKkYTUHurwEh7Lt59wStZERuYiYKtlpt1S9ifianCQKZ/vu2wFZvlK2WPhP/QkS
BoP8hQl6ViX8yjQ24ikqnm4RS/saakAJOzGtx+jLWum7dmMdkS3tHaj9XYWTfX5dTvtbb+MTzCi9
cdY/wQecn9bbBnVtMBoFqnJqSbUYvNOxjbZIodhxJwNY/683JPRhhruuWLLOVN5UlzQPHcG2jAZZ
MYiEOSphNMCSqxsqHHuELPOC1+sQGAq7KJoqw3WST/GEuNGZE63YnyidacuUUf4uOYb0Npa44KS6
uf/XyHtefG9q5OZsoxOC2kkIjw9PQZ5o4bLNc/C/smQqHT1PriuMgKP0zEzsWYm0jtZcN2Tb8kBv
wiysZgpN5Z3/CxDkvH1QUkVStWS8YRp8NvWmnh3cT9737BfNGTOXgkkpL0z4zfKnq9bXOjFE4zFb
y5D2WucEOLDN3Cxu8dCCs01mekLbx/LBjJNBfAsn7g3Ba04/XtvZoohLg0j06ukmrYnBM6u10BBq
eyDax90dZy9fRrX48VfzWBzyb0efPae8WU+vqd0XtxsDj0wFiJWLAoWDMovnimWQDVBG1r8KR2nK
4MgNoRyteFmSChIE7m+egLRgVDOSD7pTB1OEWZzZzxd/0tua+K7nC7lvo44Tm4XhDhn+ipvCNL7m
CJzhXYaZ8RtMjkBu6KUyX7MyBJRNbtjfCDIKsWcsEM8G76KqDbDs96TqhdD7XacbJmImKQfg+dmU
DQlURK7efzxCT3mDV7s/K/dZGV2+UfyezsjWZSFYh17bk3ImA9TRr7khFlvxgiMJHl+thSzMViFd
2mK+sM2qWa6/iBLTGF79REI3jo1I1T887d8sLV6ZV5QLTFuglcnegy/Mk3wmUAWH4HYZ8i52b+rK
t3mBI/vqICWyScL53DaC4rDx/U/CDv4VQ5lMxvjYKIhTcOcWo/5gpf/VoMNpZ9CyOR23xuKCfVGf
z7yhOjXOeBq54R5tjHioKSkGnn68Dn1jDyzmqROFHrcOaoIIB0S1pCCHrI515SbG5TsTpOwOd+bS
bter0uGCwDWT0BXRQC+Aoqp4Qzi4CFjHeuEnnTbvQwRZHp6kWm1ZPv1hq45Tg7VZLkaEpEB+l6EG
rBTq/Lx/8xRsxwZCIPw11NVYX1DBi6T+WwgRFq2/0JgI1oeH2sJM1fxmC4SznTfc1jaB6f3NV33j
1ezNFk7wDFytDK6K2zh+KsunTh/Nb7BEVvukuxHuIhnoE2+we+OPUNQA0S6ef66ykmMws0mc8dMp
9eShC5zA56Bh9A+28JN62Od3kt8pZbjE2WJBow92v34dx5DXpYNg98Q0CDa5iTeKm7TssmBJRhdC
8CiXWTJsmZTJ+dojx3J6huFOb2jRiJu1YtwoOtYg8HhSBbHlg/iA1WUOpcSNR+5cYftANgic9oO0
gczOrHGvNxok8M9nYpcrsIP2XcqqjuVe4xjAQsfhN//mMk5XS2KgUrFbPBg89Sv+E5wgZxee1LnK
mTuSHSN//0JlTMjVd3lzhfCXXfeHqCO4lhUwhsGkSTvwloow6EbCnNnwmuGzSiPeHZAl/aHGHbV6
ltHKA7Bs7wgvRuCGH9Vz8X1yu+U4VTz4cjugH1pIk9a90Oy2Ly66XkcgGwEq/onZZBZkh8y3HFzt
7l2i/qkGSYUjYOx515FrXJuKdzc6SetDKtxcezixS05YZvaQr77EAUmD+K0AO+Px5GCGmuPuWyQ+
TrDgozzUulIay43mAjUKcH5exgJCvKJIBG0zWluhR7wjyZmNb7xLR0lpbwNHgDFACYGChicrtfD+
og3rx31aRvJv9dr4c0Fdk6ULGhaCHBaEdJEyjuYsDa+Ky6CDDIzIRdnnk65fq95ljRne/8loiexV
lBDcxHvbXdvEnByAlHzh/9MNgaRv+H2R7ACmo2n2QnqLoHlXQHv/+q/oqSss7SdMmXX7QaehTvwJ
7rVGrBfhJ3U0x/RNMl9KRfV5Fwe4VTdbKAaYmRDiUtrbG78coijrp65eZGNIjvnnyGbrKuXe10eg
gIJQVhl2ec37x3P5tdULDIZpNMSGj9JqrlJJibqm8oM1dGBsasS5rlkhcJGPe5m9OUwhTpao22g9
pWY4tJ6Xr9eLN6fqKaOKLAPF1EFCPpcaErG++qcox802Yow9EH2efG8Vo/bpWjc40phERnqA6At6
vwwviXfKM/kmZnkLvoGpjpIvgLf7g54xeX16lrZFJxfoRrIgdPyhV4QLO0FedmXc4P6n1Zqd5ZD5
rx/N6+kbyRCe38ku8PxJztZZb4Xo34eXWT3OtGBhSHnMNQFXJ9Tjui+DbCtmOB/aPhCLL7sVRNBm
ANV4BjDEwZHo7E6Gvdl/1MAdn07+YoGNKAloOqHsz6SsB7QcwRaFWkF7UoOeGFh0S9sjPjEjMBkD
ss3bVUr58SUjVXkp8AnNkp5XbiHAgVuaD6LBxUTWUqt7gmBePvTexHk5yuxtaHZzfpUWqFd7ym8E
shtzho/h67XJttTfivjxyexZVQ6LDcWvdwdfDCwPEO3W1ijTHFd/KgSST3OCYO70dmUNR35nGtcD
KAJKtxY0SqfmOMlqAGx1GxeJ0GV+AgLDP5/ePVxoaJugIObBa886q3QjaJiXDsDdnudSiGiGAJlM
NhtyFLW5GGOjjsBFtqjFt9bSa5Eg+Wy8gqLYsGV+7veG3nezF16xn4zjde3JHAmtU12aystIrWNf
VbGqffVZNx1905KZXZcuTKLahqlpVSYPxx3/in1hcx70HSxECjQC4K04wfltPmPCE0SaID6nX6nn
xLusB6eXHeZjP52iQXDtPBskh79G9dkk/phHrQ+Mq3hMtzdB0Ua2fR9UdPau0oUm46k9087Q2crf
8lsPD7xuPFiyM5ASmTYpjagebdJZyye9y8gKMjwcZVwW/osG3GTubZLd0Npna4w20Izsg1qAFyD4
hw8ku0tsRPv2iFWPdthW1k9OGPvmiMTXa1bntqBxINZ551XzV1VgG9x3u6ejfGzkb1v64dmQM8Hm
fO14F0CEHyUIK/i13KF2jyl+81FdwFIlYQarpKV/180jpn/bgQSSpS1SdfK4kHQpfG+EY1slyWzh
JCzOCAWd7eL2PB5rM+X5rx9Y6mkUvX7SuLB+171SkGO/tQeQ0RmTNyTOY2RkEu9whvXkByDITPvJ
vFjVw6YTfgAxCy2ndfXCLD+m/5piLI1Yb9vp96d+istqGblQOtHeEvkYnZ6HChZWg49e2lFlknyp
yOmwSAZ8xOA0CHT1Duzzs/p9ZzRpbbLDFc0FWG6nH2Yo/q2pYsXRPi/iSskZHiJlk4SKokUYOtUI
s4hgkeJdmWK1rZOUyA1sTpRCTf4XpAbD8cF13XsRLFzkAmiNV4d8TdBCjEy4zxfxmd/L/9gDO2VF
2VKu0BvNAMQ0mf64OZ2Qaqe3Tpu8j+W2f98DVlUOPk79dzd4YXsR2N2NnfV1eJiXOGSSN096wH8l
gQ9Elxq7xrVce/9l7octhV6ARHeCKGwaGEhxZzRKzOZBvIbamWdxi67x+9/IiBdXdl7FReDaniGO
f3/VTmXS8VvBd3PWbapWAPPKhhQd8QUEs4kuWVILPX+AxxE6MgNg8vICg6lkuuvNfXZ9AKnL3Szs
tS0EJZ26xy+iwolFnR5/G+zXIRBgfdxcTdi16rUonKkqCHWWEQ49bFRYAnXOseQqsyp/fWzt0ucl
Z8kgaGmgoKWmKO4S90rxD64CspN6zUE5sdrJhoHXO90cxOfujuJTwuw+ZQsYrpOWPoKj6i+BiucL
mTXCUbNh90HuX1bJODC9ibTDVzKQ0qvpx3/idqDOMgiFJ7NzQVRbw6VOrnroAYvODR4O/Z9Tqzhy
9xWq/ZN4Q8Azcg5x3Da2QG+fU9rQUMgWw5en+YrKTBIOi4prTY/pppUF6qFv70cTHhmpzqWAVw5X
m0nWEPAoAkglNNW2iktyRu6VYK73kaCWqxGluP9bv/y+JbfEvLnSTzIhc6Mc0L+MGRrRsCsvxirI
NullzRLsqbrzMp6aAZexU66yA5F2fhSb2X6hHLx+OtID2L8VfzAvMEOKXbGZpp99sxTbElI0PaRi
RA5f982KbxRi9Ku4o2ND0SOQjjQHcp8T+S33zb5d78BrcLQ2qGKl5NH4DTi6hywpzCkt80EXMseg
e2zkYNrHNpLi6Uqe+Sb4H1TXFmTjH6kK0dJtVdvowD53tzG13X+MzWFVh/ciq6OSfzFzxNDoU4b4
RdKbwlKsJLAXAB9//wGrFo2BMLKTTc7XbjM9F0qn4Pt/B4owD33OspCnZkWizWC/50u7jzhFTKlc
DMx782zUonbEJsHOj7doYLyW7sUyDpYdEymFL7VMgDrRBqWLv3opUsJS3o+nBhTboGnnBUdCo+VV
98f132h5AFKN9/cXRmLNaw43Jsd9o/ElI7eePH/4VXnLceO6dbXHOh9KIRECrZN/SgRRhvu/fpdS
6iDNOsbuPm57/5kTfOzO6P6aqCkMpbaC+V8OKgDwax3QS4/wEt4WZnRzXNR/F1MQPoVUl8PG32fm
ZrHmACOaB1Wqcr/pJ0Chvxby2TbvRengvLPa88nlGLEbDHp3/31ahd+8oc6PtBOAUkU3XiY8LTjq
smnMLsaugJuEF1ogxWlT1HChdfiET/RkPVfPen6gJSg/Ed/krvY0bD51DUzRTVZLcq44i+2tG0g1
NsvE/QEh02fU2o/2mUXPmrsWvMgLZYVySTPYaYS0mWz9DsbfJSBhWUHfnNcN51/ONJ+gexSs8+nP
S2Uyj67G6IcqSwUz8gEdHOxUDDZAXhWzLbOeRmL6sHOLu2roConRnk8yP85xXSghFuhLPgus8Cnc
PQGShv7jA8KBGoRjz2BXGTg+gwdkNGEagRGmgRDCwvgXAJwI1CckITBvlQOSwcci41L2zm/znq/h
Bn6VXkggLCuKRPLvCEmcmtLrYkQWLzf3QwtjwOaOMEKJOoiXspHPbMqi8JrmQn3HLTf+8WVUHwqI
EThQ71/oGs8OE1JQ/RUbN5u14L2lcZSnqJobOLcfnTKaPOVJwVTg/XA0P8yDikLpnVBzQADvKSUW
2eXaTTEZ5PFvLC4+inANXT40mHZBWxjdleh0oX/CX12S2hIAqfPymPxGpguGm2K6uoG32k0s/thr
B/NykVHcTfOsCUMvJA/RVNjwq2q902UFcW6g2zCktlW10ksc++HVRjPbWkvDmcmDoJ63njYA9Yfh
OjQgcUi2KK6iDvWO/udhQZAdpkt5FdZnromJPRb2lw3QBqEy9vr2FpJxRMBMniLfgeSqehFlBLzt
KLlrZn6YHawwxP7rDXBBvkKWO7/YYGrpmqoejW1DDAoKlkjKv7V+PkRfNHRHiFGzMSZlrzAF+DRr
nwzr0hzQ+/Hx5L6V9j7T1qQK+Hm+vYG2cci+oF0cr0sBCQcw7iSL3K0RY3unbD9PsfdzIJxx1BdV
qTNy5es61RotFCJngQ24C4XyqVTVlVH4TEKStjJcdkfIHjwwBZuqH4ItOzFbRADmGinEHyF3KH+y
Y2kSLD1hjrseJYSxCTmBWsiPpZHLk/O2rv/9OM4IblwxtjQXD5Y5NB/mXtVMaUdRvIFz30Yz87no
ZlF2jaPQ/kVgCwyrz/F1xd62AqzKPjPV3iz4Bd7bOi4VWBnvykVVCfpgyP8je9/SY+Pc0vg+zVc+
acT/Yx9uXe8cC+7ZWck3tF1u23WxX+RRO4wlFSrh37c3GDxQamnlxRPGAfaPGq0Qn+RSddHtdV+k
7loZjyVEGmdWH3z6X3PSjk+Gw8nvgTuUyrh+iVgea97Bw2cppqO0iy9oU7jDrgDpdijwGr0RyGO1
8LgSbVPjriNsPoPsGMPeg4ZRc1gVSdDCHUapBVPwtYpfmTUA0Jd1mi8WOc8sGU1EYOgtCrxVfOoe
okKi5Xw40Tg09JmZD/Y6s3RMT5DfAFZijbC2Mc3q7/rd8V0lF92UPbY0KtIzNeSwRplrRY9lHe9b
3B3lLtoWz1p89TjIL+DEVQmYyOIJrZ9y2iE+HKwlSqEs4OdGQdDUlxO6boZQXziLtPZflUSDL4S2
Sl1z1wTpeegiuMB4p5SBWUJM5L1Wh/iAjhGPN73Tgzleuu1cHM6Wqup5dvyPMtSxW5mcbTrBtln/
satowtl722hlUhxS/iASow9wI29uhLf2isAxs9GVvLBJcARew/Go/N5p9EA53IO/JD2EreE1ED09
z+lpWo0u5NpPsLWosMJYE2gNaTDv+ELGrIUkXuqvQi4I8rhbuECmKUb+iVUopdvxl21Auihn31MV
UbjGomBd3KSbI0cty6cvgF5iJeI3yPm3u+WQntRChUSxI/Ka1u6XmfddB2sY6pm7LFEEm6uNfJn6
YObyNY9P5DFdZxYE9xOiGKvfvl0bb8NJ7zmWanfOvP0flgrU3VXJFYPZiQ70W+mXvF2kP27pYiZL
YFoLSFlFx73GJmcXllsalSXDT7SNAqbavWLCYlhHW0XakHzRbY/Mg59Ef5WgPnolX0SzF0z6mAtA
b9jueriDRj5az80cFi9l2kCoumOvUyTVIqEchf2UufyiMfE83OVyrmPvXiVA8AT2I02s1+/jeSBA
ilMtOMvl3JN9x7R/q6S3bqO+lLOHzLsl3t5JE1sIqzUCFsaXRiRhGoViIiOizuSozifNjyzPv+HJ
hpRnP8IU4n2b9OBnpaAUdLRiBw0NDwmrbnLXJ427o0f3SM9suoo7SCmJo++YaU5Q1OmhD/pbFzeq
AUcOacHtyeJlXPN4K609ZDPFEYLSP6wktIwQXz7RG6vAb+1yabYGBs2eryg53mjdeF8l5139AiEx
5EO46nFnoC+QEDoOKa3qdItgNBnC/g6pHt6CfxP/AmsNrYYvqbjtFKZdtPGIUbY6NgQueZi3ceRL
YbmjU6q+XNqjcRCGEqIemDW6FhtQVBLnrItETbOnfrTYmOOUZx2JU08tWY/NkHdkdO/PfxxdbYo+
BYGICZsd6X5VLFTs/T3IyF8ZaJNv5mlZHlCw71P7lInV6mnMD0NXH/pbE72LJ/mja7iIEE/bQQvj
+ygC2yIC3mSxSSs0J7vD3iTmY2OyHmT5/HARBK7PP2oHYo/Ah4cCJXU+F47Tr/vvl3kA2OgljLkm
BiLQiOGWqtIRlZspUXl6tCrZ4IwYdIv2+tq75tovkWaJNIThLG+SVzx1kGQuBGWMgYTCdHVTTsFi
Q/50edb3wDTFgnmpE1UDliJ0JmbzlH0xDgBl0lkddNFrSDfnAZOLcFYlhS3w9LyQDY0iYsdA+t5p
1k3H5uplXbqnNX3zek5b8unORWN+tNybO/6M6PraxgNhVAwqSItf2rh8s8SEHeHIUvLCsO/hrXmJ
/u10kJ6VrjqQRBI/UeOckjsaOgq5z/UV5zwP8FnGoy91a0Ggk7+2f+f3liEgz8wUue/L2cKst9bp
WA41WFim4tDdoCCSNoTNni0VoPwaAOY5tfHNWOACzrC4kpidznu7USrz5pgNsJBWKIj1FhwEXfLC
qpjIqKP3STUKS5r5EiYsxkw/C0xLvgT3teAKCbueFfpZiMJu037QWYp0v7WvIoB2M0IzhsIpoWI5
H1VK+aVyozwalNFu1d+BsDHn8LcBA8NlvqC6BqPDS1sMkw0nGt2ROaAB4T1bHHQYrceAszudX44E
vISApf0iEQBddWdLAZYmiTJsulhzCBeCmwas1hk6cmUu8LE2V40x0MCV57L3PZoXxiZJ+6FEw2ws
LrLLv4zCXq2uJlXf3vBIQDUjE+L26uhH3rQzuytyYww6kpM7IKfjTIF2LjuHRQjQPMsNFFUEVfZi
LbgT9UYLGfW7XkpJ1MzcK7aG4Nr/KzXOP0o3RQitEBjiKOZH1ZNT8/1zFqmog7eCjgyAX4HufZri
IfiogznRH3vmYeoQGlPqitAmkYSQOCJaYlIEPECMRKEpTSEjQwQ6oV3WZfwFg3iIf5z2REieRxbc
RZqepgCyDlrKTTlfMH02DSomq6pHQP/4M8U3QuUQf89GcvfvslJG7FeXnBmDsQPCVlaHh2w1Lzn4
aJ19ai4gIQPndB0OhHGpN/yfLkYusxLtZOCraXWVCBsuQ+RX7g+giYt8079Kai+vtXze9NZc93jy
KD57Ttueg3mad+PG4cz+jP4mYzpm80va0aYxHt3FgcVEAyJOAOqSOGThiwnC0BfxzT/miUD2iZ+/
7gEeJm4z4T3ddc7enoOSnLU43Voaa/lLTJEz7/pKqnDXH6x8+0V+lmAKMOEEHMHKYZ+rfUkVW4bX
W1CSpY9qZyTeqWvy6wUzAdxMYRQXfceYVkSnFWxCmU/eKTuds6HIYggDNNmij96RK+ficnaG8ECP
5/rx+Rls+3s/1mN93rGXMmQ+hzKrXV6VlUH2OA9oeO5DSwb7g7totqjxa51xmZ3uW6a1C0Zh8IID
KnzhLpT8k5s78jDsE1otuRAOW3xUVo9X7ByCjOUMr/StdNNOybFDmnL3nWn46RwjsaHUr5+pMYCb
IKWzkJR2b5p3zx3jFHs2GFQdJrfYIU6sjsJPsGLPJUPWVrRLYicIn5Bg19ayPhVo5e/w1NoQloE9
9KXTMgatHWR3XKeRDU80oUhMWzqZdAiW7e26xprWT1XOJcHVVTPNPm6PMEq0pqz1eIbLS7TN3jf6
XoXlw13cTCIZzjwEfDKUub7RBgQrQYdbsMnNRHRkm5LYr0QGY3FjhvcULtftxHmWMDnSgE9Q2FgX
0C8KbnWG1rVzFGQ6043CPh0L+30Y5S/uj30kpAkeeOj2dCSuO255ac4MnRHDF8x3ee2x8V/Ad/q/
htgVA2XSZ7g37CO3PMA27KBCO7g9BN0QcUIVlGeF2wr0xDBxqGmr4rhVf9WJORdLE0gd+bye1Fmh
8HoJMwgEoUI1c0ffzmGK03M8okqkXsqBCtSyloqxZLjXeBDWxdhSlRw1Jq3xXw46067Clg0WRQR3
3AQ+omce6h910zCTJtXOc8MCFB7xbRlmkKNjlTf1uC7kLGGanrQb4youc3BpRtC9PbU1H+C53rzv
qXBDt5r9aURFEVd46Iodb9HrzxeXd9bJaIwRf7lqw+Ot3x7xPHD1KnvljgBzVr/Mj43p1IQwBQ7f
tGew7M0NykzH5Uh9bLhQParuF7uTFnr1ozCTDb4xLCTyANrR7Wj+SqqePJa9V9SSTnv2QiM30sJx
qS8XFcESvcx8Gvp8pgWs6apbLAjF/BnQUG6kSCWA2fkfZ0jmKKmDNRrIU+M5uAbtZ43uti5ZALI+
CBWxTJRVn6IsZPkA1h2HLTg1ww/eJLvsr+t0boMuM16rsfa5kXkC5tmsI3glUOGZm1wFZBhIn8O/
QHhs78vxlM8SVmjX8N6mSGLTThzuMPJE9bfgkyJ2DYrv2qwFfdfEUbqPVqamr6OW9QEVzScdnj3Q
3ZIWswbB9KmE7LWLtxykUw6KWkwkotzeiu80NkM5ZaFNfT8dMpWNkGu4qwwrrLRrn3g52HtdIIWZ
rScSAp+UVsUnBw9z6C/MBtxl3CmPjA6jBv5uoM3aotAeGCzhPJW/uxoWvm/dapFnn0A8DuZC0pdv
SHYi38UZfxFuCldy1lxx1/t9MFnqH997Th2k8YjsrhLZAf7e5xH86i2QqGen+V47mTCIIRwqP5Dd
o6gpauVi/gXzE/vScuzrRq83wncrTdan28I8ebQNQStxupU+moy92/yU4wH86+oSmiHIRdI/RpYY
Sw63z8vhJ3yq3RNfy2MpEbhymDYpI7eOsdaG7wA7yN4XsZ980kkQSfctW22Lq8QjRnt/CLV66/wQ
U+ljsQY8+rRVZt9FZL6VIo+uJacfhTn4CJ6Zacq7jWEPKSJy0z0oQxqYEXSKcZFFMHzOEp1qCogo
jJzyo5wGmNbckGT2yoJIsF9uYMsHiUBxH4kLzBVIWVlySot8Bp3fkonYcvuonXcJgRYIZwZ9Xngn
jbHHVbTx1hwidYHAlt4Exl0EX0JXkFI2PV/8jsBqmen3wQIzzi0Os0Ny0/GFtkupmaDH+x1A3nxy
/iOLb8J2O+huQ5p4IRIu+ydCt8CRAnaQEdiXd5Xd4Ob7cOxDlxwk7HVFWsBoTR4GTyXC8MA5Ko1/
ktGG8Mj6vvE1nglzfGRJFsN0oN+bmFHyvOOk55H1C/S+IayG9U02ZoOzACYNXRN5UcPM9vH55ibs
exHqhyxn67GU36bA7em4l3DhL80uHzBrOYovw09P2cXoYifCSjyG1blnepsz5SumDThaGJHPh+6l
QnsBbbBw2QdwKRmPnyhSqFbvQ5W4U1HuHuW/jr+gMbty7WFA1EdkXeQIipoGA8dtt9OcyGBUWo8V
2x3HD9DuPMpGbFFYsaHeCcKdlFe4JIhWivnQelxDNFzbhTCQxLMQLOFZKQUgukiTcQJUdUo1j3D9
IW8g29aOCscPgi3LVg0WHmod8qK3bPq/IQnebbrzU259mzFI0fwcIChutu7ZfSc3z9E94LSdh61O
pohLYePxCn8/iazAGY/AArhuD9WnA6tgrM2csPxg9oTOrFU5Hv7DwXG/t3/LvxN/R5kxd/vW2znG
7D7bUD2avV6EdknUj4mN/ySvM2U244Q5ti6Kv4pMsVvAuHnsjzZzH9Ac4ovjB3AxFKCMG47exWWM
zHJFtE3ZPZzITLrnNFKN//W72PhyOSq2piDXCs51NV8NHeoah7uZ19leoEGH5n9uOJ3113QTlAOL
aTP0KID77yTOV+nPobaZIEyUgqMN5WXml9qAJdnwi9ZLkvYFvPYhKv/CaDzYKSdEqCAK5gTqxhzW
K6fcGcPh4Ye7iSt47xE6mkRjoKQhMdKaYx3oahNTaQjJhV/ZpNHeKaqZ5sWBSzUhVVss5a75gwBA
MzSHLPuoCfd6V16L23NVJPkXyadm3NU9JREcF/frJwisWouTZvxSPoHdKM+CmO7If5sqCAHUpKvl
LGko3Kva4xsZpCISuFwvI/ZurrvAc5c0pAKbYnJxR4YFXIC1CgrUXmCV+kJzCnJY55sLSd8pgO5K
33EfsNf0yoVTI7+r95QoDKroVcquiB1Q2w0ZB11xpOwIiG5TYX8iquLSRIqQr+DbU6JIaYfK7upU
b5qX1NiTRi42N2qRF5UO2vkGigDTb52SuHxzsbd4oEaWAgzBq71OoUYPnK7exe/mybfyFj3bgZYQ
V9fncTqwbhT8HUdmRsFFQzjDFf9dS9rkf4QgaR8AZm7o7AW3irwc24ynxuM6n0ZB0t19I3f5yZen
FsFgqxhEVKtZKq4H371gIDqDT+z+UX3WMSS03rjCxwwvls85OFnPAGvkgqdrEAteM0TK8tZ7DBCQ
bI4yqfA+o4Jo0zD8lt/3T1zLLtxO7tNZrI4YXUQ0L36OyP8V4ejtnCspYpKndkViYztlett9FRmJ
LEUhGjm3j11L0nwfuBksYLH3q286Pn4psX7YvvySgZgkYF9/TLlm1tvAlLptdSYYFscZNEfxiiVG
uhBPy6stYTjFUAsC1b8Lm00eFG917tpxmx4m524BKcLZS05ZrU/wYM0ijtms52R9qpBk1lAZjPCV
eVcw3ymh3TqNmVYOb4GhTpeHu+tW/Ou80I1UOID4AXEWKJ1SSQFzD3cE3+AN4JN9dDlqsZcrLlGy
0vU429hBTC+NTQyg/Ej9+GiNBgxgSHfeyjtoGTdTzWfexKmG2tWU8+z3ju3H0707dAbc+ua+DBYQ
MESBEnokHH+JXyebhCsXQ8gXrXBbjFgzfXw08acAJP3wFiQxC/FZG8pp3enkYNinIdnQ2It2WFYv
jx3JweulhSMDMj9Bs+oj/9LUrRvXkhPNaWCC4orirr7wR+Tc/eLTfKs1L3KisCtspAZ9XpK2muAV
d+UCOaEavHAcTWdCItUErggVOfMYdJ5NE0KDAomnq0eLrF+DkAbgu3P1YAW8V/9TJ+AlUrnHpznF
th4u92IT5XcK+DDj7rRUxBXsCpbYuK/qXCsF7f4HwxxxQPHfj6simRZ++NYHinf8sHQONMFl/fPb
lz9AWfg1/ENKMGsmF38rz/Einahvh6m0vnFfqyD0YB0LcrJErEtqa7h+5uoI4en9e+w1foM2Z0xA
ONxb/48+ytqrJC62lk4Dkkvf4EOeC0jeOZZKRuI6Jdqjm9ODmpqy+/Q92EjC6DmirwDVUYB4vayb
KB3qn7RGvbLpIFZMggKDNs8KeE3kWKJtSix0m+b9QKAEiwRqTl/e0CqINElOvW2JyEpFHVfm/udE
0+NEmNcDSZrdUkndxJZ70KD9PVVEugJp5BQkyQGo7BqkXS3YhxudyNQOYn7QIlouOUT0ECUSw2Ed
GK87C5loe7yqkZslYaBdQ0Q3DHqLkX3BiCjcuqzx4Y3SHPxi2n/nVG0xDoePHfx798wmmAs6Gvv1
DoZDvY4I+ymTuYIAyFQgGW9pZUkNPfWM2E6/ssXXhz7MuLLnNDstBrJWkQA6kg0RsHTyZbG2xOje
0NgsDwJ38KR5EIhm3lni8Z4hGcsSoMF5hXLZK4W14pI4khjxntOoW8wPoN8DgqctV98h3c7sB6ea
xrUzhZ2nXs8el88fel1P4A2I315tMJaiIN9pczfWnAhRQJVcgIa5qQaWBt78EeBcbNNph32lneYR
JynV37zsvbcZ99nzOXIgR2KvKBXrOR5LWS9sDw3vbuvT+lvdtCnXHkOmmpZYG+ay0FtSocXDYYgR
fOAnxDHwi+DtUtSmaLBZZMbERPjPaL19mLSHVUfkk2+3tfwWCb7A/v4bwNt9fRFZiM6C6/c6x0na
acXxRjepGTGUrlxRhxM6YLRxUkBLqKinxSwvYRrSkMZQbe0T02WQs0vymwCm9fK8k1zVWqjG67n7
CnUb3RW0OBdfqBh+lKs/uKAyPaBxTPrqlQOOSvuxpLOeaOtmMLYyexHVbQOi4SCOpXJEakbOBinT
3XbfuJ6auuRL3RcpKBqUkrT9mb7nkqCkd5dOENCiCorJiOp361XXImOZlpIzuFiUTjmcveGe4r3i
6DiSwQTRXMCaYIjp0K/KWRCH52DfwcMoOboFACypbre4WNbjXNkuMjt7SPNXzlHSARUOoRutbcMp
iP2mNubqi2fCVVS+w5q9Lwc8SLqKhFUnn9AvxNVPK0V1QgNhsbT+8JHhLPOsLYALFECAvBCda8/z
G3XkOO2gGyE6VJX/lQ5Hx1Ai6XnXMD4FIpd8uo8oxEk7A3TWnkN1v440tMcEEvD7Q+hIvuvwfeCk
al+xn3v89T8Yy+pkbsf+tzvp/MJQdDM8UkE3ybjOu5lwK00fGcp0lMQ0NLfEus+vIo8GW8s6b2Bp
6Vst6JnPhjjpLNlDzQrZtZJC8bnYPhpCbjpY9rggzKp9az28PVFCLxtVHTFF5PM7UuEjJ8cOio1N
JgBNOEZ0hHBvNVfRjH8IKUlXnrj8UPQESkqYBkIHp0Apgprm1hjS4gfXC+Iu4O93pnNIoYy51m4X
TnUgwyMX509U3IDBI25ExFGT5/G7QGQSDrHlsnUqF480kaK72RiaSaUkzCaazm71dW5WukSdvN/H
oYA8D6ZUhGOJBt+05ALU0lMo7D62CLytrdrz9+g1J63HDkMNgES3JYIg+O7bGHmwuKUBll3coYGb
nkBQTuFYg4xJtYf+JnRJgxxRTVbWCdW1/GfQ4hn1s8s7BlNEbE9nw+7vBCPts3xG2CuJVfwojtSl
0kB/9IGsmuShxuPZBlNuB27aqTLo+bbe/27dazULgPOhDF05+QjGpsFyyRbYSJZwhQ32+uIOOwYB
BBC8WGSw0JmpHGL3Wayn+D8alANR6Scm1h7XR67uGjgrN/jZWSbn7jsMVFJbeNj77jy6XOkJtcq6
48Xu/4TBcMXtUhY43Ka8VoB9FFcdR70291VQdWjunqdyoTZbl+MZsYekJSJGfUmN7V5O3EHNL++e
zGEtVoQlbMKLfdoeu/oaQG8fhL9j8bFGGRumITJAQgKgDciivdPrx/7+9ixs00f3lB9zNQ2HRyph
EsUf3w5DpEqgaM9RbFzOoGL1Kwp7uzo0rD46jOZl2Emvq20Tbr7ezc+DKq/EJfa+E+OtmFyVsXK2
8uHfdhcR8TFKFiv05QfW64ciqCzpGNJfUug7CVW/tJRwqg3hlgOcz5EnSJ8vN6RIGebgOuhLkBSM
fCvvuZc2WKlDZUkI0xrYbKaszMyxeHlRoMNgftnN42HnHzGZOjKr8TJ6tMT6/hbYxuJ21yDa8azB
0oxirfJBRTGVh0NrKq++GZ+BPJrtN7IWGRty8hzTIiVTMx4bwDExyaVJH/cCSFILjHlWCoHfaNji
+SYsKGLyQvylcXpDRTC30Eg/J9pqRqzjacL6aNSvkceJ8Ac6PMC6Ddy/AgTLk9A017gwsNDESe1i
3eQWYZDhLZadxTSS+3m0PcKOL5AVTuUlohgBJ/JWYRT3CwmgH0OSVlEqDMD0Gte1V7Dif2i9J6sX
wXjivWDDZD3GMDb3Jw1WeZrx9bBC8Zcm541Sdqvoc8w6K3Ejyu/E1kzRwiexfRhqAbqM20socF7W
oMT+0d/+8uC2O88ULBtpcKQPXJMp+xbemYNC64Tp67Wv/KrE/+eb8+qNc58zv6UTIoZugNFXSAta
16w03TmEt7re0JGK5S0ChiaSQb1E+tLekOcvnDde8L1o7KFw9VrTRhGHmu3g1GeNTId7ZhJj514j
uX5aCXVj6QyGrnm/eM49qoEaLN2fvk35Wolp6tm71neYPq4mCETCRdfS267LH8+mQEG+GY2Gs7B7
LU1zx+kYa2+RcDePhDo9QSygCjHdkENpVatw1ez3hoZ4KvOnHbMOPlxZZHDYKesuD/FG3+giveKJ
tQ8hX6alkcstgI5HXd+XjD9FaibavjmUtkb0NE5xfYfIsr5nGdyGWYId/7AFYj67MBmRj2RjqWJb
sy6COMsHucXwUk+q452nm8PWBWyXYBTcG83dQIFoO0yM7NKnRPWAclHanHLAN7PDQXSwmF1B18LL
MfXUzyUStyv7wPdL2cr/4SyLTy7cwn5PTTWVdGxaWQzMJ+1VWe4JbXSJfhCaFigxlHXi0LnubjFX
wG7d1gHiMEsGvPWVSPwT1YNmDeJMpX43nGOKSi/afJnBgoRlR9DsbcPw07BMKlT9e607DiTsIMbZ
Pc99Ozg6H/n0rHjHkoNH5WYus6cs/+an7QsJvp7e/6pgTBk4HMgLJup5pw4uaidMPOZzRwgLOlFr
7zDCqrqrghSdfpWMHO9gxYVInCbAuMEd9PG6a39yEZFzeVQkjEl6jK06E5Jr/o9dmWZQHXAYWBNw
ZnBXEy81LQz6y0I7MnHg5jPSrX0KVqxASJMqi+0HlEVlNiJD9wCtnyd8HEWNvgqtfr8vTuTbp7SZ
I/r3XjXjGDrlIGAN67O9ndWvZnATJJKzFAdsrGAsNbjiQdHKhI7g0erlVBmowHl30jZ3xKmExp7c
AGQXGfsxLDhTDBzCKA1TuDPH46qZjv2wszqvKkPibCCuxVV6CxVNNQgeIs4g4yRGKeYiVDJjmyRz
qN5mpAwZ0CWQiJbKG/xNoI/U0HMv1CQUaXSnzFz9f6qLQ16OxVZrn5pGPSfL2B6DToKKVrmEJ13a
tKiPMdaXgYB+SW9UqpuEz0YxwrUw5geQmSX8CtJ0vrVvAr/QWRpCJx7GtKtOtdZQkPUDZzJLwqEm
lIOHHmstfV4P8AcH+mC5XMew3CKAY29WfvriUczh5cohLeKJGobUFvb5+3ILtf7nFidlYiz17c8R
fA8Hoj0+/n8xy/BjGhbQQmN3vbcv+9G5qm0AZ/me6XZhRTNUWFXv+5/XVwdltD4nYoEUEeyljCMl
T/9av11d1I3pfotOxPTJyzNNh7zBurGCE6AD+AmxULEf8AOvOPrJRGAUiVcGztyTy1/e0v7MdpSG
mNWFXG4/Fytf+cRKr3k6V26WJZnxJUN1LqEKBRKDYV6BBZJZb0l90C6dGCO4eW8SDq34z6KZdcCG
Nkw5IDI6C/d9CCo/Oe9DIMmevaNZYcDa3NYdCdxcbPayCKJQyGdqRJzkoTwACIoWjzxLFNhCQmyR
wzK0SLh/23B8DtrtKxRGQ8iSHVtOBnGjVihXvi2ZL2K/JJYd9oHSC73yxiHCzU03qVRzyxqSRciC
L+56aIG4lH0Kc5dVwEAXuDvatYqSgR4C4dUlIsi7hRa0HNIZnx+V6GvuX2yN6IodFYUtczZZyNKe
lrvnRwx3fxqMDFvssGMlbEjmPW7qbZMujEnZF3Dmph2J2DaT6ZB3eZ/GPWtAhPFOJVlMdR9vWYgt
AE8bqxddmC7gwj+Rz4FNXyjdLgqd9M8aoP7UM7WCIs1QVQDGKxKJtFZ4S0MobgXqH3fv+1qRgYJq
+gi5UMPCRefpaoPd/jUgb5YFn83NYMsTeLLrql4ihSMgDqwWRPHvi/AyQA3wL5EXDayt89UtEUT6
tKoUx1Jv3JvS9cy66/dHVxUTEV0NjFS9luuF4fpEgs+VYhbPrxs/qYRCxaizpr9TFqannKebtFfo
vAdXnb0a2k491iGpmunSs2hIXdq2YfRHjFBIVIOvveltdyvS1ScJA62JLGK75PWriCCSbpPVdkhl
lTOxs+MtYo99oZSgP5pKwpxFTRGYQSKNyahLUVthp9G8yyouaZdwHt91lkuGFgN4fj9ztpMEmPx4
xa/4O/aPZ67KE8Uh6pKodH4SXIZSwwUJDx2yERTw7FLGKIGD8JdeBQrIsSYvgxU60GlXrO9CPsIk
GjT3rvJMtaSB8gQA8UqsRtJf/WlMC2bo4JqLMazKrT9vBSt+hbvgOqwHyeHTkvUVpEWOsf12D0VS
XPmtcYJAjN8P6mT02gFVOjFIvWK7n7DkCMhLNTk25iScOjuUY4/L7Z7RCTbasWdQENM5UaYYB2Jv
8rHtOjvxwHZ9W0pVgBqnzzCyWoO3HvqEuQeUA+L4LXuoocLp6HazxzZoD8d4dpBaewb8SsaA+gRl
nVDAaYlh6oCV7c/LHd2VU28Gp02qwSJMOTtsycjw7TjGrfbK+/ldNKfK08VSyPTP7o88MGQyJZpx
Wg32uuxBS41kpM7yjWY8R3XsCfwOYN11+E2vhstBk0go7r2g+xScwrMvf/l/5JVBKOZZzGnWJeTO
sYbTe2qKrR73EabWLmhXp2qX/MuZ+7on11kFJJKvfFAOYxYeVHaHQr4czLmQIWYIaM1chT/4wBaX
NcpOI9vJBX5x/q1JZnLrTiFWakAkWAsPjIcrvnVDcrzJO77EobBXUoU79JGrJprJsR5aws9ltkXl
/+BBn9aY81K6mAkl60W6u/W/avQQBWu6Pcw0DLNe6qCwH9RPePtOASuzW2IKAU89mnLxSPlVWUhI
wdPpTYgV5CTLwqF8qcFkQYCBSPvx7QZZhSiGiDBMLTU6Txyt56j6nWTI9aRHTtHCdJgG4dJo9CsB
AESgD7i2NscjnJO0v/MvbFnLgH0pJ8yBvoF91ZwY9LA6FxLRlxf8CcjfEIBp3BFdg1nwSh1Kg/2Q
m7DsctL7I+18y3JpZpNANw0Mnu5QVAWV7DIuBbw5Lkyhq/5hxAVT+sM9JXs2Pq1TMDMxzqOrwCkm
1LsPyDVsVw0UUHvdhzPn1EfqrG35kofMuMQb1AkKrFl4CeGPGwQprtKV6oOhObc94qdGX67imer5
vMohmdupPaD5jKAeVG01lKnBsEQTrG6j+NzgOacQks3yjga3HMFQvCmDJC7HtbdQKg3Doyvr/a6Y
p20jO4OOTiVAEvcWyarqClBQeEN0WjYXui+MgAh8IljPUaG4WUu36WmhdgaFyWNGFPLSEBQIpxDW
S9ZH3fHJkSDtOXM/Mmft+LxRm07m/odSzgg9ouLXcqqKVToVv2/ac1+OC0UK/fU7pafC73NvQN4i
1uiBBuqgXFuK+/vTdsrS8ZWN5TO4AJ5F1/DleXR/OuPpJbHT6/3HLDesz5LziK2rRtqt5ukpPCu7
FWlXF4Xx3T659TWJ37h+V+ejA76FNpJkniyhfiOEwbjbbW8IH25ZJl8sxpAaale0g0zBbHHZbC33
dY+ApqoOBwI30QJWywOKzjQYElSqpyUKx5Vc2rgPBZ4CBEb0pMxhkkuV49t6SEKzFEpSPwVgVlMa
j/4yOM/N2GedgKGOSP1A3QCNW9opNPNLKI8Fjzk7zMi0ALhJyR/CiL+rYJ96pIL7eKhlQyDdLU/R
cjcRsiLfQ9D0nftNug8C9a+eQIBzEmF5ywjIeCnWMU8pJ/iBue+WosqQW+NYDlvQ4fuHy9DvevNM
dPrOub2NnmuUQl0TAw1pS2YnUGLvdGq13UJWNmcSIBUpO4sz33bkoKLeMFbBVrM8YiafA8C+G+LW
TGg2ryDRGyRCdtGhBxdlr69SD2THKuUoe5FC9iYQhzC1xDnyeR6y6KxudbvcPlQR4lVYd055110m
wj7uvpvsSOWS7enZGGDmELyl5TyM8DNhgosE1XsqkgzVafZrhjce+pw+rVPcdyW4xP1UGfZy5BK0
NSev27q+NcZHrMpnwKCz9YieoUUc9mVHnDhHVtAcWeqK/Tog9aGrEhCxtDnizqZHkpKZFsZ9220d
PST0QjCz8GWC6G7h6FnQRZe498vEbFR6fTgUvx0iXv4332hjZ49aiOJeKjR+VJlxU++HvaMFGNLE
xB9NuQjpZOGm/mrZM3MlCpXunKaPfojvViIj/HL/O2766gm3tBgb/Mi+iBrZMeTPhS9km6rzHwPE
14139Q+ctrnBlnSJkaoDhYgrsq0RYmXjxof1uT5T+367zkxS03hCfoVO0iorfAdIcC2eu2e8QzNC
qADNnyBm7gVrNBhTF4eRVighXPCqIcwL9BenuAEal6G5lWzs1kFYwcw/5Aey5KT1XiFQqr+b7Smt
1kAcRXSUjd6cEzx/axQJPZiQ83AGZ4IzUNzfcTYZvVrbZKy6C/sTGl5J4hreTo5DQoDf89YkbwH/
zNjC/HR8PVtr/U+9+8sgBSi3/SjkgmF/y/CMbyHsgKFwTfKAV0c7DnbQy+nQjSYiH1lKXm+sDTGR
gj82J254cHjZHH16gMVH54a+ASd0vIHGqb5zzYBwwuWSF6xVcTwVS4dn+7xcQ08K6jeTlCrEAVKV
DgvCu0Ppr4I925ANODu6G0vSvqVKDcmPUcq5JLTbW/LAkRzIhS4Zn3DpdWfzhKemVSmI1cYf+V6x
ovAiujuooQIjhDu1JOWASuN/eUun5GWsNM2S9Rnxb0Sj9WYNx5BNUf1BA4BQVRGN4r7Rg8tj7bHd
Wj/rc/RxDWcBvNNIY9fTCfismMAqqI4TqqLvVK6e5Zv09fty1rN1PyMw0LSHSS9ADKfZCHI+9RkU
Wt7dj6mWynGDl7FjIY2TY7aBW+4U21Ei5ox+IzxAhFwtcG3swX4902WgCJtfckr7nfjF+if6/tXU
AOFYy67JV6tGaxxFY8kMdQJvNKdwZrhcYFTuix8Dog3shp773Bw+KHFuOYfUeh8grOEYHvAmeS91
RwZOUDxz8KJe/CbWmr7IHfP8XCyHtRDn78BfnM2QaOaYg/eVbeIyBPXsb7MexS0Q4iJ+uguCibls
HpAbaSwsrLVy+yO3YO3sN7gYh9fEgsY6cnubsRrMWs9se0M8KHRujcUZ35eY5IOkw1tgFzoIx82x
3Wz9Zjk9nlijyPav3rB4z6OeJzbKOG6raDZFAG397xuuKsVZ2s+FDAE60ZXVqiK1VjY5VrfIfmlp
SIUkx8I1BY1t75m5qSe9bJcgHWYUP/AQz602xibGnGIzipO2IPcTGfMy8jNaBTZG44nzQSM6YdL/
pluGOVLhWrWXiWz3oC8N0NFHpJ7wqK6g2P1s8UjsEYZ78g4ECC5F80ULi8pEzrvfmgsVkfaaOzI5
3bvNmp8mpQo+Yn/wMtP8uLAn7pQHgyU6BDH/xAhtyiRuVlJvq6YVF/VGA+7SmC9IzPu8YfzDP9KW
7rD4Ttp40NWzzweve81JShGPklV1KHVrXtwp//GR2GsWrKtwNSQSgDgWJ8wvWu969D6tmsBvR6U1
9gKuVPTrfpx3fMcjkLkTTWQa9ybsmse/ssgzYbed3dfWXMzVu3eFrpspOpQ/CLIGxwwFPZbxsHVT
PA/5YquJyLk282DbLlmT2x5X0AVRg9UeJb7CE3w3gNHlyienf28JueXTSYSAd8lgVKKhrlZXpCMp
EHyKgAH43UYlpf/0M686bt+GD4npVkdLWsfBeiOhkMlU1LmuzFGl3eiei1Sj84878XAPDeTpmjdt
NxFE/7IWjIbIiFsyhRezBJ/URxrQ25dpoKXWtyTImhbWMjWK+K/Y1BEe5diTZaPkV6VeVLaglgZt
e2NYvBDW8yR1dDyutYeq5N2QQO5ICtVTIekvwFpOXDgoVj+Wkak/wjvu2a0XNWS7gZtGZaR4cHPd
njyS3fW/OngOID2XxrNFLJNhZqGv5zlcstv50MBzKWxxvVmJmjoY/vzuoZCcsgDGtcCVWFpWkVDz
U7xDgpOSebnBuzboII9GkUsPanFeIO14b//rJ2dfvRZ8+iHPyXfiAXZiLI+fgsPr1qE2fvyo4dZ7
fT70CT5/wh0WFGScaBLnsRAcGbwa6uwMB8hGJnLgk6eROgW9daKMtzmPLuYGCB+pTqRmX/qn4NMA
lEB41RZ6IoHTSGxukMUs1fsMv+PZQ7kgbPYaDXkAGYdQNlMffE1l+MHPfKJHSfaNTUleEZtt8IGK
0Mefk5SpYXxfTp4KsEOPjX56ECIYCW9zFKKf4nG6lBsIEIPKdGDZRQi4K1q5Y2oFxFmLnYfF0qIc
b2+DQgncFAc+tYNk8jjta3O4bn6JQxDNDZ0zOXbmScKTR4Z33LCBZKnjd+LwdJNiR4ehMb71JDaP
zBfaQmdAKIZBlKrt4V0kCo3VrZBwp2A4J0/nrNWDXGmYGhrY2tU0VKLwj51ZaB2BBS+oIEEGn8qW
1zj2ox4bWfy3R2ArPMWk0k5GcqUmWoD6OBJWX4FvJRFvSeALvtlmX2Nc4zEUmWO7rcinrwySb459
XbcR+vE6QTlikvCXbNRxVfRhEBzbf8pmMHHS7/Wsj4YJijyaedlUb6x4rUq0OqSc4+f71e1UGooQ
/At6s8CNzXwPmoau588Mq2i+JEuYuZLiZekl82gLsYYm5lNCe40lP3Uli2NK79lrnFZnLM3QNSu+
bDEtz6CoSMOZiPkhH0Ca6asqau4vNJbau2sRyj0UMKQ8j5D8vvfSFU1e1Nos6hfwy0ucL7EFiS6D
05lVbFTZAp3f9p3rY6aXExqHewU2wkv7Uukn+J9XyNKsA80Zt6h3538RxhYK63O2RxcYsoYDWlGP
HBkwAYK39QAE/07S4PyQ5LUSeBDLgXBjmtDMj0iqUQaEZ+XW6PtyABf5JSjV9K4xs7CLGH9LeBfU
CaFP5TTNln5jbMEvkUNIZYV51v/gSqccNf4TiR7BVN7WRU8jC/pvwjChrG6sqvZdmFyrMBibLi1L
XZOZ5S+uW2ZG3fEmW5CvQ7pgcuCszGGRA0yhx+FFx07TZ6N7s2vBdZ7nelbTS1WGP9ShBaqsnuIw
AELkPYukHo+gizCSM00CeEJTC8UTckgIBA3ja+S107sp/guGXbZSTMNwtOtWRNPmgRs+dv8xwe8J
46tS1gyb6wxBpVpm94qnRLUxTdIxSSCrO14yO05e972XCJC19Yc5NswQsem25rIInL7khEgBTmzv
av8gQ9NvqJxbVq+Bya7TxFgH2MEuo+mo3mTGaBKFX9Cr0AQPcIHXbg2Sl6Faag1kjMwHVM2uZhva
Qde/GsTpN68M31oUUVRYIxMtqYzjFf5SMUu7SACxuq5AMfCw8Q9ua6akaeuGxTkTcAwCjPQloS46
dUMZJ96zcclh3gBgKBisMUp9BFkEW+qIiisAKVCTLXCwY2tn2+fYLLXNQcvHcIEvpfeUt8FB7dml
rw1zEabFvI03WFQxBcNKjw5plP5JPaKSFWT0MbVff8xi7H8Budzil+AfE3f6AhBZ3zJ8IIj0CJ3e
+X2Ce5f4GAexDc5pkinPBfsnnvTtCe7pxtiyhgFHf+r0RkLIPjqS+FruBtO7kIrcCPBWELDyEj2l
PbXvQe8J5/uGhhASGNlUArkud2tsiLRuQuK3axuRe8XYOLiQw/rOK0MIh7vqySy0ExLzeWOjDfYQ
m8+dml7Wo/UzJNPFo5eqUTgXLxwx6exXKhzTMpqPgkuVpr0/htpairlkVcuXpQvvfFlnHGUBrS2K
CBxI+BEb+F00nuuc2in3BcSCVxZ6f9HtuB92zhGSX7WIuBl/9z/oYsEH69+EFTpEFWU0EI/mbGJw
60bN+/Gz0FLHndUZJHbF63oSt6S9dUjKJq7jfTNp7BcfNgXb858wxto8wdeJoA0PMQmmdgxUPwTW
cOGI8dVsD8pASUMV687XdovxiSTzRUufHcBOrTJy+0NMgfc7VUT2uMFcHsUJkUCut37JFrLNU6vK
80bgrJNR0rKVPPrQlXqduxF9hNnRM9/wZJr0zwSG4XRYgC0c8NIGlgJE5DGkgi4DWQT737q3drBf
onH+wb3g5+brVo8KZ67aqey84c/6bRkkONYOZRsILs2gnthYEUFV27uteWS0nJJz+Hy1INISuQE5
XZCaxiyqKFl1A5tzHB+0y6pqoaR9ZnqDwFik1veTJbtek7pDsBQw77g+h16g9ahExmdVKflFeczz
0Qzzh0ufV+e60uHI+gXbgfv/c2LrFug7sAxXBa5nt2WSzsu7GDxwSFs7zpWVQHTALFPwLq3/NJjQ
7yEUnFFpJkvqlQNR3/+Cf0T4gX7rjfEy9vfbXJNDdw6xN2c594Q99EVOfLb+gS/UQDPrxnM8mfV4
mG/moTL0OvuUjXIBxN/aetOsZEnXsFDRTp1s194bWbS850j6JzidrB3Ld1dYBet29JX9hM6G8jiI
ppuzQunOw5aEXS7AkBayVSmpTF5bQ+IB9xaD+7hEs2m33T4MwGmOO/oDW1ZoNcefseK5NFMZH2EC
x9139z6YptrzLhGd22mIObru0UXhHmYhpasLGG6X/QaPkhbd+AHb7xs1WHqnc6YbxT8xRI2AiDsB
b1CAiE0iNfzbGWKvXcUJ8wduli3+JB2ya5rmEhEJ26Rg0FV6vZt25JMXEcEtDu6xUi2sZP0ybgPM
5FwbBhK7U2dmHJfKyzhLsz8cv3YLrU9QIhWVATWxzqIVnwOQjWIZEn9vIenOsHrOFlM/5nC2O1OB
AMo7Jxqh7lVOAcwkss/lEQrBoh0wsy4di88TXaSBjbdThJoX2TKU0DHDjkpOeJIIVp/Q2I/CblNi
qemQ5uxW7yjvJDHALxCsovNLQ9/+Ll0Tu6BQCJ9v4o0o09No9JSa5WGmSQv01fb0XMX2BW1EbMEk
tItnuJ2YKirTUT49Yr1HkjIomVHqsbnUDynIXVStzRj9igJSSrdfR2gju9XMNs98WPzKR3fvZqMk
D1lP9ly0JSQsJmnQS3d75l4LnlI4IKG5d9d8uKQOOoya6vtbwO9i+Fa4BX8fgh0Vt7EmxsSi1dok
jtWidMG7uXRugBdXb8VxH/R2ITAYxdiM6h6XGnQa5SgbXiidTjX4NmI+yqal95gG6QBRJ5F80HSJ
yi+mim3G0GWRO4vQeFfXtFjB23URrpgRFBEifmhAIXBDueOfJWB7u2DcHmK7oaLgWcw7q6dcWlBF
XNCQF3bd5S8uT6BCelO4qejkLKgJ2nvHiahldqjtx7GhL6aBh6pi2i56ngI3k7WzQKy+0T45cpF7
jcH2XD/aR6JBYn8kPhqdSuVlixS9DizUdLQ4mhBEgW1APRj8KJT4OAL6FkaZP9RxTaNlGG/7TKmx
R3M9Xfdri8sqoYYfPFY37d4d04eAV8e4s++lfpZT1Jdtlzq1aEoQfHPT8QdyxW8N+5UUnj2R75KM
2bduCe8cZWfkoszz+vnWJo1dGGzz/S0Fc6bZVTKPsX3SiJ8NdqbaCcxLdM3PVj6kLdi1cVRjMmJU
BMRHkmR5ogmrTkToLf7KO+S4WFAk8l2o3j7FSGnR/iUldkIIgeObR/FNA31lO+6hpqu7IMIH7G4/
TbV+81vjcXYUXWrsa8QNX4tGE0HYWC4CzFQq4Z5aO9t+emkwce4oiCqUv9NQeoo32ErSGgkfhmpn
b41W/Pu9N9fTtYjxrWzZaG8jpmWam34BEdKcLEwdSrPecZlP9ulkF1p70v4JS8apzLMxOPRkC4f3
u67qDYYXLRx+9C5cNb7kxtyuifVJ4OyF+urewoPRvC3c1axpYta+emPJcgW0TEcLFNAq7+HaE6dU
4WICNklp2++4w9lgVeyYOQnCzaBXyh3J5RbcvHZbcBR9QNPzYhUKS8dV1vvyyJv6jq4dgcBMDJ50
ZTF3oNhUxo4IG7DuZNvXXv0TtruiSH0Soz5u+R9ZS7JJ6rXsdsnWuLaVvZ4BEI8gFuOiM8+lcQ1T
eazaG9EbDVv1d5+OfDo8M/7AXyJrZuWl4OosXU//wOvwUDE2AV1O6BfiAh0dERJAdwrkrSHlwrbV
Na1ZhxkJU9bKH2w7oTIPIz188jExwV3z0cDNP4+fL1QOlx5r0/3RszqJ+w6XAhigE5zVCBrlUz6o
lcMRYgOnSlNQHtuYEOOeQLco51HzPzbnh4fSIOSWeGgd8vCc5777D22wAYxbYW1TAjVqz3tI3JxA
BUQyx+2ZrCmMwubF4QXMGemcTzq7ErkgYuMImZ9Vu8El1LCkZwBZtPHltwPtBNP5QnIUBwM5ATG5
7tGmgFLJU0qG969qHOh/8OCehqWmbV8QoqPE5hR2HiqKXeqgvxtY2Q41vXVoCEbRQW4BqFLi7Yl2
GLQcS6v5bTf2cEbybfe2br41VohIdVibE3QBNxFnASjsb+PSn45qahTzDRjV4nGNQ6GC8407DWj/
F3X4u4C9A+lsZB58MUn4gYnU0MbMYjmKAIDHw4Xv73/LWCp4Tk8c+OiYR55ELpfNeYFKx1fCl7Ig
XmPWkFjdbCR00LiEsYJajBqIoz+xdE/OBIG3HpmbsXuew/1lxAvYMLMYCc2AhDhqSNfgtQh6kYW1
nml2swzU802uBd6qVd3CeStoj/kzDpwNtJcNmgHGc0qmH/4io4S5eQQC/GhviXNBcJD5OQL6IoPL
B+6colZ+hiQnvMvGYxXef/etvXzGqMpzeZ1/43Atn9FvJGX2yfhgA1z7O6RakrizoSfC2krD/qIr
Tnn1BGPG7/XIrgJ5o7Q1HlL9wGFbyF94btt5w8qm6xrcU6RO+/UcZOYENwlTjVrYih/8cIsd9kEM
1KuMb5YcR09aWZP0Fx0lfwh0Z8ZSnzKS0YqNJU8BK78v9fzfUkfKa8671D/4XZ27hImn/3jVVJPI
AP4K9t+HWQvub6vNh/f5C1vbXWFulkKMSmNjKbvUh2wU7UtRRWyMUuR8QwcygwO/stkXOjy+mdP/
seMN9jnYS+mO3DJRxZ81R5Msc+kU/5sVh0dnproEuh2JBBAXSynvckBtz1UpmeVwhVoawhKwsYJM
YnAypKevmwSrah4Qjz+kZ1QzGeBD3QZ2+nsT23GUFA3vaAhOxOZT7sBENklRHMrKYhlVBnQCtSPU
bqbeaS7owoO3T6ZxdAbyuUdfSG4QZIRXBDuvh8LtM6s/s1KuCbEAsCUHIqx7RRrUQpfQKV9jVnjE
w3J2q+SyWvpzGIjKA3UphIaYRVzoRiPPqxunL0xCMdUt34iwLLdtO3obzqfgO73b0iCiv+xTwICn
1gpepABgLi76UbmLxd37pGO3OjoE+63xIUQ2cDxr8SCf4thmmOXzXW5GXlGj1JzROTu5tveQQYdk
05i/qaecZOiBeMpYut6z52Yq/oZCDJ97eg2pW7oA8TVXWrTTBNi3LCiQqTvPW7co3RIbBFM2SsSf
aUo4NqCJtOoxsLa9KSs2SyDU9Swf0DBXqVmBznEwvWl9i+Q8aQ0IxR/7wjTlNKcDb9n365cmB64i
QdQNPd3dSU6gAi8inThvr7DQDh2MOmw7fSHwo0HSdMDWCHWOfFuD1XDDc1AZiYJzjrYjikX8XFR0
AElAf53FARJh60IG9OyXWP+geg+Lr95DJG4Q8V75kTbRPIXWnSq+HS6RGH3TJsHXHJYygtypqPNn
58Tph6hPW1InKP+kpp9URtTNOVBTZXOCAX5p40I7Q+A9NCdHUwbiRZHy0dn8vnsSUJ/G5Oswbyd1
xuLiZbV5Hy1RSmzxKYZ8D4aE+IMYPPuEky4QVz1IaLQMxxa5Fzr1z1Dt5beB1xdV7fG00+DHYI5L
IB7Ft5wUqHTTRbpxbrZs//sMzDn8JQhbW+t+9bxQ0bMajsCBtm5vr4bHbytS/vrP9b4LE8WvioZK
0/jxyOtYr4cVUzPfMs80V0dQsEpQAaqLgAMVFcg2zP4ut8S3aePsGzEeDTDa1SplxvWEyWruOU1r
/PecX9zDj2CmQYzMZ36EXApq3p2vnhdAHpl1mVRs3lzyibAnLJ+hOGDqCpbmQdoX5L5clG+qbyoZ
71TDe35J82BXAIdXDYH4ghcsxztz71y6O11hC6L+7opt4YOOhSXm6V14wogofbf06dSgWXm0UZ17
rD3Wlt94sDmEMiQcwDNKnYDgBKPNh+SapkGsifa/LJ7ertAo1uJA6sT6bIYltQxn+xjjwvoEaNv9
wcb+yTzBLbtE717XXDXBiVsNNrcv+zUnJHQgjdyKGGHhM+CqYZ/b4+F+aZCSxpCOfXyYOD+ZhSqJ
md1moArhJdE2bxOVOUqfe0zUt+W/bsh7xTl6S84tJA4IOgAr9IpwpcPsKoTqSOScDEz3wuRMnUHR
8rViXQixsuWX65Ru0zNf++//ZDK/f9tNEVZ6DfR7IsOx9LJfoByuqfcwB66z41bdNbx5X0fn+/xZ
rEnzd0rzC/jsKkt7GHpNejZ06ACzrT6ZOOBPWlcUiQdMDI8LfhjufnpfQ3GwyBXZ5jAH4p5AYroC
8L1c8pcHVYLvzxi5L4IPHT7MbZAZ3WkGW3P1y5/Jqwo6H+S0u8Jrcp0tHZ0RsQUNDiTI14n1qeSD
odQrFGXEVEP8SqjdO3lirDuIyv+uMglW5ox4lvYM8Z866GxTa1D+4iuBF6XHTmueDwI9xVlPEkqc
83HVPZZKgJGg3pbe9VQcmpKDlh7nZJ/WBunEBIGZoznklIUOAhQuWco823917o/m7lmqTmniPQxU
C0kvmK8n6RSLdCd5N+CdIVvXL7FJ5kX60Vus3xWIbbvS4iDlpqlEnY6DhNxXQGmMnaqhmV5Y/l11
qjnxlbfjBdOcUVrXmWf+6fXAVh0sLXzYEda4pS6Nx17EWxV5CPldJPo7lgozcq07VFcAa//jJea3
1PbevaIQiWBdIGktldGXBA3VT0q5/YyxO5dEhLgRNDEwuVHzS2qhUBGDsDDppCfi/dpY734G3Flt
Pt1OegFDvGLTglLA7gLFiffRLK3f4FmkDsccPvXhtlLSp3T7GDOROC8SVzz3XgjNsMhDP2FqYSMM
Cj6tAoVsRoRCYCvx/jCSlSrlL/HRUqZCNqaAHRrG1k/f7KTca32jTmn5rNa8ifmTu0n1vR/oeAbl
GnUF8IyxQ/QtIi9XYSN2ymQNXzGnZQjKYMGsk4qamS+c1ZlJuztgaxi7bSt3cOEPfg+p26HwxzMs
agHwpxaRN2i+gO4wreCtfg+SdZi/xpg7cfoNXUqfnd5NudPoJmbzaHYNbaRgx9G9lL/B6XD7Fm3m
5OhEaXFvr3T8kzzmORrJcbeemEw7tlie+E/s/h0INhKGehL+EuMTCeyCEqxQMmbxuXAmkz+gyTsH
SQL5kVz+CVJofsWLuUV/ZHwlO6SL2v/HmCAp/k2oOPibOPAN4nRaWOESyxFY66HWoUnS96J7dUYM
he4hMYUYSTxNs/qpDVOAwTwYZE8+yF7tGJgOUzdWq0wbYBzhUFz3v+XqmFlwL1wAHM5Hpyie+Hfy
CUUF8iTGU1wW/iXySist7HEd/sUAMYTpibtfBRg9SFY+3na7VGvIIKJs/cgLM0QVl/DKbJbZpO98
DIu536hBT2VsCCszLd9b9TD2OGz0NLLl4+tlrTN0nXuuWXdLFZAhZ+6VFgzPeiSz/9Hj2fPC9BQX
j+SLzkhogfSYHkM+TC3ig9pCXyJguh6alh5bBSLTaOWpvuQH44S/s7u57ErqFDAcROhOObeGcSyh
3wbyttGAQ59ygOHZc/pZ/g9F+mAz29i+Ky2QemV2bSRbojNoy7Ccc3765CkyjkySBgCq43b1vWkt
VbFIvPTn40ZDRh4vfVrJTM9Iu5v0pb+c53IX/SsCqwhfP9al0zDiDzL+/KD4bXsL+8PPL9WNJrQD
cy7R3HSiuimxOCLs0dDiGykya/pvqQvdpEVKOhuryllj9CS3pu/8jbBmpPtCLRotGnM5sRFQXz8C
0TMjrSmVNe3IQLZtBgU9dL5diReDUzbanWECSsI0y7/Obi+tXDFiBRXcziswLsAA5k1vGBMNQODa
UBsvCW74ePGffGep3mDrJFj0lJPH2xbIAzt4VcDHGoXW41snczzCZTX+qVxGWcmHyHwDEXz7kKh4
/qfl+dowJOTRffs0V/a3r+iwnVvON3UyZh7Xygm6c9AJ4ErCf6ilhassQuW+CcMVl05wdsDlMGue
GQQZlVuRkLzk7y17aMd1IkcfJMval1wmtWv0+Ou5DP/g6QQ+I8NLaZ/eSg5u3nO7CvWN+Rh7pvDj
0BVpJ7CjYIm4MHhTppIFHdXR3+w0JD3je2/P+XjoJ/6RPyhhmGtvEY+mAxgpSfbBhdBVAD1FkMVE
lm+pRh0tGVFpRR3aiQnHz0d1rjzmukRiQEw3dmGgPKTTs7s/jmVIZw7Hble4DPE1ihKEddfmwc8R
QfcK6wVSvy1o9LkcsgvcNukCjJJPy63WgzNJ18ghDIcbB4A4HA4H7NtPLG17sqtcIvYR93k4AILF
mRIyq+E2tMsGWjlG+UjYSJBHXZuvMfeiB8Lh/SDoUJe8axu3QbXL+aMzV8kOD55JEkjcoqOQkBhr
LYjQqPYZC/XVCSwcHrT8SKGkQCvfbY+T3e90VV/NxsK5sMD0pOIUULVe2BfJjBA+jjQOmCoBRJp/
PfU0fTUxCBKXrAOjM0mV9/s/rPNILk0aj3LSQlVBkkbhlgKu1Fh0991zXECJsEwTkqerdrT3/0u6
31LC1xdBpZ/65rxDNhog8V9kisls/NOt2oOMUGm4By4Wvg8/+dz4ULeVS7LJTpVUeYhd5sWQcoYb
3tCumIvBoQlu8X2XvRaGcxbTYsMcZRSkodtxuShW13NQoTAUs8XCEojNydtyWwiYKEQPdd1cf3db
IpvHOQnxnXyunTN6WAV33xQZMBopsV5MqiuejhTVT5B+KjoVzrL5ftEpSHcYFsHzY320wzPU0zXv
JqT4g/7lYJ4KQ5+9Qi2hPJKQaFeqNbEPvdn31WIrS4zlMt2bBvAnnCWn2wyGFRwFfekENe6sXhQ2
u0B+SSHzDGtg3zbaSWPTVLMD3OdQxrNT5cAfSpCa8EG1eaONy7rCmWww7YbtsKT/pdRX8Gxmry87
R3nsSQCkY7TzGAPnhOicpWvFMddbDLXhdUzPR5tbk6YSXJNMc1B6sFyUKBBVf5iCHCXIqlY6WWdu
1lgnNmeHcdU5puJ8s2EOo+I3nCQwWGw4WgIHwJetdQ0+kXZ8ZIvjHKbJxUOyyKzt6IbK9LBaXr5F
12VGdlSrXMNic4/pQBaJPvkco+/U9pHZJk55ThoLFRNbru2TXDd1Z3Xvqqb/nf4otQafyn5Q9mS/
4yXxjmdLdV+vOHN0/vdiJLGYp9QHqWO2dOZz9s/UQZTHSgg5nt2ub1XVjx5G5syC7aEBe5PQqXkV
YhFq88OR40lH5kRg+rpzK82P7IXA+4/dlUKWcFvTc97VFn4rY/RpJroTz/38mNXLp8FqEZyI2qJN
ztQfyCeh4UV7HYY8Dr8mmPqjBGJ63WWhexasjuj9hbPmqhmiTUISP/LjZfrPcPDRTybOcIkOWoXa
bVMbhyLVXQYDC9d1mgOWzCDB1oNqEpif6TZ5jY2gfmEnHi/pEzjRB0Z0V70jPs//32t+lLi3GOk9
TO3skQfGsE+40rZ6UbFa7c05nhbP7KRLJxuN3IFjg0MMWwnahuO+XM0oEpbDNYgJ37yDmxcerIQn
VC6xvjg0tONOCIGwFq9jNHnki5dbZjE6rtWuPzdMLuxXZvltyhRL3PvhVOr9xhSwv1IQwr6yJcpw
ah3crG8oI5xS8u/gC6ZzUNfCaqBipApFD0azqlHKNhrUGKJJxW+NSYXCKajP/a77wlf6Hy9npZ32
AslVcwxHrOQVwUG4PQsfQX9dDXl3r55GN3WwUMJZ1lAdnhBWE/8viWlu/7dbDJ0K1AMe+WsmeSy2
65RdKf3pci/5dxUL1563LIKlxGSIA0O8s5eE5VA0ZeGsrTPalYs1UTeXGfMYBI8UoqLop4WntiNC
YFNBmPbvK8/R56I38ff7uVfxxnLs2VVKPWiyGCODAxz5rAAWdcEqfucy/QFfIa+EHA/KoSY8tkz2
KyYqsHKTBZx5TmuP8WBeoDSqjdxXn8XfZSc75BrXA6/yz90s8450Rd8juDN/d/zKK5lQiW2fDXvQ
PvEcC5wkWSjWpKdD1tCKSVyrk8yt6lAewj+tjDpuKeAWOWfJCHYCrZPArNmYhX6QqtGxwIBKRer7
4oJUT2mkBlraKFnaYqLCjxIdQZ+xBHrq4Bp9eKsjFJfJZMVWKZQcZ1Vb/kriOB20wHL7m54MJFv2
zFMMcS9Zbk5J8sLuWjxC0OGb1ziKKk2Fms1iCj3QZgVEEsbNnu1v2OVBAaK4PwI+9vs6MHJuAT0m
9wC6Vzqhmi1rxQujJqPHVWVr8p5KYLCXoBLLx761CC/aWqgNW5378dXxQ4gqWI/V5dagwWpmidXD
AY0VG57HNITS8hn21Stze0hXg57DOU8hpnZD43/BLo9Dk0lcAKZDpbI56vh14nUq+6Gji9ZdZMtg
vW55AB2FVukYUh3lsuCIQSMeh98jZqyoQzLkHv8ecA2ojoHAhDwR7jih4rnoKBZQRXluyX1BPlUi
WE5bnwX3sB1/NFNFbfr7TrXkWEqZ4qvkbYKqgq7RveJHoeWlCq+Kz0GOJEuaFtRE8NExbuja+eTz
RAcA6eGU81WbQR8rM051EVDGoP66HxCw5+wNIhJLebY3p//yq+59BMpoKOgsbZvL4tlJHStYvv5u
fqsyQt00mJKYCvYZQE/t/Wdv2Hk+NnrdpDt2up+kRSfWF223nJZzNvLybVjPRbJYO6BsJCbpyIWm
od38A6+pmNYJ1q7KfGpGar27rvnbCpsRKxjHQyEbqN/nBtiB44joUrRhk3BD5tqns7Xx0CsJMO1Q
MzzbK2vnZGBOxCwzBtug5UxIoYMTpsDntMUlrsIYgRbV2zoLgYk4O6NJhs7veYQ876los8TEvLcD
BinbGxKySFx6c8hY0D0o8aDsLLxp2FwrZieHzPe9Hhw5cxQd8oxmooHzSXoyFV1g1bLHFp94tsMp
JBf3O19T/3NoAAmgDSdd24XEtt340TquGS0MLFuYpKhOSJTutaYllFPWgQldi/ZI1JfVizANELOn
py1xjbOlvr9QgFDL/UJ2s671si0iGGNETcIbYVMCGtc1O1eZEtxJ1GhMnyimmOb/XsqU4R4Q3a3Z
qCUQ6k9bxKLWeALaVyBFfclF9TFWDMuDXWfmigAaFBT6cOBDLR8y6t6xeqAPVZSMnydkNpKL2xr0
iVw3DxEv8V81cV9GgY8dcqseVJUeS/3enOsxpjhYHZoCDR5h5j1PeyvsS3fmRf4K1DGbkC2gWlGN
ABv9g0k79b6RSz+fNyWWrpLmcwPpgA6UzKcDEFionzt1DduxVIabJwxn4TF2PjMTcIc45UlyaAMh
BWngxWAVAICMrdS2B+BDlKJuGlSNsjRPPZAabz/TCbV5wT94heBN+CmYAzOkIO9PP9fkdYeKs7D9
8JZg9fOkDbdKlnQTGi4Mp9iUwVTh6oyITt9hYy6cAON09g7SdVy++qCUe8yIHvNi1IraLbi0yi96
9IpfbMsRxhhYWUodmfEbG56I83BSFF7dLtT5hkjE5MA+Bm+EP+GYgaY3sshYe1yQGCTtauSZXL8m
Aph7NWVMnoeIAMynNOhTxg61NyIsiyXi/ED5+hkoDjWblMiuKNs8MOv2iQomiVMNU6+wJF1ZNMdN
MLi4AKffXP81Bzl5GZGXxYx2ldYAjg6jhFEstcLskDWhHYCfeDkrb6h/w1cd6Te/tYa8bMlO/lOU
nQsPqZAo5uVihG+U2aIkwqADymTONtO3NYzGABVRD1wh5hpXua6+NX+T0u5xu0ceYgyS6gZGPTwR
cupysHd7Wpn0zt49KTJNy/CX3N2QGYXj8ilJY93P/H7tta/Wjlnvzt9JIwzdkPID3zyFQss5vUhm
g0/+WD8RzKe7XhVB3ijwLOX6VgUS2tf0thEcod+iO1iKSDhzWJEOO/oYUVk3u/VN8ztCUV+2tFF4
C8mzwKSTgWEcSA5fhUJIq0ceQdMq0634e2kYbvZN1X/zwaSJkTPHPQ05x0/2Ws6Da7J9BHkrCo0P
pfvV8h8t4nOvZsViJ6QKMhvPJUeHE8d2RQL2QfaF870r110a4PEM3XTA7YE1ytMkiJdCS9SHlUCT
3jQ+quilA1PkQ9NKcfrXJgsSV4Y+kzwRnIEWCJ/B3p3AofhVsrrRGwD2bN85LdiFX/W5CA4xuEZ5
OthyQHhHfXlfw6uGQEpuBdmQ4J5K/FBat2eobSALJABBA4oA8UB6OCTLHgX2wx1YdZnY2O1Oeb8p
upcc5V+RUarpWz7oXd+Hw8sKGOkrGYxZlu1ACez7IzhWX7bU6z/QusY+Su8aJDhaKgVo97IR+R3A
ESAMb76E7kS/kH/cm7BWD3G0T9uZHbHFdUayaBI33Pi6ZUg5l8cTWsc+rzwahYd8dsBuJ2fc9Mss
+rQonjGw6kRc77p+ldvmmgvXxy1ZNW3qU2/L2ZMOqh5BbqJYRAYdbyZojW8FyPKXPqvxshIFsAiU
VS5cYkBpAahmXaQBCxS3mxJdJKF69PWsQKJHpY2avv0zsOUTBFlD4+Oag7nbuzOtPLcp2rmP6tQU
yKp54LqGfyQfVerQnk7/9MeXzJFVkf3EymoAoA2/5tnHUuECNlGKvzzHdOBQmrmD/CWysuJPY9RQ
O9X55nYPIH7Tujwrzh1V+6MDl2axuVnHM6juUjbcp25BOoJims5LwI/gnRWc+JtozpSAOCEKljLJ
uh3y7JC4CiX6TmlrWFDPapd4ZJXDMtaiJaMiN7u+KFStTfwg+f1XhdNi9ygglWE60BZpLFilasH8
G6O9eihmRtdiWTJf+WQeUON4oySfrDwQiFXAIo5b+QgOo7QDKepWNvqVNLS5ewpFUeZ3Uus/IITW
HmT8SXfo+KiouWEDbpeiWGuOIxECrbdx9AM+C3FNx0wBy4fjBFclwJxjzrw+JzOGwPWXo6IGBlvM
vHs69wx8yXm4TVD5Vp6wDViZ+GuhFcst/dX5IplAdhaOlDTuwxvUw0FZ4vAaXb5iu6DXDqHwD0Cp
TujnE7jFc+C1Y8soyPaZ3jvtoz9ZL9RuRZqbiWq5TZpUIi1w1txgVIBvqO+581ezfzqEvsy54O+W
dfJsn+QDBeshznty2g7IPjqTLwUKGnqINQ1FxR/fHGbX/xXyAsyp5jpe8TzfCmpLc/eSoh9Q0p99
oBVhOFniAIIcBJTciiZJS/lhwtm0LusYoiqJF4LIm7mp+c1EOqYR2kCuKslFuynKPDvFs2WzeBJE
W8bIFIj8fPB6Hf6Rp/fJ1g0nuJEYMZCELn33aaS2jZ0L4iA5sLwHTUaJIjjG1Co86V/N5Lu9+mLf
ATKbF9rjZvnGMg8/Jbyz3rMHhSm36vBZ/u5DnOiJpWxT4t03IFzzCbkBNMmOd7+RpkF1uNv9vr0h
UNziAiaJjnREpJd0QL9H0Hgt6EYMV/OULHZWqpUzp6mKYZaQdkaQVZV89jO7EEV+AXbETEXKJGwa
rXEviXX1utY6b9IMS50eZlsMhL1mcj7s+DUv2ynuaWCDutkbWKRX2b3E/LB6z3N8oNoXP0Q7AgYo
P7gAMbgu2ZXo2NZiere/V9k0Xvwbuk1M+I0rPyONprCENJ4cjeFzlCg51K5ugaOPhd3nTZw7x3El
tbuWqBpLvLCtltnbiblHMrghtOCM2cpK+lnkWHGl1+QY7PWHDVptFNxibYsQbjC3FQ3hGCyzXSH0
MWTxQ8vaHf5JhhPhEq5xKVK9BeT9XMhzFvEXYFPysSaZapF1Pevi5IDl+T5FjtlxCfOrB5flgypM
aD8YyWRDjUGYqBXACT7ktOpOae895MxZcZTHzDkK2v43xj0i+qWr+5BeoXuUzRrN87i0uNWOws/2
f7Ze4qlS+tiX4kbmOBm5pCTaXVg0/YPlhv4A6wqHmZvfxlRXOkzKircKDGhpHvSUhQ9YQWcw0h/i
M2iOaAK6intxld0twYjQyuayXx9Rkhkdje56SlVZwe6gSjxkM+kjLitOPV2wgZC0Hze0aw1chyYP
Pq07fQ7SEvmeAS2LCinLxJOYjl8DVl/nJ7lfi0xJ1R8Z8sd1rgIaplLQchyaY1grFQJppsm/Qcrz
Z2qXEXRxRsE1hhO4BOoBxWemm4VKf9pnZ6QdsnNu3AwG3gnqd17dc6Bj4DVjfxTUNZFsCSC7LTEo
4WB2ff47ocWVfOGqKhc3e4c1e0VyTkVtp46pZmimdHlhq2d80bYoxifwOgHfZrkDBfdR4EfeKOtw
iPq6kpevTSWDspeJlhY0eddkr7AtvNn+IjV4lPlYgHFSvGH4W0wpXicNC6vZTZHUjJ+R9foKgegB
+o5qgL/NGkwB7ySOFk6eSt0O+Hu7cLzvcl1DKYJt1DPraYZ+X23Ui/VF7DcIEOdiw3wGWBiSeFeC
Ng8L5H8A7whOtVap8+Zx+b1M5yuv32g5DUUcdCVFBhe2f3IsVGNh9uKjROuCsf8vS1GCcWepQSSq
Npnd62U8XSoJjbx7l3PKyZKMoFqctL9jKYqG1fXIalPE4CXJT7LKWYPhnfVVdz2yQ/H+AhksIKP0
4/Y6FFqGdKhs8FeABMSRtJ8F281fhvGzOa5qOy5ad0x1QJOojWJiEuQ8xvOhWJ7IMBGkyH5GRejo
xa9OYgeAUOg4IhveRg4nwmeT4hXoCPY9MbZQgt6XCtRxWKT0vPTvJJsYglPzD5GL29qTqamKZoET
mdnEksj6LTc87CN+ExK5uxdmnokAoosGr6GzpMYTyirfW3xeR4uyGLQyj5p/5vpWrx2ouJTk1APe
4+m/K59r8N0Ijk2P1jOgIE4buVb0TvqHtxuRCypQpsdLy0x8BWwepI9Esxw3asSgy8Fn65fOWUgT
p7420+G0UyRNHKktieLjRxNwYMeuoZ881fgUfJmVRmHUtIF1c5ZHFvwYW2cKu4q10yuS43jqsw6E
nhnr0XMVVP9rPBOEa7eNVnCgIMCAHjVzvNWJmAUKPBmpCMDSKUwKm9lxTgshfuJO7Wu81OjM1tzj
z+ZJxKqVEYYb9Y8s9VScnYsxv9AcKkhIhtusEwI3Rzr/5kyrDSLS6vEQzORZWZCLvi1zyDPOLkNi
mk4mACAfe9B6S06/qptL8mnKFP82jAwyXPtPvL9SpSXvLWBh49cxtdo7G6aMLmRQ3GmSmGUFc8HO
aMsXXc8l6iuM4v+Kf3qwgjkBxUICWIFE7bmiKc9n7xzZFCsYvybXP3kCFkAg24zpD2b26+E5ujtp
tb6BGgCMtMHxKZxLzzgTf8WrxYU69iqRjiNzTzkBvVgCAlzlACaq16up+5nfehZ8q0dbQbIZJ6S1
qSyCwtKFus4BxYlh6Na5ZcS+wTah5/av7RN+iy1HNOOkkp5fwxOhz+y9sdre10JwhmHytkZe0Z5j
l89lcUKC/K7XOVyEsDRGSFbuJ4fuMQ7KiVpTrcADrVgkcmLq/jBXh4zA9p4f42ijoh2mKTOw358a
Q2zGfdrVeQzxxlByKoUHdsQC41PCEl1DXJ5MBVUlC6anTmm+/j8WETUEM3SYqKTEOyahWh+MIt6m
E0HBEo1jd+Wpw5F9RBeI/6vRRK6nycEamvqonELdfEYMpEc54mCV3g+CiRHCnjmEjG3OuBju6Gia
aZna+YUs2Tc1qCrL4Wj7TPZeqVXGqv1rzhySji/L9BzOBCM06bonptYUevS8F4Zdzg5mqlifMeWt
U9Xb+mjZeeKbF9JTNa6Q+SONA7WnyHWMimxCjcYFtv0LtYMdLSj/b+UCGgcAf86Cz77Lxlyx1B8Y
pCjbEB6aCFL/mELJ/01b8DRBpNDDd/ApIGtPZNWH24zQ/8ji4UcQv3D2OIe4eZ3kg/SF8WQ9A0Hy
6XcKaPd8Nuzbf62JXsozeTF+Ij0V/ONGG4j2CE2ip3K0kIq45Maug+JuGyoOSgrgBogw3pYowSjP
6ILgY0EplC7w/SiR+rVCpw6IKMwsIZ7Us6lUB0XqX/CjyAqJqDPuC1bF9pkprdGv1AtUmXF20u3C
zfT/wvSX4eEv6KfIN3WYJqywl+mWJmteJfOIsB3MjyarPYt0n31SW6bTWNsLMYo5waSXKMc8qyU/
LJXr+EGyQ9WeaJVtiYLmMlQI0JFoKhJlqe6Lxhv1E7pQrD7MT+mtaaAGf46Uu+YfWPFbkMHnV8+3
5gOCYqUiT7MCIw2MzX2HFWmAkZqynOcXDtRvY9ySmQphUfrQPdNysCFfb9EEHVq2eX3aEgwqASyp
gW8zn5BOfi6uMMuv06TkBJgFN4REuARAuc9f9urV5rVXs7R4Kyd9AshnANsiZSiafSb9gjUPhsoz
eqZkbKhCZt1HKaPqGeeXWbAdEzmL499tYPtUCb1yVuzolfrQOYESfWxOuuSbhwEZ1GtIMSb8e+jv
BkbA4rFkMWvTyCr/iLC92vh/RlPJSIshm4aTK6isjfIrYFPjR9JhYjWyVtQDg4wHYRkz62hxuOn4
bxew21f1/SGuOPK1OOyvOUQPXhO7PzDiwQ3IKCM1+W56cNe/F4x7T8TYXWwvibVgt+R8Pd1Mn53Z
jPjRnJsHikdWv9yZ1MeOKG/GCySE81bA8y7jGHM9rYkDDJInzC4pkUgF76/zcURc+aPiEWrfZpN7
0oVBcyuSMJ5RMHMnasJiegquOKTyEnjlaInNKen1INbijVAl/SD4+VZXE6PlnMSZfXdksv6G8Ggu
8kpmZcPHtVqaZ5v44Wv5f/DXOZimqLwqDbb3FIVgap2UB9A5FpIsMixqRuOCIywaOPOl3HLZ6n9v
z/YsUsPzurfs4eePEp7wWjdEfJgzAiv9MUcrQhLzLmnvscSgGV9qhtWtjdyz2aGssPZACySijtsK
dN+d+IiH3X7A0YLlBb8cxmsHfCUHdOyGgmi8eefSd+KMALsp3qgc+lsPGOjynnFh1FxLljPJQQ83
q/rC6/ff+2ZM/0ADYOJ3xkx79gb52w+deDyXLzW5mkKvUhEgXVzLj/kTEF0Dt7c1N8kBiKGfGY26
9VezEIVuJI+bIpMCKRpFhc6A2Bw0bSKGfawWv0fBN669gNeLefEZXmp5r9AvKqvuTQ8WOS9bHAQi
QPasgB/p6yHwAKP/WQZATCfkfoHj+Y7ivgECtY9NFFbx7h2bger5xHJoRbdBnmZ2YCQV+NVKUII2
qPXpLgpWF5r4heQK4HPi35cjN0Pn6SptUspBKYFlrFzkuK6DU33jqTb5N5m4hM/twcMk/GkcrjSA
gwpbS8WgcUSi9oU04E8W+M19EsdanoxGlzexIQtrxwlIPyZEw8atzKzm6QyF9UjOZ7yVT8sjC6iU
ijWnQLbtkuByMrA2AFuZQwokJp2VkpyXRrQOAuDM2z72mPEQUSjDM9AznfetYEtt1yvJ7vhoGpBA
248PVgnLWbYQQfHmjWs6S+ZeOFP03aczcQJKwxhiUY64JnSDxA4KJsqmYFTJoI9FsPie3RzxvG+u
V4ER5J+5DCWnCzDBN7jyDF5QmmaORelJvPXAfGTpVg0NBLNl0a5DlLiPQAIUn4kvfNEirlcSZpV5
GY9Z3R5/qIThkhIGlX1+afqIw7QVrljgB6Q+ADO7AZ++gwZWCZAsR1eI6wUXvqMUcRLvKAkzaW/P
c81n0S3XJneAOESGFZv5nXDtcFc4HG6yV4BmhXWjBhG3VRvyfMmJiKsLafAMeUAIPNK3edeInfXb
hvH+IsAWHl9g7RKAHKZSHzv6Dxul++0v1Gjze3igpdbR9bBPj9MhtByPyqnW6uzvWDdduzX6xsl/
ImuOzekG9d2a5wvzMdBJu5Y54F+/Et4sqF0VGrQ+kHaaCJlhweIs+rDW9p5aVwclawUB4ohGeJ+s
/ARgGE47mhYItJjR5eOEaCSeZLaAvdAmUW+RD4iIyjBgFgs0a9kIUmhTTKskestflOf2bAhYiPVr
8l7tABsaU35wOXB4cTkmpn3AO2nVpEN97Kfrr13qp/CNMtB8dHs7IXizCgjJbFcqCeUx/duXTCuF
M0rJ/2TswKeQedRc8fAnZATrRB37+07w+6pao17iFF7Gim9HlovDf9zesLSYs8nARlIz2dErm4uR
ohVfmXfo7ZnVmwmhs4obsgYt4EzuMnjjsAO/M6EzyQd+zOybHp4NIqLO7QE/cPabbHjsWVDWSv4c
a8DLSk6Kp3hFK1Twx3e/PfHwLM6KRF49jfzU7yOcyAyvkXLjswp3nSxPB1nQcAiOIi8+MK0vt7Oy
+EBKsNP/ud9Ucn7/JnlD5PZVIXH/hZgdlS3G14gNsmeHa+LlGf1W1qez3kGOCWKcX55vO9VTEVz3
4267bT7+GAc3e/yOIk8MvfWERYbvqTL+axbHacnm0WHpB7vn0Hyi0sa3pZfLyLu/YHTVV7QDH4yL
On4aKPoqmSEnam/+n0ahGDb56IuOuhPatZPeRjAkUDwFGnGassIEA0+TE1cRbWGj0KuUdk3jWDr/
NDuog35TaKAPEcV3LYrHy4IoyUmQ8zFkKuofgXmuGAZlJDx8kNkS5FyUxD6KaitcBNRLYBiuU1Hj
obHEXbwLNYmtHf2BCnQerrXuL1Sf1MHZI/2R9FqqF0O8eio6gVvXVDOZZXQ1im+Wisx/JZFK525C
KnNL1tdYnwCky3rHnMTYa5n0hRnNzSSWKp32fcW4iNpfNHEYIC1dQACHOz41cR1+gNwMWs/FNLMu
ZIJHkXJ6rMtaopN71m7oQGXDaJA5w4yOAjdtwFg/Hmrao4eUJVGSUnxzX+rKFwTBM+35M2oZp8ny
MIDceopTvyVMqsauasmP2H4Lq/Ng5XJcJckJbbDZ5uDumQetd6DuAq49dvtH9RIj9Jdi4wgWxxkA
mZY9gIufnVg2AIOLEP60pz45773lmce8Y/Q6ka0QYeChfwHqWqhwNLHGoZLRSXCUgeqYMYAsRN+/
4n7XN/tdPLUrq3twqgbgUuctQ98Ua+pVP/uA9ITr7rWk9RPUpH8VA6kqSCo2UanlDDgwWwjntkrR
sK7zyqQw3y6FMrltwidUrZ25MoK3iYRRCh06MkOq4qvcTLXBizYSj/Cq7oPPxuaKpwoG0v2mhYyx
qczx1I9xZlC9mMPwWaZ2eJq8UfMuoGVksqNg8R1db2VnAjsQaPdS+o6Kf6JDvJNbKSFqGV4y7jlm
maDOvZ7ITpytMPTDO6i/pZkaaaRViQc8O+Cvb9w+aUEmMUI7dr+FqDf3mcMKMXmL3U6BCdzmU2cg
k3ibScZtEgmtHrVj6/gKPoR2YYJXWGUAVamYHKjZS5FTiyg0V1GHFnEjJXnyUUAKQj95+iq+sWZS
pWefUDXS8d88DxZfdCOSeQV3QYC6UpxUIdOcEv2K5Db+aLrFP66fek6Bhaf4WC250g9i0njk7HCO
fAZ7qv7rDHInyR+1b89ZSo2dCnAKup1U9Hek55B7T9If3Pxwuj9FrJsmWcvtgEd6idZjJenakmt/
IybCYgFFOqWTp7IMiEk218ydlK7+6w4oyls+6pJijeWu9dnu17xQOTg/X4BRRFWKk3ySNcOBzYj3
hfKm8pOJu1jrffrbJ8kMGGnqgNZZKVKt/VClzwKw3CVuX7MXTB0YaxS0SN9FdJKiXwFlC4hH7jiJ
0nxO1b2q48C38W35QJ4V/cRZ7YWo3oqVIJ2lsng4CvN44mlgVlSwT9lB1yKAIgfnZHjDPCiCqc65
zvDSTOvGaH4fghmVl/d+ENuJyCUXlj/PcsHuqTh8JYb7R9CTpgzdLevBSJARXLQZyz9d9F4J87mX
v3Iku23U7rz+8uSC2+BxUQxvWsKa/8Fp9dO9GolT6f6ap+CrX7b/Lw5m+jpIuvhCP0s4YO83BacL
/YhGbZ60H7C+x2TPEuUs3p5Fq3QIECIvZ34jdt7z//NgTB+80L/Ssh+ZTfZVTaowf6TGmxtvUxcn
jZAeFSLkxDxxC/MTOzbTibiq/JfzFX9XHqhsmf9qMo+/CH+wO3bms+5B8Yl5LrErv5yDbjPAIvP9
pRF9SoT+wZixEem/nhlTwnYCJb+4SYgqunWB4LH96AWUbit8MRj2MNazCXhLlNdt5/N+Un2Ku+cU
RglWAuUQA/SnDm5L3+HcqFSt5RX0ZQrGUaIM4Q4cq8KFL3bZ2V1m4ut/Oour2N/XiY4dMw2IbeW0
V6FDqA8Vw4YfEjxuqaXYdmVQ8lpxRpqykDkBEYDeMLzgAGvuk+UjfxDeDWNt3MdFrqE4qwo2Du82
O45L2fj+KRhtioOkLp8CHmFTh31mF0OpY8v/b+ggU8SUk9NNJEyW4iataBKLd8wFlE+FNkVPjEAm
C9PPEnXRHfMtZ7jx26Xmt85b5AwTuCD72i0pKvP3vt5sZ230U6YNKUgMhm+taPJK48fgPcUDnA3K
WmrHLw3sMHOke2UYzYg5V77RQNXYMrxgPZaLWynV478GuTUpUK47Go89rDPdoNUllBCAfHJf4vZd
WUUy0O5JlFCygrwZw/gx9TWdYpJulK1TD7PdMPDfdVzp/Ymxb08q5jGJGiOI7SNS4UUiDAByI7hD
Bc3wfMZ2JLLf50SWwdbaZruax3IkH9KlRjfCwvieDrd/IIRr4xLKfpfIyw2547Y7roriJgR6hbDs
5a9NN0wZxJ8bTfpwL+Yyly9A+fPolduyFXXdG3J6ttf2cOacTZf7x/utIrzbJaNHC+Sqm1uWY12W
3PjhjHq7Juz4NMW127KG55kk/qqmme6Oxnkqrz3LHGfCPkqG9ACsMZ4+595ke06DHxjQjqfg0rsp
2M0FLEMVUM6+vbBTo6twAmc5ltiKK/iUTHtI4+EBHL0VVMMSY8xd/4gQjjyNUF3PYSkVTAJUv+vF
1KBPOiYhtsqibQ8/THDGQIqop7u9haKQisI29AjOWhzAYX0mcxywmB6fY8MjOvp9O2OW0jfiE1ke
Y8QLESqIgn269lAxiSTOb/3BAe0qpyeNzuvCAc1ubEvOXlm5N/PXqEEk9LOqBObq4LPqIfoa5EoC
NACw6WhdUmtiaA4qDXYULaf7CF9yiGju/y8oOFsNGjO/6Poy/7WYjSwhdrTZ0mfDTC4gXz35h9SZ
JdQd1V3uS3fGDcugSrf9e09txLv3gA6P8+RwA+LmOiJcNRcHqVbQslpJNhsaJCc+vfTSSU0/5bRE
neZmcUnSf4yiEmmn/y+mohg8jxvuxT1eC0TLgGkctRqWR14zd3+Dpf31uXT9LRfSRmgrg2jVAs9E
aSLTo7Brayti+Z2YBDIANQyNXLWumnNBd19RhBaaGGa5Qq5vAvVrHQbxO0s58rDk0BQoQj4eo46W
+wkT5D3/37MgaLHMlJsRytaviVPieHIaNTGiQp3+x8okNON4vWu80UVy0OoNfFigoTjfIf665tm1
kumSftI+EoJBc61TNiHrnT8KD6A35ZdBo5VYVuDKVzZ5ezLGYorvcqjGNOGzz74uKi3Bc6am0C/4
D7TdQEEiRMPyMwMo4A4P8jrBJnpCwDn3G41glsYeNSpK/ExOj97Aw/IOjMmqmvky2kp3/0QyFZJg
6Fl03EeSnBzjGiU2cj4UBMrtZyGSv++mZKLiUKyjjyoxgGy4ZTTLq0gPp0qspeIO/cqSIONDnEPM
rt902eyB+j1I3YUCeL8levWppdL7QaPq912B3YBsjrPQpeN6DS+v/uM8q9P4D6LFVBgDZ7N+GSSQ
mcEvGAwy/DCt2E07h3KrClk/PoUeUqpbRTVsPvcshqz86vnny6Ny7cstsvjXPgJJFHhSrrWomDPe
Of36KhbDagsxiVv8ZITbTPmyCdH5BQ2xcqKCyv3wtQy2cGxaez4Dhrww4x3KKqs7F1Iv+VT4thAH
R+xUlgL0PWzF+kfGgVeKNjWe0NyFVeo6aWENeoraGoCPuvHM93WKbYdDdiy+6iwhMMd/+okPhfJM
mVdJLJhd4wFGd/Ve3htlT8zHoh/oyS40uKnBciweWjR0KRGJJEfXzFRg+qjmkOwX4Hb0PPf+228t
0FMGJ86hNPgtAYE8Wd3O7pDxJAUPriH2qWmHxYKlus2WRUFzFhhcBk2cKg6LX9PfuS6BdjSoHbUo
nct485cBVlY8Jcd7VH33enQfX1Bp7rcr8lZ/fBN9t5A3Wk8i3wyQYfSqMIKMZUeAkhhY1G0F16y8
TrxVVv+uY6mERSB1DG5vbGp9Za/W12ZYWhklWMD/ncSjFiT8+8BOTTFpDj2HWVCgIAmAP6O6CRDF
fSQ40JXeUBtnGelomO45yfcxUqr3J2i4p3rdUXWXqeZzyTb3P8udT38DF/Rd1Vd90ebk8HNd527Q
MiSHWmfan9Fbg4qfuUMzL+oAcbbdFR78Gw4dx84fR/1oVcj9ythtEQw+VcVAqBAZBaOTigVGywi3
t3eUn2XtOnRtA6PKZlwJBLeVNi4ILCE6ButHzbB7igPFbHSp6I35w0n70z1ye075ooNYQm0NV3Q9
OexLkrcVM7bXQCr0EcToewe5+IVgwBsG38TJgC8RcohdYZU5Fge7tbmBnHQIrSV+HupNWXOJgl85
+mcOO0Ce67FwZb70/6i+ly5LcZbcjj0Jz8PDB2cgKsBlmvUNeqavav6K9r7ha5s6jM9iWHlSjIk8
X7wMSd42LMavZfT+pEGehyx3tBGan3s0FxbsEHjV361WjH/ZQq2bjALYvIapySROB7MO1ybedtkM
wbIHeJFPnaknlAsoSF0my0rhizRos9m62cfvByFdF2YWKpCEEhkdekVmx6pdLEnmYbIWC5GPEtIN
9o0D6yiU17mvne+ah7LaNxKs/xjlyRJom8tZ7btcBPCzrOl1Wcd9QIkVZt2q3APHwZsLzFVRs5mf
EFAr7GRESTuSf4YW2qCgGuSQj9UrAk0hK4eagEaRuwaZ0dVz7y4nua9BockF/Y4aQV4KAH/iQMBb
jphgOPho8Ij5j4w5vVq4eb4ybsbEqeXBJUX4MAF+csh3akpuQVoYmv2HbGMLLa6IkS4E4zaFzAIx
e9hARfEumB0QMI6xhhvokF3HIhgwjRve2Czvmp88rsD9dYwCkxjAV60oIr9FrfUi5yVsTi1jprS7
Lo6uv9uNsk5l1w+EMWq2mdKBr0cjpORFJ9vBn0kaAu0BnDnmOoU+HdjsK9NWb+rBxunrgaQ7vE+v
IFN5Uhg7inbFG5ieuJl3+4VYEtEFAGQDqVepq8/Kyv10RNmzdUOGbEXp7398j2yWuhMdW3iZzu71
vaZbzlbT//qErZwsZFSuZckLQmh8342rP+7U4trpJmnO7AjyNbkAUBwLTl59OvEV9Err/7msaeoN
hFbe9HJy+XmZ8EubzGXti2K2kgOuY5Q9f8B4kv8usmZ1I/DWiFnQaGSRPMmAS0MYL6xlQ5APoyc9
UKaE9bF7tnddNBWTq3Mkvi+mJunPunoyEs79ikLweVfalKVdv7YeEXbXBmozSqiLA5VaJfVX2Vj6
WCloxD46krUoJYsQ4SjFajcCfDnaA9bOlcrwC89qSqkfJSm2fa8kjB3ng5kEExApMorNxOwngO5W
74bHYD08By8VZj1hjRO/XBlYD6MgOIXH9Wx/enJ4BPM6mVKQq6HyXf1M54oqacC03C/YFTiWIIul
yc2BYwMXFJiU4RCIQOuvR3RIQjJXEZBgXP05DtdX51QVuzzxOGCFN3I+iTG+y3q4Qp/5a3NO8N8A
pIAhjUuSNGgYAc6YKTj/G9e+B8MRJk8KUKTyrxQeGEa7FQ+dc3zzTFwZk4zo9yoB+MVDQr7ZomlB
IFO9Qi32ny8AkfmwthY0FzK4V5hIuQDoVd4xX1Kw9iG1lHyJr1CnF2vGpEMIVq807vcNcRyMwAOI
Bx8X0SIN+L4xbf0HpzLTEm7Xv2U87nF0dehq41uQ3EwVzyOpd0LE6IwtT4uW/zGsdTiFjV2mhUbR
SeJLV3cOamHlazEB7QHor094DbU7IXfJPdBn+KjtmGJX8do2yJoddieh84NDAIqUXOOi0PZLX3U8
FSjng/iTVFSYm/e6X/gv5FwkMj0IMjq5jBMTQodtvh6Ay4kiZ1IMPKMzFmYULhsX7+i3YwEMbiZw
uqpPrg4NOyyBzJg/BvHolpc2og+jTUiCIDebbw16785lRCPh3c6UqlRT7nxMw+HY6v36Vf0xdPjf
ClyvxcHRPWMfisGuiEVKXH83oq6FdpPH6sQMbPVeDnoc+qoR0bLPyNtppGhfA91NnptKsEFSDXYj
+EaayL4bD61Xc2ybQzc94oPESU7+jI5r6MYl2gKW7J+RPAxj5z/0gTjSwZbQfZk/9PS3gdNfBHFY
3sjseLzpnRkONDxy5UYrnSvGc8rFtRkToRO7bbZ/ngWs33KgAjwq6dyJN/ilC/wFGm/JAKQ6K05n
qXND/SriU9IXzzeSYOn3oOWfyF464NV/IAwhxOflupWOJE+KhxKj7L/8qYstV4H8fNHiOtZ9Uu7E
naBReaxV8qfa9TfEhPCotFAeo3Qx+qpzc3LLeMpjVT+30S00g+SmnPMYRDTncWWgiAFxq72wc7Y6
etl7ueiWAhBmrTqo+rrlvjIwBXLZOjgVVuDzvMd1mf2xQa9aOZiKcw0VGMHdeSa8rFJKjtGxmqyq
bEEvHLJShGBm5rqsPcBePKkGMIi+q9pYJTB8n5e91Br0m5HB7rnSnFNl4yXq0zx3/JFUZw26WXHy
FHNd5oFiSzLGUQuMVjOSSS7/kb5VesNHblSUyYg0YdspyNHwQH56wrhvAq3j/MgBrm06y7ZUmubd
Dmc70P1RbV4nH5ZqJuihMeu6AlEEfquXxhddMH77pa1R7UQ/3tM09DM9w/0wLWvRFRhBL9x3kXL+
IcqHJl5hjsJniZL7Dc5ZqB+HSZslg+HuVOGmH9O23lZVKAIU1siiqaaF5ejvof2343oUuEW52Mxx
df5GehiKXyT9QRjvUus0KdR4Ioyd4xFaePffu6kWuY20bWF61XcHWzuwGhuHkc77OfK9v89gx7KW
UskgtWyU42maAlEAI/uQjrDt0mcvFTChWt/ggrd0UE30zPNkVBAuFXUEeqYjmue59hjxyCzfYU1C
HUk53ImJvryNm4FQNnX3/Uj+J51A7+HqnAv9l57+woa87M25LmkzXfJSD1SS5eHLYoTohaeMIG0c
eFRgA7PpPRr/VcLmaUhxyE+AmQn3I6qGq29iEfoDodPNG+hgABphojtDIc0LxoYoSNJiI08DvG90
nRC/3D6BcG19k83uUr9TRLevhIYPSnImMpiq2eIuMYtoxpmvrcdPBXSL6wcJ45cdRIwZk4VfpGj4
4LByuTlNLDaXTf6eJOM4/2eP7NjjCLmO1T5SxuYzGDJR2eAAp9E1fSeV0SLFJN9ZeG2avEDNDllP
hbot7TmzKDUfv3twchwRtYRVbn3OKX93Wy0alN/oX9vwUloamRJNkykKThc5mcriBRT9hD5O0T6N
zko1Ys8WwV9Ynelx0C8hcEngjnvSY8fFHTmHmafn97oWsAbJ20YCNVkjMLOdIIPTvLO/DeSQFSBN
0Q2hpeVb5hCkzwjOf8dSOAIuFw5nCsEoU/P5nTN3VKTkPxyYB2rFtrpJEk4Hn84x1H+TRkrCwA3D
DIOmS/CmEvcdwwcq5kvJJLkRNpwKSVeu0bBcl8XjIq5UnFYD+jTVKnwuOGISwId8w52dxDAOnW9l
SHHx8hwdXbBeVG7EkvQ5Z9AIvY9us9QjkI6DkTsUTALCzu0L46PalZsVE+0Nmb6ygpXURgDHGr4n
Dmd0mWdBggBm9P8nzsD2nsPdALGpn6AFTd77UGD4xNDVN2pTMgOB1fiXsWtJDca7bD6pYtbc+23G
wLF3sR176jBwY2jzoUOU94PgawtA6q/+v5J3xcHnoOFil+JsgO44uSMue2OBn4i06XLTBO0rEwG4
MgDSrMf5YKmEsusDyIqcEzTbVrnraNfzEJkyc0uVch58acHEiHQitNEH9i0YKaa2cACLHHENX15u
45I0O6mAqSrRX9wIjD6DYoVsOO5D0J1HJpM/mwGjCcxk4gPpd38jJAvo4JiqUHnJ9xXiIFVOjbWj
N/ainPKRkt2LzuqszYV572Lf7KQiqo9jcgekq4066YcJZaseEYF6xrijiBR8mk/cb0GbSG6/7lYS
lc2fTowdkd+3WwChGt8MlhAaq5+t9e3p+u90UdB+372k6BBZD3h+69DQRXQ0dE27crzjy3MG9PkQ
6WJHVEVQp/I5EIAHSf7Jl8MGplTI5r3ufWAKyHbUefg3OOzQjRFtslWWi7ev1ol0QhTXWNfRUvIE
/q/UvJoGiffXRNsMeIhoD1+ic3HCFq1u9Ze0LO2Fgum5Wr3UK46QiHcOgexjvT+VobmIUgpBfoGY
x42Oi0uxgYTISKjsxt0wgGzUwQsreE6eSGboQ37aOweU1U7UTlAliqSaUMPyMV8WGz8x5WgmW5GU
rmWUAUGjeAbp3/Y+3VSCu3J/kblt//uPBV1a1RjGYJ0a8+XtiREkpGl2yyI/YcnuTpF9xwiBecF9
sfRHhbOilqt8oJdpm4yNTzAMhyKQvGPNq8Sju8kFaVUYNNaODJA92UUzWLJBvCOrS7/rVhR1w54p
ADVUgxJGybBLy3TX9SQl27YJmK2pNRBDJuEZ1KprrGKUiDL0LPPdf3vsH6kAKb+IfzAtR1KzwVEr
QkU4FmmU1n3GURHd/3ar47czEMxJ36EYAzzN0giHKOLgXFpTPbm1tMtULRNBYD8Qo84EhwOcmjsg
CllyrRWdjn+FIRZlwH3+7v6ffmMRasYW0SjRz8nHqP8Zgga0Ipvd5jl7LDSHQ4yWYwqlZWPVjk4K
EJrOLX4pnwtrAfgdxqIzY5mVRpErl9kFOCCdPaqj81er/xBtH+BB9Wxo0tYNG02QGveJtSDuigpN
XzpDQPvlPLIIOOu8vzSWnqkzp6exBgmmgfusIReo4WrQW9wpNj1GYxmZ3leD+gtqEYbpCE/3ynSF
3GGVcbKEYfzqAVzqu/rxKq1UDvsEsk50RTLttceSvM7KBcPuOB2zwvQWYcwM4INkQQkENNaTjULY
FxWwh2XDWTAFI8Zd11tH+NUzY38eD6AgfWuMvZM01Cu6BU4vLEiNreW/y93He1TtOdpAm+E0tOpq
6VqbiAar07/5aPwH2QI8yJnvR9QSGRjOP9CrFD2JFNSTA0wYTAuLkx8ESWrSiSAMp4/JsTujw8E/
vo3Grc7LOlQQCCsqMd+hpcy9wuS6+KK3VwEjEziuLp09ldywiiw6tWXg92+YgggqKNZNNIarZptY
7A3eP2cdIGFN2XVTRZ82JWKSqSc2D4+dbA7SMgP71VfJYv/+Vi99a88bpYpjOkFX8omk3+68xYgb
fEDNspz8vYobg0goA9Ed4pDPxhky9JKOunwhgjL7Txm++n/1WEpKzsA/tO9/HimZpFgQdYdPX6aW
bbErF9XinH9YIYbEWUB6msPiCZPYoJOyFR+t6AyhfuWs7VZRK0mr59rFNR1mDIyZVVlzeuV/1pQk
AD6N0rGFat/zm0H3MW2GBH3qZIbiZ1UntPBH8rJTMY39Mh9OZAxFVcfIBGOTk8NnUrMI/6E0Ir97
FWe85DVNWuNTphBff82K45+qbuza6on4BQPpuGMsPp+8R1MTptkRzrLjihbSPhLv2neZygvNKyqv
3GMQ6mSs3kqvSR67GAWDwU5pbzACNQs3tUshy1MPiKaw7kSTo9qL6WzEg0j58WM9Hwcr+GE9zwcs
LAR9WJQCz2GGuiLGKT2BtbLcqMjnq3PnfGJaWYVsWb6iXxKwz2yv0jnJmhR+EhmCveI7zKVj+TcG
tXrBa2v0GKvu/EpMKc89Ae6i74yD/X+TVWykDxJXCd28dWcr7cdi3esMkK3t8KAVRF4kqb9Yb3SL
TdlevFbKfYYUWtsLJgYN6ofYpchCJO8LLlYLmoG0XQxR+yNJn4j2kqfHmGrhy7SPDNvxOa9m4u9c
f+pLaTRRHT4F9+IEnnuatVguW/LcSKszyGcLBlENoa6IF+v8hdkL9mrye1ymST83WgWGUdWeSrz5
T0nopj7D2mBzbnLt+2OljUwCAa/1g3VHl1EPKXf+rzL6FMHjuUq5XmJHwoghIRhV9IjkJjY6Zwfd
CZ3JIzZGsHXQ9c71DvkVc7Mjs77M2BBRRScPq0wxFQEznIzN1Y5g9OHUAW9Yj5ieDTiU0sChOrSz
6dScAR4ZTAjgUHdh0EKVsBVXAUm3S0SkYsDh6B0piS0Z8oCZM3/orEg5iqoMfAyVLtGZLaTV/WuK
AmR53nmRf/nj1KQ1UAX3VPj/vAA3O9eMNzOYdQYO1n30Rd0A21kqWBbHTAaT7r8IGuHYtZBrF7pr
5rZAURcHVfgnGryIijGqr2FOPAlxUiO6xmoDz/M2cTNBWOPu8FsfngyYLAhXZ6j121Ad8yM6O+Ju
JozTp7hdcQO9j75qkf7XFLXieGn0e8wDr1WMoPLfvM2fX9QWvrsPJ5Cub60eQejO+qMND6entQrS
S4Sf6+CyagArvWQBLISZ0atnOU72ObHN2dG8l7k/j2bSiR7c1+vlJN0cdRp48ATc0j90/Q93ie3Q
Ch+iCPmT+5Yd6hQmcalUi8LzvjdQo4ENZOkUWTdozdwbqMgXZcsSbr2hmeRLkDVFWtZ2vU7oiagH
oxmoSXK5ohWh0o5+RA0S3nlIat8AjYx6sjMO9YF0RhGYXN+rsbQYt6xFQqz3wU/0o3RxCRSNToF9
Efe1HJqYJ53C3tZBXldig3Kylp921LjONQVQF3atvf0HLYhRmgi5wsy1zQqXPGUpdAKMTG1FA81q
EKDKYblCoiHYXrLAu/XnnaYOZQCfHvQEL087zLYld+Cl1E+Gi1F0oVMl6sAUpr9/e9ChTC8bbQPO
nN513GwWTrD1wHcfcPLcVBDSQLU8BxiFFhv881KOmhgzmHH7HCPugyO/U+Jk9YAKGmi2LVDntPO+
H01BMDZAvXsnaT5UAQuF3v1AmuB+YEKRZwfuD4gSxYUyBHB3h0AuFIhtpIvcyxGdmcJBx+RuAjGN
sv8fF22uK4EauDd38s+OwuyXk+dKIwrK8at8cFdmb962Ar5V9U53qE5dnZMXxJioBLT5hcuMkY+/
lmUufcJfUxuTPuEdDBRfgFpADv41ncq4gkKVpB73FaUJ+4SU7jL5XgyQ2bVg6JzhUIcRlEJc4rH1
62fkLxJmjA5u38H8rzQOMtgOwpkRYgOb0D0EzeJ1RtBEFrExMedc3nFjUcovAEPcJLGdNvaoOJpQ
vN1S74IYiFEEhroGvswVvPWlk8jhw2W4pT8PeqP6tleK8gTgmzx4Glc0n8fX6QUhdg+OjogCj1BR
QS+jRHTnDMKEXIHPUd/lD7v5+RgFXyBjy920Mr1QJqHOkS0DEQNtCw0wTWM722Y/9LOcJKGErLqL
HsaSeqVqJMMVSqBhuLylqFgSml0OLWGTaKRa4yOeACLZxgbZg+/QY1B67agEBoNbJzzLnCwC2KpF
cc6Svl8LC9BZwOm8sQUOeQbM6bP5nGE0osw8cTSiGID5nKAWWI5+7ab6wYrR4kSKzp69MyQKr0vQ
MP1jqoICPJpInpB2aX1z9GaRye+TKI4mI6Ql3mG500RH6K916u0QA6TjwgrOyFOaQmg/HdhHMFTZ
YrzBQHmdLZq6v5FGqJ/4KNImoV8j5CttnXm2+Arq5YNh7lvtXGTcG18pxNM12X/JrplbrCiitJ9u
Ijt9E3eSIhfqrH/7zO/xvruh58M6MFgos2YxgqRrTnYzh4RlFgh6ozRJc102sq0lNzHfWIssLC5K
HwtSD9YSl57tW0RuRlTJU/0KnLAjTyBjora5YJHbE8a+b/UKD7lQFNYC3iPl50GrTKj+ebATlYK2
LtBHO8aVs8PUnz52hetpu+CPM/iiJxSVskS5HSotD7cmb6cAX5u7qNdPu81ATeBBq6WBlahM/f35
tnRAxdGaI/xDnGdxAiozwBkEyR0VDDXsU0qaAlLcFszWsL2NWY5KI4EFp7UWaae0qqPbr9ntafJg
69cEdaBxdF+1l6V3HzUN/NMTE/juzGv5ReEqjQ35TekIGySnbPZjgO4uUAHlOTndfIMc7Gvq3w2g
/0T3owtVW7jT5tTf5X5MFqHuoR0T6yHAMIMednv+Q60F2d9WPsxWDGog8ZZT8mXEZ48gpkQezg8X
WFIU0mbgGoMyWuL1dVPxUzcHaWChfJJYhGhKMmuiIkMw3tkU2OoJSE5D047buxMDvgOzeMcvb6p3
t3teAG0snS9rNqugoyyQHlORYSPUTbIsqf2AGqhBkHRbQO7qc8aMmW5GpazzWa1V3wPBuF2DXnHP
r2T39j6/UDI+/2WYHUwvdlC7LjnMd8sxiCWdO9+FE0RNTwGKrk1WCi5sN3HQ46JknzzhIKNTAB39
WdCMmoi4InXwi1TMjjou8kaCMaAVxucxp+qwq00zel1j0eWA1n9gQJqpFkt31D31q/S5mjR1Hwah
7WbBlJo2Z+TCxDMjZUvQdBitCvJh4aqt7q6dzqazx5JCEClwj0AGqBtTkzQlH3Ecqfaod8JB24Ps
gG9/jbl/DZBxHvbCm4OFJcbVfpt0wnUWnCQBDx3eSwvx+/zzA50oekgVAowbkAD6h2rCq6Evy+gP
xdYXXy7x0fIPm3VkJWCsq3s24AK0kvPPVRB0ZTnJGFmgQm33DJ89QJmTPX4gCUXrNGhn89HYbQUu
IhSPJynyljPx+tmzM2YdEQw7jtTUXvQlzKBIOwDL/dtHmsaDcKT06MtqHWNsn2p9OK1bhNsNRFNb
VB4VPpgMszPdVOanHiNaCocDCJ9cu8sOk2ziAdmal0i+9Ft4m6WXB9FBimSIXylUWQLfUpq8hGE0
m3f/EBZfunL3mpF+xUNPjN40Y/O7qqoPjK+bx9E1bCGyuTFZY1DGpi1H40W4OViyzORGabEbXKlP
e/AE1Ro4cLKeIlyl29wcJvFQtFLzq7vld7SoSpf1sk1xuzmV/NRpZ7Lv5HIskfPy2UhB0CRKKBtZ
0RhWJT2rs6qwUzOjC5W0IoNBG+pS4VjaH1wWdxel7jNIG9MO0PQ79QmOmcHZKRfgJytXtXX+y4Ng
qOrelhlXaEZl0LDfjGYZb++6La3AnznwPR/AaE0T3Px28syVLV6yE4O1a/0eOONxYIGkB/g/ao0R
GepKz+M86BK0TqD+KGXQz9Es3phCL76FdjFvB5wUAV4PTkrFdZkMOrOoLs9hKTbopyJTW9MWeYc6
Kg0i8+U+pEeMPvYI8Ofv5F2pxe4DMbJQCOsHAfgfr+YbhVHmX5NLLPTYIgcvg62Zcf9ENAU/CPh6
wQgCXgC2XDvgKy7gwjB1/T/bXNvgsXr/l+KVEOYbBJvQMcxQDihw7ZmZO7YT3U4JZchCQDQElcCZ
o3dwe+Z/BNOfITvLG9fnRXJWBNAeg5oKFA2OL2yedO87+Npwl+5a54d+dsUPuEGQlWyi0Ng0K9Jw
FatC0QTdWhI/3yW3q+8IP6/Bae0Rjs65nR/JjploeepB9YGJhyR1jjOvcJco2gGqo018ClxSXGh8
SGpeSguTyz5i4Nm/ry62ReBYOrVk0GDRgnND5B8LTWMoVda0Gz0vo1oiWfkhAqIElsS3c+yz8Kqq
MEJFuZ+AvumSobC0U+C5QNXiR+TKbnJLqa7OT6DBKH6ZEZlv6MpWCyZ+g17igIT+n+XQ+PnzPOiK
nEBevXKy7WSEYnpq3CZMwOSGELIIkGdSVK6EXLuki/OBZH4h/lTgtYYVhaNGIlH1a3Mh1GpBtLQ1
VLSfOkh9y981ePbp0i3KWaAA15/jcfA8rzRC0OLxzoBp5TdtBisbQSkSt2OAWU8jsreFad/mLia0
oKS8YbqnpqdjZbxg72WP7q3PI+nX5iKdFZdE/slY/FtoryaP8wExd8yrR8RxPZTJKCCugIMEpadh
Ro2pS11h3vEEJjbcJCtWtgzN2j9csC2kJ27QhuzOnoNrBNA38ArTFApVm4qB6NbwZGKlzyUoLf2a
hrwG0wGbKO/HbgV12dp7R+qHHc4xl2TxV4FycVHswnxqZiJIj1skn0rn5PX0bmr03R7/5b0G9EEG
+wENa1/Md0yectyjVqQtzUoJw8J36qmfsnA0oBEdS0nVCynJsFqeCKqGOT8i0AXpTe21mfBOMF0a
R0kefiFwaUH4Vb++58IScG7o+3lhJVmxUfTd7OtgHZXkMkLveNNExKcbbmdYus3fJ32d8x2mQ5wf
ElX7PBUc3hVgxhGJmNv6yf5FJTDxzGaKT1EHJrMJ3I0Txg6CD/62PNDcYD2wfiPvZO84wHe4vn9D
qozyu799toPvN8+SuDTVJxrOPAxx5horRN0G5CCz1xcSY9+SnX2ZvmBjKuwr2hfMexQwLdFoT2af
LHpR7V8YnBGtCWnQSIwsin0iuvKupiebeAQQ1nnzS1peRFMAemUswn7g+zeY5orIQ4dg0KUXBmBj
8BjBYmZp78b6BsPe1HiEwr/UD6gElgcK3IU3QFx7bTgB7R62hYQoGWdNSIgKLhSfUQP4cdUmqjPS
/qsTfj5jq0/4mj/iKrzYjTRFgy+rsCdPiY/Ac5b0wNjwtzEwLSmxN/0I3aMsH0oQ7N/b1oBz1cNu
ko72YxyxmIjGcwTwHSC2/PtOj2IQWwMc3iaqNdqC4qQjQQrDRmHLJgxsEFCzTzJQdwx2CQ/JvtWm
9UVekQm5D5zm57YR0+mD0SMVvqsVFXCa0WGg2YuCZqNwlc60dLYHwoRfsCsIjwW80qBWf4FVbeov
cr2vbOjcvEkYhnEU5VwRCRpKg9KrInlhuRO64HCgB1GPNP8aH+2o2Zxln3ARL+0knArILdY5OI9C
xLrqXOFyd0HCerQCtgDjX+bG5E9rlEhw5hXvXRKpY/2wrd7U8daiQ0B+bznozibGvVSgoW6aQRWE
ALDpX0dTuAKqmdM7wuwbvWjyoiXiw3xb7wHtdaVtq2mm6G3O8EozUg0koL4rV8ovDOp+YFlUvHnC
dL5bPg/o62oVGicL1hT2yy5ev/9b6uoZmOAfYDCDmndYLJ79HXMhyThfJ90LC3FWhF2heOvXULyK
Ot3sNfpnAttv1br+C3cCcT0ONeDRnCc1iZX8NofI/Gh2CGr1Mk9TNuqHUSJkVtcie7BPAvkvuoyx
AuEKev/vpG8t8IcSvKVrqBIRwOC8gU4JFOy4mpg5Nz5e/92GEADTnZaB2t25cOdJQO1LtIcDj8mA
PsFqeE0H2IqQxzxFVpKbTKUB6hPEncCjSS/3j8DyRNQ1QiP+/7/moL25m6/FYL/euFu4VFq8o4Jo
FWWc8B49I10E8nK2ZcpowZGWIdJQ3aSy+v65tZzXItlFXws1im0T2SPd97NhigDAoktmfflfjB3j
ZL7UhtNXxTlRwD2Ql/Ci8Dd0ELKK0iXu1tlMgRkGPuqDA6hg0SS95pb4r3x6OGs5pdimdLY6B97M
HEwIdzTkus90ffJ9Qy4ssG2lsACXTcLhB0UdgdQx/RSPPomM+kxwLe516NtZyMw0xWBJBdzwmhxz
yLauzliraejVgl0y8qLRbiQcVH/4VjOgrdlkUQm15Gc/286FZu911QLGn4NoQLxb6/m4HEw48kUI
oaiLFyonr0a5uileiGbnKirTVjRx8OE/68wzL6psXkW0Qz7Rx0G3B11XrLj4C+QjwPE4R6/E4kbf
pEJKoD1Buss3g903QRURzFc3xW0R9VWbd+02EbZnUzU3GxqiDGmaC8bU/ZEVkT3h3bO/My0sXzYb
OXkAjRQaL8pUrD13z3J2/4X/bI/726nKQ1y5EJyaq8zfUGfzHPS3s5ymYOPVqFVhcfCqy3+yE5t2
QnCIqYYHCN5GL4EWAsdfFFERid/k80uRwWkTu6sxEJjwa+jaF/QgKzVYtt+z71ub94StnjYnSGBI
3t6FKtIWdlY9pi8fLvO6n8jrhu21r4CqcEwpn0H1ysJaG7Bh8+JXZ/7ULBqd7vgBgaqaNs+5s81D
47IY2ZHcGjoYRwoOdzmzO9lTUGLhynvXHnCvs560EpF7PZ4g95RqzF8HWCPE2uNTWrcqlhRuhCQd
DXENlrDIJ/7pjS9VPWXMtEqzZ0J5ECApJSCDWvccu/GaIHP+o2VBhduX5S4I3+sLvvBrXikGbYRW
arxgU7A/ZbWzkt6Mye1DdrkXjfQHcu2kB0CGWyZRTnZI6fzrKzX/nawwyM6IuUwGkp+yTv4bKFjy
Ba2cidvNLG13urCdhD2PogzHVaRd94yujLpkhD1so3716k+dGA+EQOOg0VdrfPxLkJIvsLPyw8j1
cjp3yBGqAlMLG6gwuefpEtaro44tbdNXblxKQ83Oh4PQwaL3BsXDF4Ag2AJi9sOamGxFOpuMyTNa
pD3+8zC6HftUwNLbW1vV201quKpwXroSPtxWjo7JlNSgybgz28YxhwmI8qeNpsv3uK738fl/VrC5
7U5m1+4b3g0v+KsPoe8+LVkmAdxeAtle+oLMja6l0eQ7c+2cxpJzAoqi0VwPCwPkUUaRFxUaDJIT
Z7llmARXlTyW5A89DDBMfZC3U3f0fK8mmzF73aLdMpo/a9NU4x3PdNKuNNYwqgvKUqdseXSPWP30
/7h4j6TLeZiIRY6/emkldZyCHVUxjCNJF+eCj7S3dMo9ot7NsgBc9STrOfFPTY17FmatI7Pa82bA
zb4Cy/OCklxM3P/J7EOOFi040yWoeg0ojQnDohuGJandE+n0gJUiNLB32XNWu2elpn3ZI/3JfZU+
UCpIGlJ6Wl7GgqZ02r3hcwxmt63aQcOLb5gkceyV58f/d9QOrHARCJksPK/iK9LISCCDaaalZMxl
nG64QzhnDIW/3jEzmVTbVjR5LU4Ibie57cB2XEuK/3tDRf/7AQWK7bbBcbFcWDHOW7Y5PLsNy+so
bttCpPqJxdHP73h9RXdmmLRH16iYNNcGTHkduDbxW7hXoFNzBIn7AyqQo02Bno4SDWYeBhfg8wmt
uqS4AowlDID7d9xg4AGAlsjsGREZhtgoinWFVRV4m4/pj9XZqEFD+nkzqsOKB1HWrZpVlk3RJVAh
go5CwD8Mr/ccjtMoLmP560GIzu4R9xz1slnz8s00AhUrhN+kJPnYnKwYbD5cwOoLy22gr9L73CD3
l62YeKKi2L6d1koQOwKErZAEAhLn/LAqfHDMM3BnkcedRkSuO71ZtF97zGJpuY5OoJGE/HmmrFHk
NQkMtQdlaaNn4HyupyXVEhs2kTL4shvJFBnegF6hC404LoNKKGa/LoqAGYqOx8JgsbZt6fymcwcW
7FSG1gn9fvzSkt4QS3a+FEE5PsAxn/2/t+vXEkGB7lbEBZCI3MAtOH9Ee4bme0D73PWyP+rHtjV1
yHQbRj2MSf192Ja0YqC1Xk8MWfdRxQWM+e7mim9Nfyw/MarWGw4nVmfAlYOoAuQqBttwwbwlRNLB
pwdgsrALSpcDhK2P5Yr3lmA3pf6ee5DClO0ZKd07YtRskN/SNxO4eoqGQsnT+OiLejt1IG9LMvp6
v7ADQlbupBUp9Av+ndlDuOBBqRwNXAqaU4Ep/glGvgg/6BLkRlRmadcxdXhYxLpHIA/hOlTXIM/a
mU8bMQu6hjy8Q184fha2EK/5scRf5sZvEK6pAC3fHXoIuVPYU2OUT+6VYh+AELYbDWa6TK9hsUuw
EzQgacJ2XoCx7Ijd80DFQcC5YBBQDJn3xqQjfB4tDMy9MVdcfnDOGt7Bn0J8ktWiJWylYBahX5wV
fDgYtYjybF4WBxT9em7zugINsQr9239mHMsAvzsq9UjHee9Vg7tUHMukPI4IIGN8AWl0dEjeLBmG
AMGjl6CzT/Hmle6tg6nzYolam2bf/l8rgzwCKNfGrX3MJ5kI9gi02mEtewWyVcP7AzK1sYPcRupB
3hXqRInSunR481zUulkg3KExmAwryTC3PXN/+vc11P8OiXr9hy04YamrG5LHAOp6mSkqnGJUVvO0
cAX5qYMoZ1EhG5CdiEL6trJJahZTstSgObhKiAPVVdAPX+1Rv6ArUuHzw1RXNhZKQwiLyKkZRYXf
Hm+8gYH/WCJpVFHlqQYdqAWimn9owAmnYN10a1VWnj/Gsdz/oiqAx/br0QWCeCK+AnNBUeJiI5EW
SndXuWhVz88y8B33OERXnvPZOOz+mWSw51i8T9qqHkHFxzGFDDWAJzy37YDR+Ezg1wQZY9UMw0gr
RVJvuc6yRGip/na+/wb0BykeQxrt+ddjmL896tpML5bzV/ewHlxgJ5CSB7afVS8iSZOO7v8Xg1vA
JeFNi2/L3Bi9JWBJsJftuHS6g7U7fqlq5K1QbW0nvFxU9to04Fs4h8ArEn061f1H/M2eHKoI+ORS
Jcp0kqd2uKVnAFOp9Y16BKsGKVNJ0GSDzI7wsEey4duja3RMnoV4JBiOBOg22aXiAA5kqxk0n4Uj
taKGEn8ZYsjrBPuXOiUg7qM4EStXYs4ZMLjy4pu0x/whN/I2hfvGIV8dDareIDWiH48S0RceIfjb
a5EKr4tOU6pvhLbYTf6I2RLLvxsZdLLg6ozbG9yv6h5j22ShQeGrtuTmZ0R6EGpK2HqEDM/ehfRL
F7H8FmrcCjn+kn8A4EtjFYxZLkK31AED1dgsJqDNtsDGDVIDqarpOWeqUh6nlcsqF1jFg1CGaayl
pUpuv5s7EBuVOkZEAQna5M3xyuF0iKTOPmZYrs8zUQy1vkBF5aQ27YM+DBwdv8znH2gIdwx0ox7H
OBO7nM+oy3IDMC5WeaQ3F9x6AhT+B7uS7BpraPbrxVPJmMjDWkd6fp+R45hjPWvs3KWYojv7stTR
7P2loVgX2BIrl+bclUcH4tTKEDSenClB6ChFn5yfKkL8kSwZ/sum99hBapwHrePjzO75sWpbzwk2
RwGNXMuS5SvuZzduVmMg3290tlx3dW5TXzCrbK3LyBhmJ1VHxkarARyq+uJGTMkoa+JcdayUepEB
xZTLx3kcyXttoQimlH1XfIOxLs6l/nL0WyICRNWFaajE3ExMRIqE9ORh9TqShar6Z5F7s+m3urq2
vOCRjc204Ei+qugu0ZZEmsP++JBMUyryDiTfO1kyctCr/UDxfL2mrQcfvJu+IZCFOyrCVRh2JrvM
bNHpDdb1IXQ/mkWMTPJPj/YEEXTymLajkPMs/qfKfoge5c/rDRQd4av7yYAmR7NPzIU5uEMqncPq
+Tlcq+CAoLOHzQfjhS/6uUeEHkMgKGX4lCqp1PD9TN9YAUcpZ/Lk7cPLlJ4TvKBMhBkJKdg9dlBR
gkwqS735XGBIQ+mrFs7yDQxqSOtLErwwYb+U2NfrbpECoS2I6ugvexwsDtdkQAC2FmIWvR98X2uy
TdCPt8DxT32nhKvPv+QZI9mFUdB2M4qytLILr5bisbVzd0TknQI+HF/X01xS94o+iNJ+jcHhthk/
VFjoOXLH4O9/+NLnfhKGl789nvSd86TbIHap9IiCrAz9dATpTKurvB7ClhPfP80LEfu34FxMWAmO
82ypWPO9ddAqMMo96mrTYtSSvI9fCoeUkNmc1DOQaGpVEWFUc2EYyldToFi18d+l14ANxGPq3Szq
RyYC7vswc2x0m9FQ3PQ2AU+KEGcHPJRo34fATq7paEXG9tcjNWW3vGMblbXHNlprU7AXM2Du42Ct
jXoqCg98eK09tz4uNEUcseISihwITN/79QEt3FlLFrvdwUqP2rTPrt6VcpQLcOeWmJ994lDd1YTV
Rw+PyqBl/KAL4cm2LTKo5Qmbb1pq2F/qTBUEDxFUgzOeGBCE+K9jp3D3wxv7gwi/g5ijCTnOM9iL
HgfuQwzf+egbb3n7Jb4yopicMxysIkb80yrs6mkmP4zS4CJOrPIfItCL/Kg9NaO12ZRLCxdwVFIu
QjtoINVOTwx8cUHNNYqYEq+gvHSF2sD1fGZFS0t7FPP3alNaaNjgr3iBCHUA1MEkmAFY/Pp2hSpZ
nhnVOV+uMDrMeYuu2IX/lkSvbgTe/JMNcu/Ha6GIOZHY/HF0ZmTWiuCN7ILsrmBOK22UIRZFi5+p
k8BB3HtrVx3X5/e0F+fX/UvxELapPKGZv7esAFJe3cg4lNHZVMM348x0jqDL1FIMi1mPQyMCg29u
Bn9/pbY5bmDuvDGKJPiTo/BWKEVQzws4Q0eOWKZIeUkjh7i6oufUOA+1fkAZQUXKrFzzF1r+EYaF
RxePxWabBQ9HSlgRGWK4X2cJdsTBbQFvb8eKsX5ZVlqSkFbAHjMomntUhgbRMYEpoSgYo6egpUZG
uvmdEMB7PaLOnyz0aCHeEulW8pTWemgs3zcNd5b/W+AI8YPWHfuHBCrP1eV1mPOQT+2JS0iXJrGu
NoVI1raa+ZMKDzFfI0v4Szp0kNXxbly+al60HeODvzweeiEXXzPJ9N2pLZkDdYgvKcvCmyBhD8Wz
GPhv19qBFX8am38sI44CvK8ryK8Tl7ILZShFsb0Cvv9QOkNt6dFgA3Kugqp43/Z3K/0v2foQyYl+
6P9gBTCX7tskQjTLwnexnila+nF0ez4c87WIGtdNg3dw8nh9n+z1WSCy5RPRaFl+7UyDtefs0yUW
h1p5HMUlwONXBgtz74Kbg1CRKVJeY+DB+ZE4WK/WswG1v4wQ+7oozu5F/3wJYR36qceprZH2hCG2
QQcTJsD0yJTCGbfRXnobuWNtSkPSW8kmRYfCOCUeEkGmDIQmdMnYqz7TlfMRmAEIQ46eY+NDXCzI
tLAC4o8NtLXsGCpOygXlavn78cLHDZkyQjVr9GoG3q2gRlBHRrnhFzrqhXmgW+0cxGuBeNvb4JNH
jBQQ450hOP+2/+2ol9c2oOIdlMbNJmQpPuRwMRzwaiAkNg0Jb5BOuU4eNJp/rm7wU4nSGP9BtLG8
XTLi+ZbHJVDvSvzyvt22uoc2NW6PbNqBoLDlKnxLn6rmwRSwJBiHachphDbWTZ6Bvm3rLk2tBAQp
AK2U6ZfQLoNvHev8zi5/0LNNvsM2d2pDy2hGU5WUTbb3ACk7dSv/Nh4NdW0qs2+IpwZoHiVP0cI7
EuSzK7jak5atm1Hh9oo+rAb065VnNAgVfDbUiOBhNjsku9rmqmTyixGscVBsYa95N7eX/DxgRfbg
voxlDrapVR4SnIGCAEzLLHR6FEXnXuBJGrZwbSlZ1jXKPaIRVADzWXwpmhQHy/jZg2PPpgTnv/cD
8zKOhrH01Ib+RATaVqwVA1I19mb0nvTmNqIAniz/H8zOtstVdGrBWxbDPA1G3ZiNatxsu2imfGZn
2jP+g+YTzS2ANCELW9lPq1LJqn6v9kgqvESv9RU2E9aphHxjK2kWcBjzKDvM+yD4U7OnReYRjj9X
g0x6QEd1gpmRLqpliVPhp5bgCR2gw8s/ZWeo9lWMAL/JtWP07drXTnGl0sWM2dK0MunMu/HXrNzR
wkisu3H0PEvXQiFHIkEFGgxeSzFqHBGuTmv3oeAIHiDDtJK7UGqkOzi+hxqo+GXOi2vS1SeD4Z/E
+Je1MFoeDRN6g+YSP8ifNgYORVJfipRUmzdrrtm+11AtyaUn3cs7Mwx6Fw9esKopxMtme1DivROS
zebmAgy91e/T1XfyyNVznx//sW7Icqs8BnpZz2B/bHM6k/+089XUQKDWTuG+JG5Snb1rTrUZooJA
REtkBABvJ4Ljq5rudzm3n9kYK0VrVTEEnRc7iiHvzVrTts/QR1Zk4qTTdMtkVfyjV1kpP2fyT67u
5EWSPBwFjix7ad5eu6h5GjJ58GgxkPqJSuhP3XjP2T+LhW7GH3NduQgWE37CqFF3Ud8T/854ADI+
s/NTMyWuZQ5s2E4Jb+iqI1lNfRQpmDoZQT2Ud96xKSjDoThmz9rq5xRyFZlP/I+rNLziCnm4GPT/
I/mSaI37hB5AsoYGn1DxA4uUauN9BszmlvVgldeWGbpUPEjV+p9uTOqcHUNNVIdlfCR6r6jhucnp
9qbWNhxFA10klgFgeMCdE87ZJ18HDHJ8sQXaW/QO3gxIvUipKidn9Wmraqyf464ZMgui/X2NXa8L
E0XBC5jtO5uVWUGh4tQSRsxQPP77sD76CUVqlSpJlvT43WPKXPpGe9L+vPZ2a4DO0fJLXNzbccd/
BpHDbSMBpfhL1ery1AKNRQqPiQyhVQdbAgk0sl8GyNPbBOXMc+Fq9UsblM/oh845tiqbA9Bi/SHb
UTaRAcx4neswbw3iorReNqF6oykd7qlsinIA6eR8vLe/AslNub54MD603CbZUqbQdFbENzdVgZGe
vhd2AUM914TauQMcjyKe/apvSXhMfzVMg5MGL9afSP+VBFx7rx9VKAEjErFJphjrj7YTtPTw/Paw
YD6zIMjMhBM5aWuEj9zl601OYJdAfl6dH9ZesjRvgPZxVnSMDw9fzG73XCfLDLWoFfFcpjXManVY
WLZZBV/aNuY73pRwxtmrDt9DJKCz5MqL9RSeXWZpjJWNReLrh7mcSmsrzTXdDCkH13lDN2xPYmsr
umZRErMP3ck5YHS650jjvWcfcfylbZefO6rL9wgs8+Kifr2AqXX3pGRV2dhrLstmULs3wLsfYbb/
KDfVvqGKfndVLldEc04k1HMgOWzJGYKl16AFX18lDufC+v2RDlORXuSb+9+xTKeZ1NrNswtW2lkv
x7cZNcAsGId0m8Ov+WFeZGdMrihZkSMQu026LCoO88zb4JSnp8C0b2w62lXuEDRP8JBYPwukiKAL
VOCQVhsGtxIMe1mimKcsgIpa0ayi5iy9e1QazfViLLon962qjwkf7rwEWeA0lKplW407aELRIfqQ
AO2ZCctdGcJiAT5BcgKQcPaEjSTFPeScc5JWukeyJkHLU0hyTu+wGk8siOaMXGpvTL3ML6Nd0dwF
w1NtyTaMl5BB+Jyj7fyMex/E7qfi5+auO58ebDQ8ijwVZvNbD861k05b2VmMVE53B7zblxrSXakp
wyEpDYTYFgvJWPy6uA6dGkf+z5wLwOR2C4hpyYytb5uKjrPSs97BWKMab4GsGsY2hBwJDd8jGny0
/InEXvfSLHmqiavbDGDCLX/mWtOK+132m8MqPM8Q4ApVHhirWDjPn9WuoS57GnXd8HP7KJFuNooT
5bGzR4Pl2/QipdJTfSoeEpVY59jQrmuKVogvfxIlbCHuqej6DjFgrtj7Lh3bz/oJK9387cWSuSjL
Voyb0kY0oP4ByZA42kjXR+CpmdcYQ6mgGzd6A8EuUNeUcfqE4YKKarBZYC0KrIddC1bBW6qY6wxq
074UejYVaB89Bes5TNlI6fwhMHFuRGVOZcdM8k1TWYS+yBkZBzvAqVLAkb8xdLeXMKfH4waw55zh
oG2xHn49f0uNKrO7l4TFCg13trjES8F6gv5hvSboMlceLn+CGNYylPNrEAahYKm56f1hCuGVXbm8
vP8dYG+GFN+xj1Wv4d+grZcdCg1PBElPQ12RMzmxp62Qogs5KPdb7eYB9I1XP4NlA0aelz7FhkOo
dcXh8iyV7wt0nPQJ6UGri4z+IVpDxjj1judesDkqL6w93IwD9vbcBtzmfkA6/q0oSqLa/gvEc2X5
TLFlCN9g6ZoPPyrecZsTyHHTfzxgb/TUjgloqkV/fAeAmCo4UZjBhfcjL3eqr3x2Hn/809wpYDgl
7G0NsWzz85USF4AGzy2r0/ACTptwuXppXaxmC3vDfIHnQtOJO9SbFVdWx47pFuBsrZmtynLGOk+g
Gl1bScVTvXJyBKz7LobVLWjQCyRlPPc/fvi1BwA1WvPErUJgZfcM1dGbicpWTEozV1enwqYVS5Wv
1xwdXY0mU/sUgLdzWFdtotrrIcGPxM59YX6D5boeBVARNtk7kyzwqhph145fV9DtWDLu6v+sjTR5
AQNYq55QD3N6OCamNqNkc7VX8mgFxLRPwDxlgbpQTn08z+/7B/1YKbs9eSr6yzmVBpxV25RRzsex
vWGkAFS5DEOhcq2V5+3db8V5tLsd6fbeWiGmH8CoL2LoyYTAoKIFolC945DgyzCT/BcpFMSDrMAF
6F+RvL7Z9vk3bkxbRwuUs1vi+jJ8bXASMBjQT25NfwMl2iw5KnXjvN7+KjuZn0z2DBZC7np5b2Qw
NBsTGXsOByeg3II/SxKWthrEiXokuXN1Z47AyJKzj5dlGCeqzR5URja59k/DkxPS69hJMrJokJTL
9t33gyvzXEFZJILCUHMbyCNlH557bT15A9szfzAZhy+cjwB9Dp8uGr+ialMcUPSuMidt0beRitbC
chrjQAwojcEjw2Do7+KD1ScPa2ZESPq4TdqpMYNQj+rnKfnn0LLdaTA2KhmAH5JwcZQd4MtpVfte
yk34j2SusGMFM944u89rO+zuixefEgz7yC3jJO/Y+HWIUfh262AVu9HcVrClLQuSY5v4qGsYkbTr
zNOF6M53m3/a8kkJWlOlI5DauGHTQGsl/Wrv14vOr6G40xLv5CMjYflpACXjP1WsLTAnJz4Z89xI
o5IxhC6KI+6D/JdGqc0UaAYMU7DEqn9JLNXXru43WklnG0IJYO4ioRaUoMMtcJawWbfE7uSEVJqX
pXoZ2HE+xLww86ges9h7ByL/5p41ctBYll6s/TPzc7t2WrAFXd9eQ4PLm8RMUmV6qkZHgy2RGApy
n4ZVaUkmCFB6jcu9H4i8dRF0+nxKcXFc1tQtEfLhGEkL/LgCPKmR2xwkSmFLxACHzN/A1FvQU2wW
bpDmxUd1U6SH/47e13zl1GbzP0wFmuCKHeqasStwO2AccVM4FssIImM4Xg//rEueQkPV3KgEBn9V
MtAy5eiKjJi0jOMC9SRK1+7P0KuGque7s5Uib7I+UDL0BGCnyxa3Rm64cgFeZmvlBSEtRKTg01+g
WJcnfzYqwrbMK1WI0JB7dWkK+r0lFaBHfUd5jLWg+V+KXHRxJZVPnJLLMRFk5g8Q9QipvuRKTGaa
tNOM877Jp1YbO7RfLbTTM/qNDeqC1cB4N3T1Z+8lLvdRrPMUlA8A/GcMWQ3ESmYiRjAP9eZEI+IA
abRFqCORqlqesjSEqanW4dpgU65YjxTpzzd0H+nlhYnkzIXSkAVsoFS1EHt1yMDuUDoDUgortLL9
nkeGRk6nDtGxXTMdE0TqOsEvmG8NDe9Y+N/aji/duOOnpUZYaRT+3tWUvtVldIVfmZXDOGYaOAcn
w/EY5BwQ6ZVVMTfuc+YDHBYAw6HdHA+t8YgljUwPkXVFDpLTnNL/j+HBRdo22MYwCZuBkQ3qSwtG
wY1jZn8IMlq/c/z6YEK86y37bL+JPERcAgOIC15v9lO2gQr1Y/zSZZzM2gCsgdRVnpZ7MTDjiW7B
9Kx6hEfebLgf7/naQ6BckGrxhF01qDHx+HRkg9yb2OTCeA3yyVJje35uwNJFjch4/L2VO4bh7DvY
8iY6kqTNtFS9wJddx/zrvlegonXI+hoAeQIZSiFkChO+uNCB2ew49qffONBDfYnSEca56cyYF9iC
Llcog8Qkwjv5GY/UvnkWgvf9zWtDO6//fpkCBQYO6in/Y7N7V5fAkVTHHlfBXuiwzrvtsJWYjgxS
m0PtaObPN/q4NGgopT+11zyZf6o4Vbr+L18TeaTYV/vz7f/QvBJfs6t07zxaId5XcL+hz45cTEnG
stSgeOYuUQjtehllr1alyA4cz59jDZU4AI6MM82Q7Yn1YVR8izl48SLFS51YcgJmjc1swmiXqW2V
bEFBcpzW9uU/5XOj6Lt88S6LWCfkBH1lbUfFmH9tlwxPoJoMM54SoW25Opf+Xxunx3irxs4/sL82
mdDoK9vAyf4LNoDm7qdJgRcwA0asdIJsUlUtsbLc2Ycx5W58exGmkooHJ9jlR0G2TTvbYvjS9knI
TcjINR3xI85nkWpVcQ9lZeh3muq+32HqVB1LfFz90CeTZGDxmIGinj3/1+jmd8se4/qCxW4t8cak
VJ1s/ZAbRLOP95BPmfZI9Pz7tI2ofraEmeuPR8bV1b1N40xpdl6p33HNplETrJ8oNxScakywoVih
TbjM+Ifg1amsLISrtjzBwbOROSfoAcRS/Bh73k0MhmqzMS2Vfb/vlLL1IgBLQ6GOwdq/8v7raYoh
V1EnrD4JO/VUxsyUMCq3PWIZQ2ke3VVKU5L8JP7morSRG+akgZxxrUKJkIQx31aBLM5HsaE0wTTj
AhTrctkgHv8UWgnIaKaPcBYPuLI5ejgfK8saOpFT/igfDwfpHr1hz5ce3W+9ExpZVa9Z2J2qdwLs
CYr0aodqcU7Ks8X17RuqYtTmCtQXEKcZXpzZZraHin0PXyiPfnVHew/3vdn9B9uBFXRbg1Cre4TF
YPlk5sC7PySbC4JROsFBQJCKyt3+6ekKsibS+B+AxgPFNZ9Ig7PagvKy8iLPdEitOdO10KY5tn0r
88eARjRUFxC+9b6yXOCeR5YFYmYgDQFYUYfB2sWY6ttUb54PYHTPuY0O5YLKH0Gc3JMRtTzgEdqR
K5DFRJfoPChxkbU9GXOMcCxYw5rGzrj9S+Ss4c4LoWBHpnPTtPLW8XDhoudovfyNMQmit0AqRdmL
G3qCKjrg2Fgs8ZMWVorZPCJOeX37vE3y/tetje/lKA2eJSM95sg2GEYzg7wWOchPUu6turAjjDd5
qHpqglJkXa9NiKY+0Mv8k6SYJCSRs0SBMeff82R9kekTorIrFyMolC4sS12mBWIIaCbgw/25NdBe
v7RZt0NIL7SseiMSAG2CEU3z8q6qax6MacJ1DT8toytkCVur5PhyURx680+i0ywC6AuMMSx3TFl6
2ZcyHPI9+909Rfcc1gEOB7CRNI239yJK9N549m/agSNmupqeSk7h5jiyGNaVIdNCgezyCWiurCa/
qeD8BQuCbAc+P479I2coeYbvCG5HvYpdC2taYCgACetuhenehba7yEIB9Q73oExo3keV2dRNZbF5
Ccik2sqRW0tmRPx3mpXIDb4V9MD1aRyPn8jAE7IxeLFPi2kTwMIK6lT6rVlIX0eLwlgnuWuw7nWb
IHeJr+5PIZQnA9jjF2Cu8URxc3zwTWK3QIvu5j0w3SneqXPxTFJg56zKHskuCbnNmfD29im7Y/Q2
UDts4SD9xdFl4Vbaiyes95PrAorg1CNReVnBhYaYS7jW5KC5ctbyfAKQuEp3fHe/PoMnTYvqHRaU
q+6VaS5wszYbOECvnA1Hk9Kf+85/ipmWrbmqP3kKVGz6Kepk0ji8zijaLDcfvhfdk1j/iS4MPdGA
UZabYTZHW6J7ky2sMWQA9t/K7CsQS8CIKo0IpIrFuCfjDIa1IDiYJEkxCw0M9JkgBYO5769OQhQ8
x1Yfr5rrgy6YNUXyw67tQ568w+gb5e3c8jhUvJNau+jpYtqWv3/jptlAAj+y7EBni8lTKaIKwkFW
GGlN8MYkcitkTCmUylwHnBJq/Iq1TbjNPG9ABXMB5pItRfUDBjmcmLTFI4Jv7QeYExK67vewiN7k
VwFIJK+Wbo+NegWwtP/3MdF6cxnre7K6o/Qfaaq0Eo7vdY+7xaY62VQao4cHS/WO4bKOggrioQRc
XgcrTx0FzzNjTPsvWSGjhTWyjn6lu0AFa2aP/qIcZB0kWTj9aPcBZZA+7bQQYuOUlqujngAC3imz
OgRQcJmT587XbrWAfvqxiNcbG20XZaGWa7MobuK6jSLdwdYi8SEkqdzkPrWIACqVV486hf5yTOmK
C40GEtdtj0jyRCFxotmoslbJ5j8ZqiEj94IfTVze2p7hg063Zlsoj+tUnp/gTnWG1D+ul8YM+Dr3
3mHS4rI9iJn+Jkypi+diklJU4hNjAKqnR6eIF9HRMStn2V31n7rL2uu9vos4+RfTjCispF7MKt3f
Pu66W12q1TD21m2L7YVJ2oPKer5NASgydFjnyBH1KFoclePLvuGHlc4MwhLzhnWOyRWrMQQebWsp
Ne33odjeBuNqZCBLJiALFeRlA5dp4MILbYrOrXJ3TOcH4RTDOsZj1A3XV5QMb7BpiuErDbriMbeB
Fzq6pZxLdvF9A9K3eMq8WFnSXwN+MRxhl6yL5gJVeqGDGgL1oBegA9GxzNYu/BgD4pTPQdsQ77r3
pzeLhzpyf9HFOrpTA/jB4uetuvrgUojgqd0lAMcNo8yDGcaMOFoAwzuuhvVJtQxP/oVDgUPcd1wn
HRIcniS57w0ZdZVe33no8GJsdt/POU+uZF/Oco4fmsHNrS7srxa4KW19gaoUXm0YisUI2BW6fN1J
7ZRwbtNVYyPp2FsZQRzijw6g3e2nD8ut14t1i4mSVjSELh78dARkZO2N7Zsr9wptc32L+zUG7bp8
N5CClQMJ0BOkhNbpWT4f5c73AMmTdIHR4zv0K4gwY0KZjnl45VAeRCD4B6CCt+b0ElIbcz0trFjc
wEepOLJNFPN/mNnfP6WLuODoZ4++M6YTJk9qLOe5HBKVyTBFBR5MAk5WeHRVEV+9kuDeUeVMX8h3
aJrfFMcZCNF3e4VALH54bOkv+7ipdJez+MLgG7Jyc0EPaKUf1v92Vr/TvuSpuTI3Z2cuiZAXHdek
kq8evltRY1GHx9kpZxA844BE4+4WuW3JtMbzYxFilLZ+bh3ygztuWDlNDY9LKO0aMRpeEHpsNt3I
I7C7JbJpYdBDYQe22G8Pec4oWBsoTmSgM3TZn3YDmtA5FGooOU65DRvPq1AAQ6IcBxP4VSFVtJUM
1rRJ3mXgNXpghbAHyjH6DkfuAHpbZA3xpZUj5qHWBDVP5C/3ctAFURtDZ+AdBB1JDxKZuafgNNfh
fxkazahapGxUdle94RfAWjSd/l0A4roq+2EW9OQApAUp1oYknz5Tl8Cwb4ug4cMd+yx0jdRcWio6
4OIZb0HTjZeL4Vp9oV/lgWbrv3XLafTzSHEGqSPo0MqxgAT1krnG64BfW1EP1N7Ve+MTdF517j4m
Odr/1eQ2jXwZKvCM/WoE7EiNbkYmsFmqhW8s1XN3UAgznRGR+VAuWO7slRpTfCxaIFvvQ2G3wPNc
dQlkMA0iBvIZ9e7MhpDPlXb1s3Brmol77E/fWwVqnYMXfSE5+4jwr/q4s3Hr6ZgSY0F7n8ErxrdU
BBQhDXAB4w++alhLwqXji470Bx+HGQLoMKOWhud2t8EwPs9nEREpPrR3OgL1s80u9fyL4PgpVvK7
3x8DKBGnq6/UdgbsY2ZCNP4un6h9nOdGPQtJl1TrI41kF/TV6oLxAu10HBkTKfbbUwHlR9rPaEF3
xE6qA5W7sdTmel4Z1l5XArVS04NUlaB1nfq6p2/QanKRn00ZG9sQvMEYwwxIL1sDUizmm/6NIZgJ
VFdxU4lK9fezbi7Fp7u5CKS3iYsUd5MO3eIjwLKdPeMv31vNDvkx849IgoNqVMuQin10BDThDYGB
JTzHy/ZI1svMIdfzwB5A3QVHGKeLpd8kR9bQXL2xfcHZ0bVrNmPMPaqQA9lSnHNBRSI+scuRnvIt
m6XmG4l2Uh4Gl6AxQZBqtmVa6flFh8bQRip9nAi1Ylf9f0UHRGfFPR/yAjHfSEVPflZf6iP6PAKj
VK8gVK+gqNvoDJl1gW0I3uRe25HYv++ZDjUAzYtFLChW5EiRjmC8nInBEUUGWTCUuA6A6815rdZ6
uliMjrlwDdR+woKveSssFKl9QEsy+K3LYLQL9pEw2/qsLoviXiRZbD3F+CREQSVSOHt/kMp7iKgN
adp01Axg3AuXNe11qwU4AEfXt3s+EB/X9oUI7Cy51Vh021OSsBM8GyVArabi//SVfc0gk2eCM6Vs
XvvQhFRXd05eIDi1EQaVdYkRvs4H3gnYOCoiyxxz9+5nKZ08klPhb6HA8omNguN8/JE275S8Q5jw
KheDcIF2QD4FKK2d/6v+XONmOgn+rHxNicVHr26Area2XoM563TtiLDd1J7wiBA3zDzuNc9LCM1T
0pNkpeVRBfd5ln/FlS5yYV+2/HsgiPoAvCjEKibWgHvRhajHU61qK/9qUmm8V2fwT5vz2Fppq+2/
LCXaAB3wIYxvrfmybCKQEvdTQ5P6qeIq1bfktMn1mHtiQEkdcVlYWrjHY8+C9qpOaudW1XYvDNCx
1Sh6pb3aQvzzccdiJGwzfFt3VSV+0OVXr9AQojdD01NZA5twE164+fj54etumU/1RsbLYNC8vm7r
0/jmRnB7MEawQbECj8N8VHmn8AILBDNsHDCLaCBhfeAqkX2meUTJWgNyORkR02CsBcUMMegRLMV3
woxj0k7NYtjxv6JWgKVGRpZlQJHtE4lhpvh/tHkYt8KTOWPqwK3RfwnUO4B1ow2jksQbJrE3srPQ
v4oF99QfDm/nKntnWJ8aCJ6fSIJMDaLRxjvxwELIyMITclWZrEnSyrFBbYv8LQg0pC8iZ4+8saut
6/7ifczlGbt0t3dwIaT9XqajcODfp026+G3UamuLJnf9u2oc88jGjYVQ8BrZzSO8rjhn9jg9BEA3
wYXn+KII+p71twgbegpC4XseNoYNBjnrvcbTqXF93QwEQtmlKc5fz8kh8ChlBop47DdxKtBx7gy9
77xYsta+UKHEvNYr9h7/TxbxWA2MGrLSDoNcPbCbxj4FON64mMY9LPo0SI2NXsNPwl2Oz9z+PlIJ
qnZGQ4YhoZSuMTc8RvMRWjXfSaGI7njjX3fQH2iF7wCAaSbjz5qmIRKWs8vySXyDJ1uHcZXavJoy
ubMUkdGK1mKofVegQR3Ugd0kWEzf7hNHT2LJzS2TJgmxrwqivHz+0hyJcGfMsjDLGjgY05Sjl5Lz
LmV8hmdwboCzTQuSzvaUPk6ey+D66CMq0xs8AedSilR6ZObtFyUUpsx5tt9+DqduXtrDyWFSF8Y0
CjwOH+vejbRqtP1KKaEehsrKld/iDV/vRm2OlIH+0EuMNSCl4w9FlUP7W/5N216PE4gsAwbIW5xe
BM4NF0SjWK4ocGIW7qHTINWbUfv4Lvr4ZjMveQSpOFjW6kREVM4YIbKSAYBIBCFSy/cEABZgFXuc
VqkmV/+j3cBEZ+UOJCMpuOL4XMitCulUbP9S2bWutPKvFrQnE3SxRFx0S6p6CrjKdsSitXn7ezpZ
2RoxxVxDl4dfijn60yfPMr7pj6UJ2XEJUNSTYs/L6v4+nK9/mnl8BQ4fEKa/KKHgZ5JIjl2RfOZf
kxIskttKjppEiguIiUSb5bgnjLc7HVSMgSrWLZnAqCdsV63XTHDykx4DN2IVPN4mRto119Z2ID6L
40JEuHVI3Go7rj9/MdiPmrkRGN1tfqHbEsmtFgOEEco5RDO7Q+UXkFL62d1HibsuxVd1I0FQrFom
waZokypPY7Ya4/VCVUHVCfjn4Hks+mI+LgaQir7gedANAtBXfz45nimMcajqDJGEUqGJ9CAOb/HE
gNXV+cHvPuSiof2Tg0UBLqRFmWBdfwQb1dZLih80kC9Su0j/4ZxrvuKklk9HVPNJI4G3tNGnFw/Z
eRkV3J/7j3s33ziXSRAVDVcmI5yQO8Kb1Z5TTjgXElHUxsSjmazSKUw+l/R7uyMsYmgov6AW7MyF
C3a3+pqsKBRnmKAaGKZJyqZgcOM79AQsMUEm7QNYdtElEZ7H7S9DmU/42eGlddHAPXRxa3aHMyIb
RwAovuvWAPn3lOi4EUtscgtlS5nr0EozbFbZdANB6XHrUqGrF7Qgeu+YliKXTsODY98tuhg9v36x
jMKjXatkwr3fR0/WGX/xMY/DA/NVm9K5mwyAcfFVXuh9grAw6amBDOegtFIaCHpLGYcnJT8UqxJs
8jEB9+/YNWvq62hAvc9Z5HCJlkmpjw3dElnUl4HjbA9ug7vK6jL0NetNLA/etYu3ZQrJ6QXQjbY/
GhF3SfdoqWC33tAbCPVlHanLNgXqnod2x6jtidot4hojMiqcHDZOcYRvpzY2JyomO6ZR2AIeqHeY
A0n8FrBkoDMRhS5uIfVeYryyH7rhWHO7h67/NV3zd8TOvPNDdeo5fFsjjNoC2amEvAeGMj3NqA7D
2Jk0tBrw8DaD7nicX8MhI37M6Dx6q+Erme8ZpYujhp9vnPDYO+EKA9DuJLkSfRWVKqgfPGFIluXu
EZtrzCUkjF0XxzXHL5NLLCnm32DcVKxfDZIOlcxsTkBHvYHBCi5VpOGkhXJichk+C4gwN1vqHW61
ATUd61y3FFxYZf6jNGwYt+17abcudnRkap6KJESkBoEgywxbiZ4TZZkSlSPneLJH2GcaE4Pp1O2I
u1srOsyTsxOFZbkslwNgsl2e/cq8cmg9T2WzFnWryR9n283UOtuzHC5jQalgUko9P3oVz0Ru/pQ7
i2P1cHHs0OjL9qOf7A2E4ArPO+XqhpZubOF26dC+saLirENqs0Uk2ne8GvHsoHjVv8kU+ADjf0UQ
S5dWx2J8cY+E2wPu/uG/ZtuVyW4WF46BByS9Jr0k7i3pqIO4pBklMJYpzIoU0baJprwd/a09MYzq
+mhz6lNFIFzXTi1HWk701AZz43xzlohDkye4j5ETcceXlrjOZF53S4VA+gprlgWzHePAQOQbD9f7
nTGPvkLRDndR97lIlklFijw2/neaVr+r4OpVO/qFltqhKI7sLlPhTyZ84F6cBk3h0QhEkik+3S7k
nhp4DvL5jZ7rAxVv0eAFnpPSQuFHbZFj3WnchjsZ6HbkW5kgub7gmTlJRgF+u8MgeHeQYuCmExNs
Ze0uqNy3VGh6CVq2/xcIhBAmbbKx2Lp6xDmB2mEzcQfDx2l+OphM4aDbMupsL5Yb8knApQDbTTgB
jJhLzBO8FBX/COnr3Fj+GfpX2sJQeq/lpm4UUZReypa9nnGMGvGLlPScaPGVeLo6Xhk8s7ksZ7bI
OkcaqBQJWHSsQARtG8nrA5yESzNPc5pTGknK8ADXLguWFChDUs15X7JJfYgEuxA4nZ30pCJkgRfB
NShQMotDgrdx/aOhsREpqqdm6Ti7+pm6TSUK2d6dAYfQ7ix5Hm1FSJoNe5m2/JJZKrtPNnKmSBr2
c7gQOHHoYf3FWYjKVz+x1CYgXAE210pyqC590RXnx82XWmSolpCw1155hC625eIQiQAliuHRc+gV
txf3R8AMtQz3Tdzk+kz8MZXm4pvf26nM9k6Xc90qLjfgeBoAhQd1C3myGAmGpXJF1ys3sZr+IlYf
x0MVgLiVCTjXxv8h+1TvtbSUbHsKgrAyGj9ErYUnpIJ8Hx17Ww0YN/PWzpTHX9XSrUvY83wCKo7d
Ee/8oyLs14WCxx3b1t8ATsBpOcc1WJKbg+uVs8nv58OengqonQ3Tj3ngaX5jOmqUpvPL4xkOanpA
MMbUu4fzsQttA4d3BxMeLX8zX5vosCrOIIdFc32gnD5PO/aiJeXni5rUS6WNnv9dk0skbHbbVGkX
+EeWEY/LXarHrYE++4qgDqH9nsgV7R5FNAM4gb5M6KxT7BXUVVdX7FuolbN1+icHjstAd5mPvy6U
/MnY+kjnt5k/IwxEcgr/19GaswveNGvZ9PffonkMVCFCH5Ngn0UIZf/sQ0mh2y0+TAkssUOeIX8f
nV+/2lIQb98oQ6XBfbTcVsxfegoFMghy4n/GsySpw3t3xCgTRlfnuka4tRGVi9sUgYJ1Fd2MqGRM
FHod4NbuMUBAhwEeMawKgfWlp6UG4fwii1BHmkBq7IxFc/9rZJCHwFDtDsS3MNI2MP7Ryf9Lp38A
zZpG45OpVTlb8fGfqkob7m2cttBMn4eHbtQIlAJD2437Jbzpi4vINyGAItsXyFMopSPaLmwzfMKC
2jg0C9REivmj+VHJHQGaX/k3nYIcHFetolwg1Tz3B+Q5/Th0lL5lfWyNEq7CpmYdudTGhs+Igo3G
POVosMA5xVU8YxsZYRTXOcusPm4QG10X4c+qRNNAPNnHeIR9Nryc+P3RsEJOO7rNLM3a+0MKCs4I
GB6xRP5uBgDBc/qPd03Pj8U1V6vSK3CwWXRcrmHN+zPc378S5ICzb7Fefqxt/gd7z5a+9VeHOWIL
FxQXxrxErQ/za66mvX45qMxgY4ssj4yGhjuPMh4l7IZpxVkpxPAAIUypX13u8myFQIHLshV23Bae
b1WZuey9VnXZtxh0scM/vODieWLrtrT1e8dTfJsjn1BO1eOq0LLcUP2OgeKLyAaGP4h7LJNjKmxo
E8+BIEshovuXLj8qBwh9UkTBcZzc2DTwt2++KmdmV8YEW4khAh0Mwb4VF7kqQS2KIknsRBbBia5s
2sDeDid5C+sn1LDoGw/+yaAHvqVFH8zZq1p20dq5fd2GWyEidJV9KvXAVAD4UPr6kLGF4q3diFa4
OApiKflI/9deYcYnX4j3JAvLUiVzKd5gFs+fz74NsdhG5Hyc1hkNDZJdgLjIQsIr5dxBxST92px5
aZ8CNrjmUjZ7YpuUTN/jCCD3tjZbq8zAvse6d7+YVZpPI3QjR1BkxIe6+8t+s7bMOPl59OGQjoBQ
bdB4je8QctBKW4BwPxF6yGtvMivnAzRjcocDeCr2Ud16+y7x8bCZVYU27XbKvlrlSe67hEm436gt
6G9HVTer+LnKA0rwxm6BCfceutWDHPUCDnuczVDzoeLiOFI3RqkL89+xGwFqn75JkaSKx8NtrgFF
Aqy1qvwUer1T2Ve/kHUxHNN9jYdrhmiuDqTTIdG5Y6AzAHFe//hHeqt5KBebaCvpCFXKIX4vGJGx
Kn9GTNNTQw3w52F4Pb3H7QSz0OXLMWAWGkwUenFphDQqqcUQBiJpiD7KNUjaXQdgctM7E0IhDpAf
n1TQema+SwA9BObxyJiDwegQ39N4hbX+p03zh47zW+fJdy4eYlWVdM2V4F6y8GE3mRQvIhlrFRW1
uZQX/AD/bi1alhyrMQNqVFpqtks8k903nLZVlMPDZKx1+883PeH37OQH+SXuVfq1R64zPHu3QDfV
j67W39CY8BABvQhskrEDyrRX4vR8hGzgO+N6OvaBm+G4WRmYCzWO00lRqc0+RPXTHSgWaDL9s9O9
fdOduexkLwSu2J9WfYrbUOk5XMhXMeS0FaNEZsFT0E1pGevqx720FRjgSv9MDwQBSrFXw59PK1qC
xit/NGJhpxpmkvzw0OjIidarjmnzwvk3FQwHerr4W12ZwO3bhMBX32WuFJDknTAL3CLZOFCrvDwW
bmosmdbpUhb5iN0yxdrSWE1Zca8j4gl2OgAHtu2Dc4uShhQ7T4Pql07NlmpWGN0rbZJkUltSiuRY
sksERZKUt11NejDcc1k0cgc6VoXSibOAHxiplEC+kxVslhQo3oA6/x0YgpA8kzqUXXvSpRl4nXxE
uijT6jKumA0Bo5NDnEv7f4HH1BDPdfSbSW/licc70Mx4vZ9gsnvcI71ZqXQw+taDuzH729bo99Dv
/QTw3as5AMEO/GW/+GZd+BFeqC4KvlTjBDzgYo6rxeYqQaFqDVOuUsJG9FsO/m72cbTO90sf8U31
6Zk5UHvc8b9DNIDG90lSLE3yhWhtHU31vNtPD+G/IrGToKsxwTHTNqHxyZYrVT/kxF+wmM527tR7
5mrfxK9dFnJou/6rY+8SPcw43RNYjNMDQSKQDgQvLe58sCR6lDv1HDo4EWvPzyn21FGyn2C+1D4c
yE5B9PLmRXvqA3728Gp18Uh1VqHdp0LGSsEKlffyd0pjaYYRKMHxhzei+57eED9TqmoQXG53I1vb
GPo6wCx20exlRVUTVPhKOANeRQGVr/8F+YlCpe1To8LvZVzRb1xSfQbaO88qxn47ePPT02nCab+i
Fb+C2W6bA68bl+Vhv+pPKBQc4D3Hjsfp7C3U2Ehi+P7MFUaxbOFpsNYfMywxwppXYW2enwOhrZjr
RhQB7Iz3ESxy0zzjoF2Y8XHsUSo8wdfndhYWJRxWuFsHYnbKmodg7z4Z8pkkloOA/PuZftIsUD5H
n71gdcAOGkMtXPc4Lm6rbjS91bDg4r7s0DvGJzDLxCtKqWxxrE7nv/8N3atCdd6HPjHXfw8mHY6d
NlFwLH5Ed+mlcRU4PH8kXckqR/lUJLV12TyyzW0d4gyC1HNbCGqkqWzjlK4+rcW3wVRjSci/IMot
UaMgI/BfFag+F7TJAl1LEzeYrhSyt+AbzwJDfIIRJaPPFE2iNJqqdGWA8260FMQRxl1fex1vwgOo
tdlEhnPt5HN4JXLy5N2Ktwz407XQPOFNQsk3BmgjLSknos/PrEyxDg0ozz+9V1qKpZZ1bry0fXC5
nzvWdpvhdXVPR6CRP2bjqTtMhzVY4JDSp0VhCSlzDT4pnVaqFyjUl/D8e5LnJCGsvBOWMAAZN5SB
tz3AsdPuYuVNd3qeVpusmegz2Pz3+Rr3pqQcrahAf2BRFHrdt7P0mSDdz0cCghcL1nDYcKDp/vvW
GFVapV394AzYI41GTR+crw/x+i1hiRuCf1BiXkS+2GzMFMgaZvtH48qzZF+V7O0qE8ZBsxRolZl5
QCq2tkLnXcUM+2XmQ1hUYG6+28RIOWOqub178t3pKmrZLcxHGMxOtd9K9jMdDpH94gKvLFKEMa2D
IKpQBn//9VB+NGnxyKzL2OaR5x5ijR3tsB/U9YzjDFpXQTJNczdr7H15CnjO74dn1SaN8q9z/dfR
U43d4IEV9rb4RlXha2aXyGzKgSmwbkVfJ7UdA6BAfCVuBFanGxwYjf0wKfjiR59TUuUH8tyBqCMu
u+VBt6VRv3UHBsfyZYsbdPFY6mjsqG+nEa0XxqEEEBD5MWCO1rl5xCnTPdbgrOlDJVsIca1q9Ie1
nN+RAJE2y+FQ5/bTNSZ2Ttkn3/cJsqyPtmLTNdM/LM4OupazIww/eg3FXFBLpLV6mJ/DYMsS1LwV
7h+sZaPs/g2xiluNKhKP9yfT1go0HD56M7BRSbx0vJ6T05LhMTkKfz9QUfErDIO5w23x+ms28PaR
n976u3diGHH/I4S/As8XLtBvyCCN2sxrytPhqysBzKo3IMv2mCzkOlxHhmg9kuqlP0veAvzl/JNK
E73reiEA+VSOaFcr//fQah0tnHQBJACHO4+Pt/KA0zI6aC1x/xrvgJ9O9sbHALPQRieWgY9jNZhI
MYF35u+9DvSZx+ec+D4UsM1njYp9VMuHGlNnDS/VPTUryKWCRGdYwzRbjaX84lAA17OFc9OUC3my
aJIFIZ8Py2DZultm0KhE44ZHZQ9XnHJQrZIrCUh8oAkt8at2ak4VwF5vO3rrNr8epX9QLc/IMWVN
gA7qsB6QPwTyzNSqYc1E7pFPHUsW7eSKE+gslxsDc6NsTHeAbW53tC2Bdmpvkx2nBGzfkaeytDGU
KpbQ2RxofWQirxm9/dCHR3ILbK7aIYFCLrxt8TfXD9BpS5MslXpAYO2DQGr0DVY8uQCjiQ/Excnc
pB2RjENpVcvB8mpAX4kCxcYUAvUgoqwtxfc3qjLD0y7feqqz6pe5Ts9NB641mmXyGKVCJw+kImGf
I8eOjovA+/pmaPDNTRHI/i2hy0TxnO4sDL3TwuGH91G747nYKTZgHViRp+chPd2pQT3eXEYzUy7n
9xtJvFcek0YkEXtnSO+McIUHATyYkQHolUSzYViNJo2LNRqOvIwJn1HMKhV8wo9C8JnDfNB67uy9
z/c3zpVYvIz7xa8QMCzlKtt/ntyBgsjWoSBnNC5buDgQztZieq2GET1Oay0FfdcfQvk5E/orUBEu
9NOv4FpRCFsnjMr7a7vaVpsvvN3VGXROfh5Uk7pCuP3HFoo8lNStZYbH33todzr0zSYymFZEDoMx
PWHisDULysp1WaclDMsTedjbJo8OFvEl0SZBe2vQ3MKiktGv4GThbSn93OfM13So+1dhaiw+fMdW
xThGdDRGmojaNjIHCKQPr8HpLMrhRArbxFqLgNgkLpLxqNpAIdaGL/Ztai9kOKyYxBjEKnx88FmR
Z/lVd1uBn3iAgmxjVgUYi90OoL7eUSqyh2ehWVRKuOSbS1Hxcz2JbZF9HtKNv6n3uQ2kPqZ5Ojom
BMrQMCWozqA2CjcfsH7IrxbGLakbR3QSONlbAr94Msmr2+xUPp+fjgOm95H1KWc4aVIxB1N4QdVU
/uvELMP/1TtcQE4D0yYykJT9BiWictHHfcVBi4VbakMGKGRPcKeFCEblov95c60P1IBo7VvLokBY
al18oVDNoqkFu/q+Tls5eqUwMTAkoqMQHMARIlN9k4wN8+b9iY0gXzO7Ylegh/lAUA27fryV5aaa
O5H+QeTc6Ca7XUZGAQpR4qktcBmC6bpCG8ZUI8j+4Qj/Nu0Wt8rvOsgu9VESbXo/kFZ3BJQGgR55
kp7n5LU3PgCHhhDsr5PwlPDwYLyR5crAplJIldQowXnwI0comnzeNz4rK8Z/CcMAdOoq5dLwNsj8
l6icKJgGp9hDNZOOSXHXWKZj9nI9jix7h4D/upoLnRiWchqgla3hdcInQqv/DXp2+W/8cRfvpuuF
wF6EJTFVDqQrxH115MltQJKSq56SUkPffsCiOimBdQOQT2DXpJOZsF2jXIIW6MYaWZJhKsoHNB9v
me2HiGi4Sm/S0cZ1tdc5KY4VT/K6SUDxamm+XWb8FDdXbc9moYY/cH8dH+YblyLuAihiujwP89Vz
pdnTSea8fO9pTrr0PYCi0ugj+egQFHh+DD7rhpD4bVECd0sHSLKHlADDTuTcrrKtlGBW+uD/cAFP
h+/vFsHBX2uOwBGH/TkdBouFe2LaHycNV4BPbK3fWHPhZinckm4rByhLkOhUAb27WVEDiA6dIceY
wfv6QeBR7Bi2awrScYuEmoJTK1F5XBi92tOH3y7K0dizt1Zal/Rl6n5UJcYvvSbHu58cWv5FWwvT
SsH8CGShEzjycmDY/ROdnE4s3UFV+YTI1N+8ZbH5RprN1ktP/Uz9DmWZfq1FRRDLNruQObaG2fUE
qxMYX1AoCrfc0ZfGbSNeKeDHR8/vlqqxsUJkexIQRff5kK3kKOskrsD4SKXGrqViXFwbspC+GfAH
wNt8UAqMIsVHN65zwP1AuTJ69wiUE5lsxIICQgAN251E6YWq9B+B31iREaBG0zMDEv8aiCvj5knU
cJ1XO3TurUqkrCZ99Tc8rl+8HcWXz+5LMPleupN/5C6pLLcBtOUitQA2NQl+kG62lw59uGRc+MKw
+WFRiHBsXgwg/sS2ATow/6H4wvCzKzdG6NCz85s9ovt6s9b0RssepLLnrFvSpDI4I5EjbFvrmhRD
dGRn14KsSWJ7ZbzoY53fxJwcPplQsjhXvIXp6T1xIyQlm/C2UUZxryfnIzE68KQmowsf3HSTMiyv
h4lDZT36ZutWchVgTsybBdWny2xjEkIgkxgqCwV1UpX40QzAbv10arcXjnYBSKLP4A1CJpZOuVXE
YGg8vdSuyNXNHHp4P2Llk3Ld6PsHVh5btbtHh2PnEFPL3WTxyRhVR4hDyoK2Q9RWJ46ZYN20G6bN
T/yFUtbD5oUFL0I6tFnzo4rD3nreqgp0heXvXucU57MVhR97PtS92Aw4MZoNpIUqAtL4Phmw4H5/
Pz+6E9RfAkg5EOL0vdfzEn+dX/A6p4AHSXiQbDAkzXt/fuZlnci2Cy8uwVcWT3c9at5Tvk9H7jVC
7+i5gCaV2hjksSOS12JPvaJGOPkse3V22JJsWLhQHP1AVwrjHXVBcw6Cx+PT67a+WvUbV6a4uNE7
LN1jqdqDyp02mVGmmh0Hs1Y30/nqCvrS9N653Yzl4UD4tFS1KXIAex/X5GAMh+ZOb4LJM5v+wbeV
DYtSsbbsRQkdpD8uHUCTGFhwM0TPZtr3GHEOUPL/0HJzAliQ6YD3JpMClyrrrGcpFKLSws2MqJDi
pA4/UAr6a7r15DAscY/gpN9x7j4jLHC6K0Rd3Y0zM/Lu+SjwUZPmQMroKlDnql652Q0NdvvFkRWm
Vnyi+unOeKs9l4sAgOAJ8hpHovBOMEYk+BklB99IO0BMmuhOni1ubWV5KahSReIjIEtw3jx/1NyP
1JGgKwY6MkfdSZ2SHBDIXTsahSf9uNA/yGheg99FcLV9mJ53qbloHQqkwuBxcMd1t8hJAf3ziUbh
VwWR3ctcpO1DJKc6fwQpCyacJ1LiaErcPfZn3K2yNHMVlEgNeXnDMqAw6l/7ObdROgE+AXPq96dC
xX9e8+vJSPLn5Jf+KCUMzOtS4TrVbxPXTH47wPLBBTR/Jgmr4NXlM8xHTJpIt9JYiLsXt5ZyCHG9
hu3r5D6Q3qNdbMKE3pvgm06tWCEpD6PlM++G9DAskstKz+hcOU2I8zrwNF63E46VWVcOZ3278nOv
IG/puli2yL4RTeIKVC9tcTS1HfAfFW+zjeskfn7sP1mEQyDwJHEV/2B28VzkbiQUr+Eb+/Hh1w7t
kByRt/YsSt55IrIJMlcMo9R9FPORric7qnduOZE1L/kBktBTedMdALsu9NKWVsyDOfyh/keWtAPH
QnEif1k8SDRTR+qreLPaUInjY5z5cweuKgVB587YsSv/9IrMGZ8QRdG9C/PrScsgDz6xaNbf10b+
t2fDYw4zgY05fp+Tinn9VRLUNYCWbYlOMRs3Zk0YHwtrF+ubGMr/PPpderiqm3jporSDXTaM2kiL
3qXPoyQgsgd/AXi0nH/y2m0a1TeSkLE+NdLXlsdB9f0jmp+GlJYHskyPzV0eJM4LBRXJTBrgud8/
vJM5vluKmItVHL+RHmljnf1Tt0p1E+Ghsy4ss/jSiMuVKz1eLfCXxTU0Pri60LvvM6ePeaf5rs4L
UqU9YIq4LzjXLu3p2NPqFKeGYbZlO5V9xcyHr/OSKNTYCnlKCDfaWJoKkEHsQotwhq16o9PtmR8x
rH5sjqs8FXxgvO/w8xp+XzlPF3MUO4qcJUunosElOmvrdA4qxkVj2IgHHGJj0z7+MBRhdVhCOhwV
BknuAyfcxug9F/kb+gfa73xBxx12QLbqabM++aDcXlkUC1whUDlVAxDEPmJzR5Xf5eoIgeep9QCB
kjNInkrtmgOEwzOlWhVZMUyd01gZcmIUhD51OJvrfbmsjRSiAp9pRde4xiHjfrYCaK2RvHUdSyNn
5mArwZEnZ06O0YGq/7IHQ+Q4P7QYT009zwm8m9YOm3x0DlNxRjnfZYq2ZNZ6wFHLjWtYm3lT6IaF
Y8lgzUBPlezrOLXiIdKDxEyNhe+wBaD0YpxNrPt2/EOjviLt/quHns06Xsz5OlPDBEyKVMMVS75m
lcCsvRuBsFoiRCQ1So8FGefRIAona3OTAwKZVWv2RQ56vvYOzveMmRo1TCKl3G0UMvqA0WI9wy8L
EN+Mnw3FuC5j0FbLOCO8hJVkX9rSAixPH7ZKpPL2Uuc5TwRj412EA11k7VR0FBeSqaqTOe4KTzqE
XF6jpFfGk32pntc0v5ADpm91n5IH/DOhBrOxBnxFVRFIWYFEUj4YttQw5wqgLN9ZP7Em9XZZ0nBJ
jgQhaDPGt1aZHChxkTzL749v2lE8xGk4NiUC+l1QMEJNe/960lhwdqD4cKanhx9RbT02efz92PZj
4A5zkXsVICu4hJHbedd0048pkZpLOpFdgoLZDEZEoak9B/RdlfU5Akugv9k1bf6X0Dd2ssoo0Kqb
pfjhFClIsn5iTjm3dRcrPkfKQ/n/UtXeM6FGduYwZMPHvFwfaGRJmygtgCkA7Y/CeLtqLHlQc+nR
ZHtuFBLFxYguE0qjsBV2q+CQ32KbBl5ddVtZUFHgbNn1ND4BtSLLwt+kjToErNcKpxFdf78Ll1EE
IgdRRj4Tp8lzzSIJ1mMQWeM5m/B5Ve+95m9p7Q9A15FRmm92kD/an74A46F+jrzPDYjNL/M17SWa
lBCg50EAk2QbaZ/ugGZsO+vOIqwmJ0VrysJbbvNHLINJknEzTxLOk48TG2WNn4x8jDwWJ+kJH7mu
5DRCRdqKGbELJtqlwtfcm545KWyD3d6eVIGYN882FWvTrDWVsd4gXZomUJvLGUqZDFhVpT/F+h6T
bIXCUczC9pL3Ijmlo/cetCNmwABfCECCZ7lHCJeVv4Q49jXPf2lNo7Co3Sl+tJ8sKjcZ6RntsEU0
6BwIsvSI1EdiBs/zPjqgHmqjMgQ4RjYW07krO6+Cw2mSVghmMwwI3LFJ4PWEKJwWkXBBCUncd9NO
dCCBWDTek1+72cr4UyB0AbBeVpPOYaDVtS9M6lErhkeQRHl0tRv/5RflGDs900XVYfKEerNpYvsE
rhwgDLp/qeq77uG9jwMRlG9v0X7bxrBNBKo7JJRQX/0CHKMbChtkEDgKJuZZ3QNxP3P0tMTh0x0J
Me8Dr02eHxI6dpemD4sT9kfBYQash4LXnuqAJyONE3RaEYB1Z17+K8vR6Mn8IbLMknjSOjLacVQk
Ds9W9bt1/eCRktCyc2rZaV0X7HbM9JThdpMKeLxJCHPERmuPdgXGvYnpKQVqu+PFGusRWtGg4G1R
Cc4B/t/9lPwRPbRn9P+wr3OIuRmaLKuASGUVZtb7mGeSBMrNZZFAKCPhGvX7pxneOn04gVi8zOuB
aWlyIxkFVKuFC3ygvEJAe/aXOMx+CS5/p7xrZGl11KfLvycc6h+t/Ww1N0mndmae5rfNpf0aNDzv
ELpn1V5IY4qg9j7qvUWYL7JG2EcLC4h1rJYfzJJwQozkQofjAr4fWHPEl/3AkeNKJ4Jeh9GTIKqg
inhVyZ+/DIblQC2/n6awzb+sFG6Xz3vjNyWFjNNSNSgYsDFPXpBetKceb2A0Vc9NPTeCYG6IrWbz
n+wXApajA7ZLEafgH+bLTzwqmvvpMFVeIGm/lT9DNh9xQQ6d3bmJDPyJukVHLjZIPzlzD8CwERou
eS8AUiQ2qPzUxODbLpsWUdnY56mopc6dDzhUb2L7E0zcBpSkiqQCgRWzeeJt7OqONT9RS0E30w+W
CvdifjJheWJmWsczovtdO4k82VeQ6ehl74JlaDF3TvXjeBKFYGyIvo0SVKHzDisqtfiXqGsWDNvR
mP+L0orXbnZIo7TBYxEsiCMfmGZCQEoj9eBKnCcwFsVx5tbUeecEaOq3sVkXxVCfXBYzS58Qx6lC
QeQvQJESyXSr4BBHPImQ4X2jcVCvkF6W/SI9wgaeMmOoIsFv60iDU2ULYSviP9spfe23SFRu8S+w
es6AV0qsPgbaCpq76LLAalXs9GRXNfDabfZIIkZ5K0bs0yYcI+wq+9RA6cQ8ppRT06xtci26H1ej
D0OGvv60hi+LF6K5IMf95yOWMnKoVCKaxhAEelB/LaL4wCheTfBU51QX8hym08jpcpslQwb4qtJt
abF0tABMI2cYqxEDxDEO4kknsFgNRDhAM7hZmccNa2eXz2eXdQneELRt+qwx0AtjadKi7mukuNQ/
OMgHaLVfdXPE5zM+dtMe6ATT7XfQCnAwcAmI7wr87AOqXsACYWSNbkQY4fo0MGVb+Duqxnv7jAad
xmP7JIbrwiYkosdyjWmMeQ6NbasJfQBR4QSDQFcCYROc7xCFeBxa6xSAkNiSUfpi1bRByudkhyPI
u9GZYQxtJv1aLL908SwejG/9fZieQG0z0guLK/LhSXU0AdUpKh4df0862w67PTrNE+64RM/RyyBr
1quvW1Ks346NgMEel2xRv6EfPERBpt5SmSzDe+iBikMKz+6Fax+1LlsL/bS08K/W6pDFf98lcVdy
4Hh03O5E3LjSZIh+jmVuxHx1aCLx1MwgkCCF1iQ4r0LuDBWEYkJTO5MjTX4+QzflGKfSqEb6ALh+
x2Yv8XVEGNqm8qcTgcveVkLkvZfSOefoWd32jQYyjpp1+4ant8eubwsm1fomSQhkE0Q59EXwMwc7
gsZn275fM7/hB41/2LJR6Cqmy8c2jrS7doh98vnEZYBqqoI9hNe6l6LUjGB8NPJpu3YMPtm3Zqtx
LYWbEBHOSF7yM+oGNjUJlI/AZjCSS6qxZxGKzQIlNBnNpD2DSrDBTehzzCp7W4XQXvbqmPaqenjV
7Z7XcXwP04Z3n1LH4MBvtuZn2Bma5iUPyuxFwn7nP9G0oma8IkVE+U/+37dqnXOLWaGHiYtZIDMN
ifq1Kq7tWysJS6ZHV8QujGqzw0vv6m1PXbpRH2tsIFpmDX9QXNbFV0tKoG2CSKa1+QT+EEwaCoIS
DCHHIPuZL3PYivFBcDAYLLJbpQUFSBITHFVRAXVjFRevHLhdZ3zAbCIb8UIv2ZfmuNNw/1vokZai
AQLbjsaTvW9aXE0olRj20Ynh1Vy+Pz5ohA0goXWZB1grQw839LzaOJ6sTRyj63G8l15dit8UMNZc
BTr4l6GDmJWoXvvjOOCnetv8//ywGFW0A+zAGGEZu8CVumkdzFqjAj0D6HR+k8pYYZqcSEDyvKSa
ALRLauO4ZuGWVZQMUGJg9GKaAY8RoSHVfvHnGUBktia8IXZduAh2HVyaNoHthZfEif9xjAPukp9a
j2zhP+G6J9l9oMb5Fo6pI6F8fuNWNpCs6L7P76n5txol38W7UmwnBnsGEqzOjcXuuDU3T1XqH4H3
CLZ4fawkTogeCngx+dQWlbqmHp56zVYbjFY8duMWLIajMGwvCIAYe5eftctPKSjcnG9bZCSNyabq
X1qE6zncLBRJmEfJz9cRYorvr7Y3513VdyXfFAPRfaVVd/Nkc7Vf/QzO/pQ06vdHpcje9k+dkfky
zhu0quei+SkJR1Z7n7XfN41buLBnY/ULjUMnrgFv6Pu1FXvsJECXL635IkqvFYVMeXtUg8lAB8wj
d0hq1kPWp7SWdDKMVysaDcQ3NVGHywwaqjS0Mb5FEqgp8Jh02ciSv34W2JYw5O1EUddM0sMYjNOB
ctHFTj6u900BNBzLiOzUdkKZ4cRQUWx401yzHiu9MC6GY5mTA4Gu6dKe7qCT1qrrcyM70ryYxRQ7
dyPuVfhR/kQ+Q9hWSac9BX+3qPHUI3oloHgEbSOt9sYAK47/B6hZhveqSjk1TCk8CTgHtWh1Hsff
47YDrOgTGkDYuRAbYAGkagzjxoWoHVqO9GqoHgWWsbHtKjtMdSxBAsRiTsaUpiGXxdWitYhmatfs
BnQxcROWpeg4TPfuR2l2XUDXR0PmmkUoIP6TAHXZ/0YQU0EfqkwwfsFoq6TBu4BhXqDRTvflJ0XL
oTj4SBDAiXV7njsx/n6n35CsGjLIQGBC27o9mtS0xr7vxU7+QefHe2XJpyeuwd1/08bfDH1n+dIt
TzUibtWjpr2mwbJJpUqnETIPxoophzkoNaMY5LN4RwE1WHIMc+BwI3ki0FMFe0B9SeH3DR47BphH
DoTzphIxgIW0xM5Dbseq9S4jsHqAUnRb0mahNPxUKDBvJYjBtJcAYibti/K8VGnFJ4v23+EzPXny
eD+CqvwXiWWnpApIgrXeAIqg9GGy2IGdxVAsScJ5hnMfIlqiPk3NFcAXQcTEFEbJnRWAlJspbCW2
otCWtHk8I+KJqYRqEPZbMYSWU+9vNBEJy01lo+hmkWob3Y2AqxhP6+UV6t6MNXnwXTg1UJTGhamX
kDygO40D/mIyRunMjrTzqOcx5ZBIsdtRASYoV1GNhiKaHzVUsKn+FnFrFvJUNKWalHgt9Ixq/k83
XARmEYhETIFDb1qoHhGbJ6L83ztzgCsPDF3gRr8DhnsclG5hRxA43eqdtf04Gj2810IfTckR9cos
kNZplohpWhE+1ZNLlLACbe20vPtqKpZB2KNWU1ew/yPvTIaAspO+1hXOCTjwGv9LIBcTjAZoVrI+
B02WpQ3q3Dlq2pDYs6ytcicuKhQnE36/cfl3XO/A1f3BOwT2TPmeiiJ2IbYhdbdrXZJGWdpXXI1/
67jW90hAxyH3IMoJWvw3Cpy16R+rMhKzFNQZQAs5Rv4Yiz4JSNz3RNwScBMve8fiQnSHVFBohdPt
Y7cVG50m/6b9CA4qPqU8DpVagKkKLIN2MVuod1dPic7rhtpQHRUiSLZhMvmHtUrHVGa1xL+jebB7
wrp1Yy3EsrDc8kAmWAqgBQvnAuynbJnE/n61uawx7FNUEi+ZDu3A7hQrhemKHrGu/Yzdkugu9ixZ
XEEU3BH4abBphngFsnLdtDYDFeBfcADmO9DqcJ81MMHBY3p5gkYS8nSVwv686IoIpxq/PPzzxxM3
p9z4BnPg6OiQCG3e9of2JiwGFA3I9AbYxUro/YygD2DAQEp/yl0Wlma2w1S9XwW0KdOu4r8An1mG
b/bot8ROEzckIoVuRBPOT3NvMpUWvfWGln8TiiSq7pcFNCU/houwu178AHGNwteEiaA1iJFQL7CH
ASrjQe2V1bGdBrS3F0WQg7hJGX+WImZfI14Xq1yqOaZAd0fn7drLEybiktLUBRL7IYNxZctw4dgf
CN6H5DRr7NnvrV4QTb+WOobt4AZgeCLvLnrvAPFH+VbPzJhXQc2nCCxF/9Liytehzi0AfQvs3wNA
C/PmOUO0SprpHCRNaXLkYDvlXHvF8EaJItNyd+vfRY42Mi1vMfGym6pHriKi1Coa9KxSQJ3I3ISM
pe0HqOVAxKNOBzrj8Ki1Hvly6dV73Loj5NATJABsvhmA99KKQCj+K/TOiL5/55EtYrf44G8QsNF4
X9tA4JJ+59jB6ok+MG+O3JKmg/7hUuirz9XFnTJUsZBuHhK6od5myZIq6RTb8vXqcJSNRKP10vkA
J3l0F2j3MYNBbx1acqONOxpnISASbg53znyDVCOoOyIRtKihtSu+cbTphdgDMfVEvC3HXpe6mPeV
FNQ9AG0ZriT41/yz0gW+6VmZXyPmy9Q2xrPIF3QysXyq76S+gJSwDkl7KH5fpn7phAGmTubWCvGa
lCnr4iomimhvQ4PC/ER+Qai5waw76bzlUPn5QAT4tc8n3MUR51RJo46GrYxKtl0TissdTC9q3RWL
k9+Sz/1QRVqTYsQJCfrPnUK3W4GLGwXZ1m12HVGp+hCRm2pCCwwLNnXi3398OSnehusmCOs6rMBA
sn/01QJu0Ev3Hl24escAXJcYYcgWa59KtH17aQLpzZniGucQgeL70ZAvSFHnl4POHsGKn6IQ3iky
oTNLstfpib2b2y7Mh80sx3ukdO8T9Xjty7nxTBdP+wOOrsQAeorPc0kVO2fj4PDOMX/zHNb3sZ9P
53lg6SqGWCajUSGVBvUCrz0M/fC0j6IXZYtzu8S54Pm88/fCq+W+/MwcxeKyYw9zpIsTg2a9+4vj
FvjV53cf7XGYaRlGCw0BK4IQDXqsdeL6PwPhkFHvS0YNONISkzjG7wYG19yku9XfztvVFpvc3cxQ
P+/0dt2pYt5nAkzj+uL/mFFU39OhI6zhgLZ4CK/4Q8Zct5OtHGCJptn3bhPoE9xaBqVQZkbBlloj
wLxy6sflVRfZshqxp9A5N9fGFQd2N2hd3jO2E30bbWoNPe72tZ2pJRwyPxglXHFB+X1tW/rvTiEW
icvAUHnILUZC7SJz25/K8pePBEO+I4X5Xkx6DyowZRvM7Fnp8H/jQFfOwEhi2+br9KZC0uasGUd8
u98egP5UPHvxCzZgKa7usxXTw87JPgSbM228cF20VjnqZIeLessbUtZFSW4UzgFCD2hh80VPsB3f
v8jLSzz95WBtqdk4u/S2ej/XRQqXYdpHBYuYCzrN+0ZijSqKLYzz/YkwY+D7vfJJAq6ZMUJXaWDF
hPO91MqRuqZpJCx0xRAkkN0TegHDgkkkeUCTiTIi3vyVqrD2AHwXhFdNDrlMZG1UAATEvGZ23hup
nkDfJ5uouRFQ+0fr9keKxfBO2SpAuKJW3LSg87iNJ1RWKHxnyZFbFL6p/PVL6x18GOMN7dQ1AV34
yB7dAiKGJPeB45OyozeWDBd90DVdl3h9hW9ZxO2iWqeeyETsjB5p54LoRHp2gwJaz882pATOlqB7
dSqBsCZGpileccWaOXzANAL4xp9YO4iSCWERohPwmMjGxiFMjjQ24UMAhW1s0RqbC6zSGYuGmET8
pU+w3IwVhNjEhDEIkl/VTWjWS6nGdj17nVuO0iTVMD4YaIW8AvXKZWAEJDhjoM6437dyinu2NK+n
UrTVNjxQmzuHvuG7wuPaojgBs2v+thHbgpagjHU9dAQYFNw/49EnnmxofU2KlQ6BdvZASDNoG/hv
eGXlcy0qjivPOJsFuKWolOJoVodPeR1qWDDOssJ4eu4+XN/F2yNj0FOQ/x/q1Pmzl28cspns8N1Y
bw9YGjL3vJEoEC/8WdicuFGShcmpN8mr8OLaDyonPZLQbqBamxJEhYrcROyO8elYXoJygoAbDueX
dgqe4uS2yF45prtgMYyg1/U6p1qzofI3rEaOqtyP4EyDhb+vaQHI1iUwtZoStZtbyoryGg/ARDmi
aQBo1zPCgpEPe356JCSsXRbs/oEQ9o0S2O8XZa7ivBCsjmc5RkFghfvt5LJ9MNxtHB1eQ7R0Cv3z
/0vB3tV+ZhAXFlHwLHBckUR7W5X+udxLZpChfbk2bbeaP9oj8OPeqpQuf4ozmjlLce2o/cTgzkjD
UHjb3dSj4T/xdoUz4CMXkkn3cl7TxjBoq1XfllASTZw/KcRUgMC1JJvvH6maHfHdtDpn/u0MbLhG
QZ3sCwqBYB8tN50OaZXo42HW/Q18hjV/p6tnYHkqF6kn8e61fEA6Mx7rsT/XShcl6OatvWIbg8Tv
L2/2jZpQgqAyG25v09CWh+b7dEbukamRzCS11oW2TEsfL2v9KpML1ulv8l1+IOiKnvkGLFuAFRXH
2Iv8OvAWsNztznLgb02mcx9PIEu4wgvPg4c7n4qzMkAHYpgfVHHsy6gsaWnz3Jk7s+j6FW8jTluO
IkWu+vIp8kTSKP2juIdb2e82mTFu4CAXhChFOaZ43VwIfvOs2ovH7FeLPFFmEuX6Chl7f7X+MYJJ
HfVyFohtBOrCZrJ0h+KbohopfPJEDnAvo27gALWcfmbIvvMChurxnq5Mh+h2Ivumzu7zbrbGLrho
Zd/zVnsEf4sBaCFRW4SLMRwqfQ3bgIxhbhUxfRoMrkxEL2SsBc0XTx1n9OV2noeSDoDK0Q5fWjXM
kbeOf4gvczipxI1GSu53mlenkOIiKJprCQAqrZEM6z8LYdyqaJMLgy1s5vtfQbQ8NS6IjZwtZfDG
BiAweyqnifyMqTjEqCneSawGRbXmaAyUQ+0MbD6ZYXajZ2wnBNYds9XqcO9b7ttqNlwTR5hcCHRa
Zkmj4GBm9QSHwYfnLUonmQ5GBqUsZKZwXfynwiZB152rf5z2gBOUw6khvAUrG+rHrgTc0/R7nmLa
lVyWios3s1TO7C35DtUxU6C1wDesRdNiATyVr0F50pBW/HyxQqdZpWaGbkU6XC238NaIof+eM6A9
NgtHcdF8QDf3PhB5LfqfGwzL9ZGLyXLcSzhtmY0mIAjUWYHbbNW10mrrBfoX4Qv6nfPVFM22TFEv
PG/UYgHDZdl5YCNegI/QYVgz5jFZKRTCdGqKNiC9XJS1a9pBvvCwkMDAFkbMNQoJ08rVqd51JCWt
CTIDsrlo2ENajUq6/Lsvh+YEg0RXRRC/7Rv2SYqoYMI2aJh1hYxOUfQAngsnfAp8O4D1kFGy/APW
xRguIZy/cfYOD+F9iWe7pqJYTHAkGOXM/pckJ3MaIptNf+Dbg8ZnubCq802JR+qQwfEQASMpg1XD
P5gaTJrRmLAzXdUW2WWqE4dCqXPKWTRI0/YULMG2iqfk8BnrIQaad1nmRoUcnRdPKLlyONRrH33l
ScO4C/ixVkbMalD/edouctkX3edXPRp1PyY5516NzHoobxwCFaG8AG2fn+vSPuc5MTJxS+4Z/Q85
kOO+1QlG7NyUSkOMHCwSk0A8X+hSzfbDFjfyZR0k+U8M+0uQUSCCW5TnDHmGuGXGOjfFB01Lui+V
DZPraIg+IM55xqB7x5aDkmXJU7eqCg6R5rp58lIHGdJTtIMZVav7NON0ThfyQbZT+pmnk8gvkP4m
R3tbAQamKkoq4RxNK6DrzWSX1NWMp0zC7edWtC8FUSgCA0HNibM245xuHc6RbO8k6Nw/3oe1tSTc
HFlSS8ir2QBIbNZK8CMV3CQgTEK9FkWLPxVmMpHznzSFxonTJdGxScVRi3OC8F+zcrUh+V8A1Tex
CsJKjIIY9pSNDfwgM6DkZIDLyhlcx2hHiN6debBq0TjmtBdoCumfICBs7HLZr/QgRv4LpB5zZ3Vq
O2CQ8KJ+nKl/zqx71ev2bxvkioMmkevuPYxytGDYLkTM/Rdy6Ce/M3QtzeCc4XVJ5ZR6uf4apA/H
qfc4tDAG4/qyXFSTkR4LltKpBKMBRPIkjZ4lra22ZBoyreiA1tUGuiM517/ekzYs2IuBbVXMON6z
SXmxcA+75TfPJGhWNa/f/QJUoB4L1x/aQgykrF57yQJGEBomBGDiqeqW6FrHfjlw5Gtl5E/3iyqb
3hNGEckI6deP0oJucU/X/1Hn+AMzqBI8M0aR7Z6bjy+LQHrN5YA1SG5xjTDzMPPR+I6JVKOiNIqy
BeO8OsvCqGKXnipd8zijKgdP5cF5QF64FJKT2J3Wb+52J3yZc7Q4i3v+nvg/IYF2MRebzXJU3ENh
J29YDIyhDi+Bzg3s70IE1/u6Kd4UZRM+uGPhqsdQ9utkIq+bDGX37tuws0IFXnnatA72BQKcuQsH
HF1490f+hAMlpCrOaztPxw5lBzczBE0tRy0Z1Vrxao/kChvpY7L+TzSRLU87/eUb21i3G+4xuhpb
Tap4pShQq1wbI9J9gSdJHo6EAd7XSLud3Y3oFOcbvmE+5Ewm7e16pU+EJlaMG7CQCos6HV/bSPEf
wzCg7I3FCMHJjcTgc6Nt2A1JsxH2TydNGT3RGigF1xMP6/aOhhy23hmJPGuvqqyMTRRs/2/LH8GW
FenlqPBTr8PYK5iW2cjr/9vtKlsFdiEgY6w/m0ymi3X3l1uqjq/rg2pW/X8ZNHfiNjROtPPgdAmM
LM4+1eD1C8w6RehSDny+jb0owXjgKQ1pChpDoLVEUUPmQDLoG4wfCe/pWhOV0bQHZOfRRhYKQxSj
FMlDGnlP9Am2eUtBxkRKetx7Dr+H0auA2vu2ZSXls1Z1+DdymPFdUOTp+liHdUKRID35ftxHVZqY
7Y6pUr9X4aRyGN/Z+wYQPBiIT971veXETpAOZkehLpPThnKuYb9+uVtLn82DHlNnusIhOzfHfOrD
Iczovlh+wfMPmC4eRwJyvT2cOSK6LbIz2vF1b0wXBJMG4URLTAXaFmgm0rmPoG4MWuQWlEKNUYl1
s6H5TtgixcxMzZGbU3C3gDsDn5t42h/7hmnk7/9FRAQh0VXqIOQqhmtFefIywnS/nS64R0eE0TVO
YQ5S2mELa6xu/n4s+caupeab6ydgbgs7JFvljtHQq8dh0j/pYWxcEPpZm7E68vteB2A9t1o6+FZd
7RMOouAmiCSi+v7TiLcaB2f1SHKsoUvUhGooIxZkAq/UC2Vm7UmnvCVjSXIrFSbRd6IR8GOEVdZ2
6BqG85iFXwJrbXGwdejz6ozZOx3cpm98nn2Y7wyV+1S9ZdfFMxa0ktEAT4s0rjtN2VFBoTOFv6c0
SH+7SqZha+6Z3hSOP6I7A3qs6+7FTL2PEqEHO9PBKW2Xjr9y2al6+xurIxmAVKnhR+li+YUDIIvC
ANGRD+gc04Km/ugG9Ta2INg0zZKyNBJvsk81RJ6xv0RyckfXsPpi6Mv9LN3SQbFUtHBibugoHk5s
yLyq/1UtH49X2QJUgXS0wA7thdMkbjdvC4+9krrgFgJjROtoVFNwvygizjON7AYCcDu2S9QbZkGA
ssZhnHWIHmIfJHvJdKW8StXT4IEWmjv2GlDCx8mPfW3xf/zEwYjrQQ2cRv1pvm1bNdY6p+3pC7kO
eLj0ms/URtFAh6FODXQhBA3EokcmCTA7KN0xgf8siUJTLjgIfXOEMyRPomk8UT6NgXHIggj/pWXL
HDrKdB+snaUbRjzW+nNlc1KCcs9LuaJpe4nmBPGZRMSy57yGBcgJcfqAE/zEwQ39BfJYKl2Ib4aS
1/GdmVbifhIw2UivmyT4ClhxqWSP4J/tGyd7ybJ5E4NfgyXAj1jA3VB7X6gFf+B60TA748dh7013
RVSSaJtB8LyG5tqHsmI2irc9/IiBC20ZvQouoH+TS+fVHjU2FeWJuxg4KLUlJy0L6Y+Xli5OZ9sx
F+oyw67SGuvk5T9ZAfsKj+cmKIRUWe+E32KwpPMqtubEuFmGwsKVyx5a4hu4G72C76dWphfW9wsx
D27hXk00sf1TNotyLgpJKal7PjadHicJ4g9fmc8YSWaxnQHrk0ciS4BwgguOn2c1oU+XD3DwwmBV
zyVXKXW2974L1+eTwqtRRKwx+0X+MksGITIu7lf1zmOYdYITlIP5ermCG9nqkVC/uIRd5DZQ+Ie9
fLWpulGdgY3BnnHmHsY3HushG3OLrolh8qzEEjBr6wDqrla/2OJwIAEgSyH07QvY9TRTZk18wrWN
sepJ6OL9oi20QaV/9u2ZdFLq2N8/wkewxKSMr8Fuz6NYOVs2ydo/Oml5XIHzrI781nPzGDPCKmxA
Z1MbpaOEYlkqwgX9INEGYlMc/nBdc5ZPMui9WI1RJ/uW2gO9wybkFctSb5/PKVKTn8ZEYClY5qjY
5x6iCIWekq5Zk2lEg48z4ScAcQjsh7qRAiMz+2J04ESaxkG/C7vIcQJtFVMyinNpBqzyM9+vv7p1
W53UJfQmBkisI5wafbMHXEvfozbnHat7r32xCf5N9CVfFXqNcFiCTDEiYsh+nCUFfZocIfGU3MZw
ouhLg6x2LFX5H4h5dBBcKGVODIUyUA078uksr9bNk/CD8y3VNsPFOSZ25iZwkVLsl+FQLkkDsJas
NXJogYA6VbBoNaIntuvcrEuS5UD3rd421KM++GsysvP5QXkUmpgLm9UEhxF7l6kFDwR7ptf9cN3G
0FGqBDTSGMrmZfWpm+GSZ5XA2ue3e+R4NnPRDQhC7+tuOtL8WNx4/WJejU4nXWNVjg8KkHzaItQL
z8FW7MGi2IC/qaPpNPUk/PR7i6CMLYgwMO6ohOTNavHOspJDCO6n4OeeCweIMaxIK5h6zDN5t81r
LGOe9FQCQ3lo3gno1KctsmwrXKCVtulW1Vzq8+vtPcBt+uClUfrqFTJEo2qNzeHqXSv45knMijm1
c/5RTBexGTzW/ckZ1HTzucm66oC45Gdon3cFHkhQ6S0JQM5OHlFIov04EM0IVcuUqobNypuw4fyL
e3/IWCkB2xrdcNPeJzIGHzO9Kooc1LFNT/bVxpQkUaHVb5ZSej11isqfbj/Dg8DHc/Y51l/jiz6E
4yb5ySFKdNSlXWhsceebG/5iwlWrv0B1IjI9GYA42hESb2szovnK4DJL5uCvMOht8mcLEx1H8rQk
bY0F/YeGiFHl8tGSMj4drd6JgjMUb5gt6cN+6NOd4Jqy+OsUq4crZLykBtkq76frK/czn6m6hGTj
DDfDjUjC6VKa/l4GatDk8IrrBvosqY8FiyP5X9f8wt+3EMihlSc52YlDuhFkUUn/D7a6W0dTm11K
1TUP169MizJ/K5kJNu9CgtlzF9Qbnqo9qHnr5DoUFPkhBamS/l+Wrd5MG0EwXGyDJztE74jg+tdM
nIffr/IzT0JpbU4Z8XLErL5zq2JEu9KiguayvhyBJwuGznfdAF8SvF7P6pBAgMIUCvV9zNeZ/w/4
18RLUX9boGoZiE5jE+5Vt6gOoUt+GJNFZq87Ue5UHN9R5mjqkTRqfC9A/GpjiUOJvegHreqF7FaT
uDbpsrgRmofQMdaUPBuUiZEMQKB7BtTAkh5yxN/F34aR1WsWcPhYfgIRsdicrOL9pzG3y3BQDB7m
pOA9Xz2e4m167vlydukG+eapjIRoZWAEcUeRef0syOSkRl3jg78+MnP6NnnBw4Nqu/eUCefp/H+V
0hzzRJVGMogi+8ZAjoOMpRnTHqoK4hGlb3FfkoD6BWxYHOp2P+5zmmVViPX3X9Uh8f1fXLCO4EcH
AecYL/R3jb7IJqiGFVW4euLPKUYqzg6hpQLds0/dfM7G6CRMuCJZxK0kNrdYK9VJ1jxcxYmkuRsg
rqUFudfl1qgFFZG09qRLJqWV8OQ1G9i5xsODMnG8y85sbS6Udumi3YGG7Gn9K86HCGhqkDUEYbWC
8wjnfya0lrw90wsojh4GCEUCpMQFOwuehe/CHZMgrQW5OSUqnEBsOyMxJFpsIn/VxgywdqMPMkWZ
3k2zNn5BYSda0J24Na0EsPLySYUO496u5pWLzL0UPTZERV5ynPW8zAZuiUCeEypB4DnII0M3euT0
ON0f0pDiv4eBXSPdAYk+Q1wpEWgEMg08/3LXB50UmqiUTH4vvoqbXaOnMQf0p+trHazXlw9rPlGR
Lrh8jA2O/7B8kcQjVfnZJe+i2f2Mil4dTunbnjRaL39xOL4RnJhp0yiQSJdfkoUsFlomEqkemny3
KyUtdrfPQ8pW+UC6Cym489C305fPG8eGVS2hrNAAB/xwcIzlpesvpY54Ky9jeLeHlLQr5KSJo/im
bCrkIfj6spaDq1j15hHczmy12Uow1r0MioyXsUnJ2EoLH3tgmtA/zufj5kTLHDoof6T6tWJTzrHI
santI1WmRiK3EAdGS43ZlC3/trLTjt46uMGWhABJn+20Rlrv7CmwpJ+RIpDqUYjnZxBF/J21bp/9
sM7N89f5XOUObbvAuA5dYnhQB4UWFsPcjf7/xG0XcT+mKqv2Cvx4nnpHkoYuO7uF8COkDUw6tdSZ
ytSAa26gM/A0OR9FEmQxYg9EZYjcmu/8NSAq5461rHp4Wff9mCEr8UazLog5tDlU/VaRU5lE5lLJ
TKI/yqZbDXlxm5H52zD6GwHaqxwO1Iqqdw+kdHLz4QbJVo8tiRAJ9OP4Q0tzMKAkkq06KXbfgbuc
ShE27Zn+d5Nz11n6pN10gyOG6lRZhuOksR/mSK6fUIKWp99eJdugyNq4kskWcfEeGa+0a3iWRdKN
TjzuHsTeKuPdT5SDt2vx7m/dwn4d/2zqQxl9dBgX64LD+Jfns2Dj7IVLmMaa+0I3OQjtj/kHwDsN
lAJtA2od8bMhBUMXzbB3eABMSXqFneDjHbhrpKMiXswhPlsnWMN+vcMOAe0duC6gJFDwmB/6BAHH
c6tJrcoOBRI2Ii0N4yWdtokeEcSwRJDtqaxd5fumVF72S6fvmk68X1euatNTGi9SpFSj2xiOP1ps
ZcYDv7bYahZiu8eePHJRd4b4KzRq3wwi0/7NQIlBvUB5H7uIsvshVmLPLSkzhSx+kdFTDFElB6dW
+fYOd3Nl2s7LE85K+bjl/i0TPVt+4/9CG3rmM6mGqt+LZ5OlLSma2MpcfkHigc/Tl3H0C4CnwFYH
dv8DEUr+ewnANWsg8rUco++JzyV3WWq4fMvxoisf4Y38hjwQfwPHBTMJeMn3cXE1gcrfI5Jvocwr
ml+1I3fEpGVtNmrUKCkYslFoVpWkVfS2Y9yX8hHqueQvCQOm+kz4ZeDEac/kzBQaTo4MhzrStr0h
Vj7J51QBTxvrPveX8MS0GMLD33AKSWn1cWeut9LwtgYUyEXBYpSUm/LDyNsb4bGim/76ORL2jyQU
A6O+BVwHxY/W2aeEKDirBhnaVu9VglUc56EW8a9dCsrDvkJbTLQancoBcO6SAfyHT775dblAwK0t
wI/e8rfyNS8CXPreKpg2mqfrTLIxz1Hq4OLCwK3aEjVesxZvLwuQOiA+k2iX7XcA4gwF/8NA8l9d
jfSDwswBBhBaCuvXVq4miD2gLLXpxL++9VH/Qo53eJV7paFp/2v6qAiJU8Wi5S676aQajiJDDpE0
PAFvyT34VejcJKW7lW1kf4SxdIouN8tZxS/VsHcUpJ87V78QeF75J8t1y9nLuuchOnpcWtm+/6xB
+48/KOZZzHO0NhLVupj0B7KHkRNaYw6ukVeeC7fYJLfG43cnrfdwzlNs2De8g7SGNNxceSsmqKqu
A0bN578yuzLu9C7aOZqCOM0t0YR/+QqCN4yxhahxvoza6QrVzzWaafQcD5g0dARwK/Ultrc71D3k
N9Ef9TAnZhieoVgq2jm7tmAgowmIluZ8OK1YdTvVLhKwaeT8QqqccuR4v8FYhRHhY+I16miM54pD
YPPV4AJIJSgJZN1/+z4R4Hvrcqtl7AdsRd82VSxdFkkLaimOquSc9iZSoKwXYRPxoy10bxW2eJkS
axJO+c+kE0sCjp7fmbTloa8XArKLxl/U111MH4Rcvk4ykVGHZ8QW6FYvl8QiDgfmboYKMNQ1cQD3
hkUE2eXcD5upEaJBbIXCAGn+gdbn+3uiCFB6dtmMWgz3qOfweBNeDiDiYbvEBYHMmN3cH4CWwChB
LYd+e4OySG6KXoMBwHr8GkQjddbh2v/b500ZY0IgbGV5KUaYI58mjgrFeRxaPmn9uu0nDpuN3yin
LbHgnDGKBqDkzdylaGloII+iNBSjGlk0PlOjGwzomUKeKBDsIK5he/2iS5Dr5LdtqvRInQM58PSZ
OXEzQ7B781AmtOBXq6AfP+dZeR/xauev7QJTRci+dz0MbSx6M5qxXlGG3urFQ8HagSiiPviZwXOo
RrxZ0SZA1qJnoyVN7Le3KgcUmfU+KHnDVncYNMX+kTDWiw+sMC4P7ydVMdi/1WV1mZOK0U5Semew
MPC65AI1E3MPR8J1Ayv7QwgdryyAJ3BwrzZtQH4ZWMyd8Muzib6W74aTs+e9SgXXPThnqRD0Fl1Y
8/ayKSvSDCJzL0y6HEgewrOxmq8oLtaxJTU6IxO6mFWeZsM6rDh3gfUsObOZsCyr6cU/SB9K1meU
Xz5WhBB7TNO8S2QnZj+Sgq826wXMXE7z07E5IbTFq/x4rieykEohgIRPdcXQPRQq+tgt2Zb1CGpk
ZPncPgUwC4Wfzrh2PDzKIEf3213PK0o41g2k3KqS/T5y+uEJV/SR50S4Pnss9hpicp7upqaqBvCO
L+exaxmhSGtWW9dUiprQz+ms8Cp4yzTYrnd/k7F86KH9I68zKmzi3VjQ8lBVmkHQ70G6XNvDRxe4
lX5hR1SawOQXnCRm7DVJti7eRU/FJ4SbsmQXQRhoBa1RJJyJVxIZ35pNlmZuaSqcadtZ+6I9xCCO
KXX3+tM0ihp09XdWklSYR274CU7IzyZC/tz0TPkjzE9b48TpxIZRqWDTK2f0evLBGXnKW8FQc8K2
/d1R96chnGj15i7kU9sDfNpQaEVegrhd3g6ISR0/N4MUjoXYaFlcbD2J2AYxfI1aUcIOc61QlWH5
xdpc/1QjeuTO0mEPoMaKgRdSIxbZ49b62siVUctXf8FKTQEcqEg7RuhK7vJ7S5ZCi11CjmSbka8o
xSc9OfnyPksFDWdux/eT253SqWOhsGgJqymXgafFWq2WB9DntND/9hSuCGIzqbMp94LCombT65ZR
gjfkuZwVVotm+vOD+zyvIVjKPVSXL4urzyROlkhsEvOaOtJT7xKY8MElt70Bb5HmZ/tNZK8MvpQO
OflFqMFz31jflcDSIdwdhMoG+zQoxdCpFeb0YtX29A9r0k3E69D+6HHr/cri/gXPAi71Xnl6NRnr
k06J18lqUT9JExTfivTh/OgEKr1/g9f9G8qccubfETYh3dP6t+OWUbOzGfjCXPcA+VKElyeo2IZ9
h+UzlBFulL1rT2JPv7jQkfpJ7Ny8sfycUt98gd7b0nZtCPSMSpFioW7jADLdWv7IdVPfb7GgD2MS
Lxbg+aU15E2+B3OjAKSwKZMrpPEXcNEFi3st51OfmkI9K7JGfIXyXWQqF3tzN6phkrl8RZKm9R6M
wVr/qIuZvwxkVv25jrk0WdHa6GFaebCyJ4okevRxKy7Po3yDv205Hwzu9E0fBUTRBNQ01eZlCQ2V
14HbRm6P94eV+d0Pvh8RP16dZhc1WcqsIW7o8s52PPgL/l/GD6E+FXQ2RJVvgXlYgt+3aH+q55xG
R03bSLomf9p6IfhwQBZwC/yfsPyD1qXVpjlVVjGz6dJFzbBJ1ENvSYxVBAUqjzFcSgACJiIPvuFB
aAYDu2z/L7Bt7P4zG8lwXLKVr0IvTWH74+aljCnp40t1Cn91yKuNkadX3SwC5HX4Vgjsf26I9gtz
QlZ2qTu66IsSJM8iA3XcObdSU9I6F9VgRH/doH3H3vtEPNSBAwo7aUsEoTTIF1Uhfk4i5w9Ld569
zfh0biEjrstOulnU2MeEeACExNqLrCJ6guu/BNOQL/5KvT7y93Yt7EzQaNVKAh2GrtVQH04S/8rx
ltT1fMin1Ga3w0xj1PY7H6J0FPAKfY8H0Kmhw8FLJyo3NgamhKa46IDQWj9ymsXEjeFQmI4qJ5VV
IjMTMJ+HpsW6xCDoy7KtrHP9oLC2yo5ScU3X2fLB04MCKsUp4/9zF4ExkuXlrXei/1HFqSYw/Y1G
VGnNWCNcppLMO660fWRQADeJ5Tc/29KD8wiR3OtNAM+U83ZSln5PqhoXw0CFMVMug/46M3ukYk+k
+FPUOS3gx55OuAEDxtPcx2yGhroB9sMzPowAyuzXU8JZltgjRb5dnMAvIclj1nzykctjjToylJSQ
BczLFXQFhznvCzaWWvf8z+nvUReyGPmU/Czy9GATo+74ENH3v4IIirxtG9nQZIWHBglkhg85tNBx
dqh3bNRG4tnhoEXR6b0gRGv/LRynRf1v6HD4hyvrO5XIQOLoXBYiEGZAQRMEcFVFinGBnsgZ7PGi
YI5JKIDA2UTstoiv//1Do/gKadPxbt621Ug20G6oxHZ1hWrRu+cxnwxpehwpkBn0NZk9BC5WNDB4
ilB79Eu9v3SgK8D+QOBQwhEt6vODRB68x3J+UcDPvHYPuamckYOVeHulr2ki5vw8N1L0NXhx3499
H13kM/fMPP6aItHDDTwBJUC6lKNlxs+KoEPaQlqXthb/68oQalKhX0zJUWlKjqOgwbVcmZMT2JSY
8pwoufrmshjR+jIKJcfqutNJaESCcMB9u+qWpgLxXV7FobnLFR6BJwWuQJS24zIazRQtkd6YGH8e
2f69YC1ZhGEgwA/3zIyCiaZwbKT6BD+854WDTydNyrOKNPOfS6QF9nlbeNksPZ/iz0lCASNuF7r3
aRa2XnJASOrSlFOI+JvBtxDvNWszaowNdqKZ/UfJq9OcIv5Q0RPQGJHQUHouiCGvoTbHlDJQknqY
NU2Xt0mY8YxxebIVWAPWyU69ftUBFwWuoEqtwVIzYYiCTWq6Mqc17sC0BJLfFcC+a+5hL8CIRQEw
rUKAcgyPcK9GGa/yYYADzlVVEJbmDEHn+reMh04ozJlNBmcLWkbjoVyORJ1dxV3Hro9lLV8u9XNx
D1z1xPQgBFd7oAUa5kUIYc1KwXbd9d1JGxBLqdkWIA04gpZ/dUlG6Sv2EuepzfDTto/0j3p2zffy
h7KDIA4Hhzzwd2nNfGIDsntS8wHYzbGthV0F72NwPHS8m2wjqARwSA2ZUq9MCz4OpIaIu7JxncyQ
PtqLEA6PXuXAyRAKYn1NGeqenf1J1WQPVVDHuz1sKnYPmqTUgSjOJDh+iI8oWfmhFnOc5smZRncs
2eb5bREW6RCW+/5jkh47Edfx33aH7nQNrUlDX9bLq9o+e5SfhiyPPbLM+DAagMfpiIoQpv8fNWgb
S+GWvP1mxQbDY7FK4IlCEFL4Os9oYqoWumvZ/wOQe0jQD1ZqknEenQvxsoirdjqnMk+BYLcwG7Dh
fq2SaFYadV/Rwlk/oSZ0OpsfFZyv5uHgHqP92PFJFWyWr/0x2KyzLm8TENEn22OcFBQut3IqphRr
yhvPaYCdzXH5baAeVPeDL3smF/Kt33rx+ooYQGXfRhw41DgLdmceujgfBlBvFUa7CuT8c/B2jprF
kZ08UtFpiOVhTNuufUBmjPxdgb+8A1uMffvcuDjSYpIoAsEEtYVqkbOA9U1gTuyfs4x46EPccoXq
DfS0aCzxFktVDNYDsy0dW5ZiAWRSYUlK/FiN1lpWJ4vsQ1N32/Wdeyjf9BesQigf33hxqDVQBWuU
Zzz30M7O090ogIvoUXZe1UP5Yp9brlCQfmvwW9JCPRUbKyWbarxBe26lOqI/zOOvlDnfnGrrt8y3
m+4ss0Yp6fpPrynUQvydCxdRtcXEgEiWB/Wzwy2WQ0GdiDR99Jo4Pqj8rRwYx+d3Ghrnq4VTZ0mj
WN0PktgHKrTYzU9ibgCmTAqr/M8nh1xD1Lj9nhuDz2qrPfGcG7ppoE4jZZ2kjtXSe7Kvfcqxnnxx
+Ag/CQ0gleVx/9yOIYkt9VJtzWlGenxbtYJI4J/aAkw0QflE9Eb6W/FCAECRY8hktY96T7Sleo80
vbQ76+Ng1ICMTNlFo54Y/53YiW6Cb1og6cTQy+IqokCSAcFcGllzNApzMCffI0AfEwwaO61OwoHY
e5LGB5wHPlNPj4JagNoTwrNSDAD3/oW3rjFispBwSBM1CEAN6nMna+FRTXJq9Sxitv22p06VcYnP
wDxnXx2XviKOARU3IYwKY1mhibmVHLEZAkKXXh3srbEO45jTHRGRfoEkmpUPc4hAhvYRicEUGJ/1
OzlbeOzJod9aOUuFYfgHeMr2xT/rqn25GM80p5nwPhaDq901HW513FTUry84T7MLEzYc296ESySs
mmeir7V2DfsyKj6WWyoxpAJiYH/tAZPhYaQ5K5gP3sIaaIj78YBhnGOxsW6ZypbHn5oFLd2JgqxQ
uwQSpgdG3SVvqD/f0A0gXFtn5Tu5SGQlDucPjWfWb7FF7VBl3mKGt54Ux9kgqHrLzwT39+HUAPeW
R504mShjBCAPUem5C+IxgrGD5bcNZE56EQBHdFEZEt0DA5AFZxUhHpVSzz6y4ToS0oFEHFlnxZ8I
/ba7LYJZFKKL/2vmLQXa14MuiPob5A8AfuFcn951djD93dia0ctc2coG4IojyxII/yknbovOZFn6
HsZNxHu9BV20dcUw4nqcUveRLYjAnrXBv2NQyGJNOoRfZkxZgtLHDNhsiFJB8jUE8ClUQO/u0zlQ
I/V4s/wzpfc0qbgrsNJ8ikOcR2uKdDv7fsJv223DG8b08lyDFC9ItGcMbhHBfGRsbNEP+meW4JS4
U3YsJIY8zFUMlsJCMbZxJw81GqpxeJ/j2dkm1IG7JIe4CnmiV/5B7K7QKm1mpulx8RAicmPVczRJ
OV1O4Vmkd5B+qYGWCM26MElqwG0NfJE6oa7vDhWwkDtxHj2pIxezT5SZoJfLvDkTsT+kcP1beDM9
20GXJbR7tysOZkEzefX4DsYxSeexnTlUEBZQ3an3bA5DwGIgq+7bvUoS3LNbnizp4Nt4EAjjBwaO
FnrOm/eFYoSOIF2zQd24d8vmrXR2LWmHnqL3o/8vWwKVIJ4gQEgYZK9ljAYzOOHBHqp03qrkclhm
G+zu+MuB7nLQWEAcDw+voBYiWaispf19PmPLEppiqZogU5HBBLqJSiR/xKNH4XRpJY8lP09efjme
PsSY2s0+mVyk71qZQILmIBriqU+X9JzXK1N9mVRun71oy97nmD1lg+PLRwnBoQ1vy1Yo5z/bMA+S
JB0Wgjt8TffNV/NBK5FmPknj97is+oP6KKoXFhQ5/QjuXjPRhTKlPa5setyT+RqUOIuoPDO16dqB
B4EqN5fKXIYrmu/pklEdQEEsuVYLkiYaVEzY9hmWIy9nu/FlyxqHUHCkLhXqqbUBVs2/nWd8FK4Y
ESPg6op05V8uy78VBpjXzU60UvDCoAgnTE7VHe83a48HaS+c8EA1hCg0TJWImh11CAhjRxsXsAHh
vwS3+y+Y2iqP+561NoEo73TLSESap1LxGkXLsmBzeyyV/u91mcJxKKQEQS4qUXJ5jRJgpMK26syr
QvDJyQO9uFtc5d/eanQEuevafBdCzfqntCVWuZWkLae+fBR2CYyyFicOxW6Isfyn+w+BERRqFVaH
BDkeD1qQ2dsCUwI8x1P2M/klalOz9IId83GtSvP58R4njPJFv/l7ltzWA93skbl12qdU5jxyIS5v
WGkhcWQzYefDYWILIL8ScoK0JUJf9qEgg2sLJ4U5tLImbIABB11rTJXAqPgnOEbJXuJiF8t0g4MC
mM9w0LyG3Mt9/z4Wawowah5ytCYCjMpi+9ObK+ai4HBNwY1gOjdxv1E5QHInEbon8GeXl1afcWq6
KwdAv4QONKP0j4L8SLfnhpraVSYbXqsOVjsU0PPJnzw4i8pXxARKg38CP9nwBjHndpO0UKFIOf1P
34P280HFb6Th2dkD56bS/Zi8T/+E3zUryUlq4LmdrdXdbkmPOqsXyYLbo4gmTcV1lzmV8aJ7pZi1
i801LH2/GklPfY01efnz04eeZh/rPDoMSFdb7wtMOKg2wSQ94wCN7sPooZlglEUCVVUTG/6udWik
cDH71CKuuNGzO4IhCGmXy9ldQg6U/wzUD2ZRJiDdX81Utn4G1KLa27dRj4LZXUMSmhoRcLJTeNRO
6MxwCig4hbfMmPHXrix4TLqcI07wdDL0fOqXhSt/yTCmBspLdoNJ4kmZVUdu74KyCw96IiP7l21f
RLg8eb5V02ZYE8pGUTzmf7/l2X2CN82+DwqQz16S4Hqa7In6XrBNpSqAoBfdhfMCGUjM3XouLsa1
0A/FVTzD/fem51a9xznP7FFtCgjOae9rA8Jp8OMzKJjPpt+Ed8uqRehlGcNa+zTLAGtT+w2T8oMo
ihawm7nAjUanW2HAtK/EoN2X9zjIY3gm4mteKy58A5x32eDIUOAD9Tv0H7WaVFlr0LpZPVaet7dF
TgsCdkYH6wnvCSXo+DYFFnHe4dSSd1B4A7jW6Zc0aTWbeaZXZHb+GBSg38XOc05Lkmgo5XHSr+UN
Dg0oO4ZDpYvLrbKrxEsG+GMM3dhgLkIB/YoWSd8HQYpJ934Eg71akVvO/6CCm9yPZ0desGhsiBZL
VVOeIyagLy6mO5EFRegTBMDKJJ0rRSTSn8F9WersZ6mlmkDqPrkjbYmkECMUPGtisF8KacLqI2Dc
fsme865kk3ba+/zN8hODyW2IRlPd2XNpAwvWP2usWXsG5MuWRgGrPmRE3ofZ/dPNF6skbU3t3lrl
kfWdUTCz3cuzPw3NFaCMFBdGYw+q8Rv/JEFKgSNL7ZOJyVi3O/uijuZDmcLAPErwgySbeebCuxxg
eKcZOvwonjCVVgAV+Klrm1i9iTiYXijl1srsLAXJwXfx7hjfixKGUoyLm7DeqIeVFUQN95UYo2qJ
RdJpNZsWtPS9+UP/wEcLrj2Y9iwxIHhVqMWTlRB6H7cg76dsiDu7tD9nGAasCPF/yuL8Q14oYIK/
htG53NsBAL5O1r2/Ss4Q0HmYcNJkI0y+13t9apT15k7W5OL9aqbbBjgOl6Vxcw6avTpRpWvC16Lf
gcikuzXW8+p7JFO6Akn5Xba3GhBKmpkba3mkJivOV7jE7Q6mQAyr3iynQqrtlx330x/Grrm9dZII
ZaXX9Eyz7rlsw/wPWrGjBld40dPZOKU5areOpVc1CERot81hnO/yRATzHmrr8TI7zy4ES2fj6EjN
p6/Lt6yNfg99oLGSFlYeBm9GVRTgv6dFv0KpZ279MGsY8W80KKpfdgYjdojerqQon0Kj89MZ95oT
q9Lf7Ty0O56mTdtuje3EfQUcxXkuMPFbCU8yfvfpv701l63888HRoy0i2Wn1OgKtYQKmgOKzzrwf
Wgk9B6Du7NYptouiF86CeC/EtuoKzBg+JMa55VHpC+V7rK4URhhgB0wFOUIzMohUscIiP0PgeOsw
W2Vf0eCiJiQrGZhcJr+Lp2h/ecW2yXaFjDP+2VwFokoDCThYnu5+GpqgNHVY8gYKDNr6zrEhe3/Q
lInqTG/42xJfIrecxlDXMezPbpz2gSznTRPgasxFhtL1gZtY7o2EM7ICb7ZJRwmrM9+ZhRTosU6n
QNjWv7QztXGdn90aYQ3BXBBAW4BZBYMyMnXIO6Pxr3l9Inv4JhLj9qnBHGSX0eFRKSJEhBUHuQlJ
paRTOPePqx0vfw7bJb4YrIbKCOhwhjNA68LSRED8nlpFOQXp18SnFLQPduMoLaQB5ZxZWMjwKrSK
3vytPakWPH8f7ZUl6cODcWmpoS2lchAjNmbit2TgdHhhgb27eIIHj//OQCtRNf5vKUhpKjuOu3Sb
mIMUyuu9N6J6xa5j0ZxZR6aDBQ0jw09jrhDHJiBtwH5XjXK24ECSGkUX4Sl4ChFGV4fldz9Zu0/H
rjNKAma3/2QN8ouwDBatOXk5xtftuDV5SQnkxkK4s7c1of10OlA0pGNMS/80fM+1RjT79IsFPM/e
aun5vSGEZR4exgrhE+rA0nOvwjPuNpWhSEdboJGX0zANwqbnpSYR9RLoT3dtAfTVHX9HixSS7eOQ
6cuaMEdwUaZe50oPYLGtUUnmG4D74+0N9HeIcD0fAjcbv6mglC1ZwkbHah/VL/R3ovhXSZywOQjU
welxILeFoq6kho1WJuHLQTmgbx7uCSHNZbsFQW1gpzAUyp63XAnFsP8FsYYiWtNZ+bYKrD6Kv7lA
UD6K99kq/uAFA5yc3llM6eVvizJ4sX15K/umAqL5XIp/PypFtLhLJt6yjHosnYTfNmzrAw2AXvQu
grlp/OoZic1FeCSriRZn5huGYsK1gR2FzWYIFW/P6krOikvhDaUiHse95+LsGj+s4OT5OfgS3m8Z
bs8btDBCAKcbEJF2LNCk6nGCYhXwWfp9j7SxtX+MUQvOoo/aQL9anndbhF/TZSDZFe9gOYX6NmKe
5ZJI6hwukuieUYB91alqLG5cONctpISlhnvGZXRQQVd2PJFImssvIc6PO0Q93koxGRMlpGQcgAZd
NwjzVJhZCrlsyqRIBRZes8QdMwFVxpJythvwRdeQ4/4yvNkSkz2eD8aBXtNvE/x2mgqyuEag20m1
PWz7d4MO0QojhI/wu6N//C7lOwnNIk/J1iecvJ/sCyYswaiU2yD6XEGN6RuZ7U556kgroZ6MEniu
fuFDLAMDPM7Wpw7RofsvGZHjLY2lZ4ypRM/WaTkORtqOPUgZ5aI5Qdyri4EAIvlRhwdPj8GT1a55
SEfmEcbSgbUR1tNs0Qi4xy81llcCCs4QROch0hAw7wjC4M9BBKDWbg5GL3kApYUoAMjuoPTyrE2D
U3aB4grwauaxb12KlWata0KWCbQ8ee5fEOu0jLCv1nz2txhXE5T1zmCZq1kg+NW1gPR3eqIqHr2t
HE80SRGpBAoKLNBv2Q6R2rpC025wZ+WC/dihsHGlt2PL1DgROOohrKtRwpHKNYhG3wKneFiSzAEs
6OYzmU9MtSb1KsxJhEZc6/sCHRytTmVL7LhvLiKxVPQbcZdDVhvXiae/uNsVUqHa1+CC3k3Lmken
TyONfA8Tzca/FDU6WQko39Qov41JhGK+ikzWtFIuIio7lRPum6Y6ccsNrL0sRrSnuX4vQ2lEQPBT
sOlUMNyw+VevbI2TVT2Y2l1vT2c5K6zMmi/ccwqDBVUtecvxc0sKny5xveVwNH0LrjrvylRiiZL6
8j1DWVF13D9NWm5lUpPNC1+tBSQ57mjwWpsJR57mORNc5yy+RKFtG6BEQFNjab6X4aL0PWP5G5pM
5RsxYshx1Jd5eA+ZPloGD+jlTdhlRhW/lyM4PSD22YbbaOMSEkrXNzZHo5pMfVO4/D9JlW5rvzRx
jLi1X2q6y6PemWr2WacjJe3asic5sjv7M9dPI4dl3aWWLXxqOa+5kBrndHNhSBodyECY9CLxsbzW
ajJZuitWS9CPYnO2VITq0ssPjtAYEnrbG2p4lIxP2x+GEYNhYXQQ5chvAiultMtvR4Ot2j9ezACg
J0+U5g8ABS9kQjYduaDmfEvld3pGdEk3kZlIqxKEl+LueCoewByNI8gSY7KAu0zhVC7qLiBlRc7z
aNNvqa0xvq+bXmA+sD73Sl4TL+zC+8qjTjESwAwhsPzFecs14RNWKAboRb3oYxlnBoJ0vJUZg0jc
jcsl2bfE22wZieTAPzfe0NiN7+99WyuHylKhT5bd4a+S2GqSW+LYaRxUCGP8cdwF5DnnQu0alW8x
FUuDHvzLZWaAoZ6VO8URLWPrUmKve0C20ND3XZU9i8k6TRWmNgENexqfO9eAolrqUaNQynhnLqFW
j8J2qEaoeN3MNCAYEqJynqMVAGsLvA4Bm86fL/icmrZUGTAUblU89ufVon3BXQTeKENE8vjuEyCy
LO5iQFsIW8Nui+EjCT6kQtXhj+WPCHQrjygjMIny1vHfDbSTvr6wS/Z109BpWx+vM78vB27WqtUM
Dmchtxm0wb8pnq/jaGFLu/ypp4DZRuSGsU6FKtfM/cjWlSbNUQNcYIwNvNFlWHCqfRXvgsXa5nbJ
mejpOR2dF1n4k/p9CLdU61x2RR8agCWAqCQWaMjIZdX33h2gtHbqHWRpZfYbtiMc4NzuGEEcE/I4
pxHRHjo09F8JXpatXJOo8/wfTsEzxb7B+QtmfOAex4anaH/RdnvjeuhDn3Q5FmsJ/ro1oqsDzDQC
ZNNi0YepmZTdjPRtdkAVElnYv2uGWpNLHF0wuK/hKFt33JjKV8Ayiaf4fRbMUgKCm3jf3ckw1fQK
d0nf2+KB+a6WKwNPDa7psIbu3y0jsGKidpD09+GzsXudn6rIG+lCOvweuHRZ4npJlgzo75ReYYDP
qu36azmrhmgDkOEqqk8XAl1aPoQYkIS/XsQpry1+pB3RutpdRaXjIhXImUYJVFm/IX/I9ANuGaoa
oAQhMPMbunRlQstpH0tHhLJSjNCJlqPjrL+0mKWe6Idq1/cTenHd6Msp8sBsDTtUrLn0uc484yXt
O0nDN62o+0P08C2qA3oJb7lGdSZtjWUPQTSpny1flkf6C+KrAHwsq+vKnMMOPgfm9qzslJX/Lo8D
2zjKArmGcd9RZhYJYVRB6PlVZ6okAv5dZ07o86nMXM4OEIRTZ7O5kXQe2WVjB2anKeWr1DxwgObl
2QGCSF2cGeWQWxG9htXEB9MMsMSkv/0Wd0MMZXEC0CKHwOBT9vopd1Xew5mLblwFqrFqaPiN9a24
Q39O6Vm50Rq6OueMCon4+JPgIZ7ASEbdZFJndaH5NJqdGW/dDLCtcsgr8Oqcgh7iNut2UiopsZYn
BNi8Z9Pw3tyQSutaPV5oHuljzSTWg/a/EChRU6avFuWImfLhBNcesMuIrvLKByxDyfJRLnoxOCVn
vztDiZPahB8X1Ha3RMWJ+p5gZWk0plG99kxq322ErfrFvaChDq4fcEJDhdVJAy1OSM7VSkX4VtVn
6BjCdRRNI/KCEK/GQEEn2rxnQvlvQWgAZ/OFf14NjqW4ZZI3CmqhsSXUBKUJoyxgXPzAJPYDO9+Z
cedYD0Gh33fal+3YhwFm7kOIcSAq95frJp6UXV7j6Y4DYMDo8skjGGXv28Ozr1lD/3ashkKBcRcL
UZxFOqUF8Ms3cz0JVwQS7/u+9PYR/BtHEDiDWqKZBLahFQr96LMlhXNHNkQPZ4l1FeuLAZUhqkmh
PxLUHdpVt4ZBPFjXSy/Ys711dvU/I1FxOZLg/8pjvcNh6N8HDRw4bey+f8XJY/yPYZNNSQwZPKb+
5xe24XWDRKU1Lf0huPdJCnnCRb4yhB4O7vcwpNXpyv397+gIdPngUs4DK6lAkFMn1AkZiJcUvnwp
eoO2BuWEBgHVkDbcUUU6j1RSD1o3iFwZZTYIoAfXURuTg1k6BE0tLjuyn4BZEHwyh4anhmmPBUTW
shv16yftByHjqjADGHd3EsMyt4QFqj/MszpHpcez83+4UVLCyGHj2vARptHL2E6igtRY85XO7Yi5
VAz6ep8eUbFCUQk/EuJl+lpy4uyOK7x1D5W6aNly/qaZPv/cFmgk5LhH5R6UAg8ykwFKRPFCh0rk
v86PhOWePwJTTwGilkFL0Z3iRGRuG5XYrXevqcCbJ2RAvL3GUpHyjH90XQgOSGfHUMajG9TZpTWn
JZ+ErIYmqJdm3RFNaqvVzh4OcsiIEuLMJYc/e7SkS+0o1ccJ0BYWQ9Tx5XnCUT2OAgNfowD0ymNV
84bap4uHWeVHDfRn2OTggffeFzbJKbEkb+Y1JV2vX9Kqf0MX3weY3nM0ORGt5aneNtoBmphLPkee
8YVb+5wFmGi7gGMm14VrJgZjYML/8W+pTQ8CDQXjAyihnGQAW0kuh0le7ccsyAdhxc7OW9+E6yWQ
xugxT5oPXZeWUWDFVx4IkeRQiA/N37FXtSg1Rpcpb86uQLzUxMA7T8QfdbyesUKJp4v5BVc/11k8
Xd/3sMbH6ybYC53bDTu1kz4vFGjsL1p+ZQqW31nAF2NtTjYfp7uRxhCW/ZOm7eEPO7BTr92naQK1
O7ZL9PLcWkK+axvw0gf2y0575hSaaeBiLwfSN2ax/96tP74y2tgJuNffj8yvIZ1qzErhuuRBCJPU
Ix4nET4kOuEd74qOJWTm2qDOSBFriUrNsyshv9BD3KjdN9xhN6C61H7Bb46mJWMop6dOSOvVNJhX
385u+Lm6NwA2JhSvkJAhv5c64meG7bG/2bhFjna8V9MlaMcQFbwnCSV2/gEkXHkgsrZ1gRDK8V69
0/FngAtAII4v3jkJO2rKCA0SQ9HoXv2SWi5Qr7H6R5lva9DBU2jBZr50eYI1+RqqJpmB0SLxWR2k
FxIiKCbzBFde2wrVTG/9ytMoMznm6b71xYRncLWxSDcLp+bRSEPhdHR1QfId+NVpQzgFgAwsr8c9
NmdHemF++ToVB78fBJRnNw/q5luDM6tv1L1BWq9seywR/es+RJ0vwFfGeC4n7dLv6bcqCDOoszvn
ESyt0nL71upmK6Iyi0c/V/6e1ZxY53gYHUCDF7vv4GZ0X0yGVf6VSWqqM1dGKNJu6YPfjsM+VHgD
GNsD/9oBQKfRTa6bhP5fXADSQU8tHA8uBBVCs9Gpu7YZY5loAkUV24JE8jO9cNL8Ck4SjT85ayqD
dBAgC5XLLxUwqNFwN4rz1EdoViCEVnLzqSJT3Rur2GjqPzXknle2bn57E66o6R/SxdTKLi2ZtnFT
1bcfRASCqRGvz5XfFFtw6iScCjwG+o1pq0mhDgfT9xB6kWHswg9X3YCp1T84i79wCLQ0d6yAp1GC
z+T/HCSy3HtUJOmHXaN1L/jjZ4iuvXqfTfoW6WR0fbfhFv4dsJBaUa9u3k/i3TptoO0Om/9LLaD9
/nnUOzQLoqluPGe7He1ZcPtci5vo7Cmyz1wSU7A3WVefuSuvOQ0u7pQ3mK55ECIPQ+0ZYhCV0Mef
Xo3kvcv7yioGDmmt584lboHJRUQC1x1+H2kQVME/laP8I39gbiE/BxrwJDsg7Ham+wsS6VQyXDFv
MaLE251EFnCrjaneIEJF+8cd00feiBv//pDlkITTxRFLZc5gOdRwsIe7ciK/nWi0XlhOQOORyidw
fS06HJI1hC0rvpAYUNg9z2B2q87hV/ZZwYY079Z8ZZkBal4hcjxqnyGtOtyF+kXE9B0ARtIgzMgL
rzTp9Q98kBdi9id48s7YxS8PEvwhFe0ClbNnzc2+VhmmFXQKR7qSOE9rd8W6rPPFDrC56GemxEfz
k6gcgEvMD1CQXiBeC89wePDFu4ro5aOTd9ksmnpKs+0F9yMqFNqN8JwbSgCsO9lzrjc+VIyZwunc
VE8mOd7YJ7nFcFpNoj4f5mjqyNfIiLZ+wEVh+c4/ZbP8UDlBrvf8GfT6WcGAkfprHW9DkdO7reb9
DDKcD/VsE9Y02MLfkqZB/o9HXAHPGN0vIb85nTFU9w/H+tH+QCC01g0TQ+SPsPT9Hpur3A4FRsfQ
nk/gzMWOWFi7elI8wRu1OUnTb0wBhzc8fnDET0NNyCIhk7kTwsxescmdlZ/VGySPSxK6qSYSUKlh
GGuNdlXcDYXgI5bpY5TTw2bE6Ls90JWTwzJLv700FFzSb7q6lVm6Q+g3HcMqGq7meeKvf9SsH8Ws
qMcXtaaATghcadn/rWh9QC0Y9GJA9hTi9IQxr3RuW1bD1R0x/rZownNZgYdY+uUuxgGqgy5rSj4O
4Wre/44BOnvJ+fQcQj7lL1JVbXlmD0wIA20Kn+7fug9B+eiZ/jp02/r/WxmO0hmhjiJ3VQsOGvFP
xwnxzsIpMnUDL1U18Zp3SaPwW5ZxfWeUTuzVXPfrkEeU00t0Kq8IprNEuPERLaNT7akm1k5CYPRt
xTCj0f4ynT2yWpX0GJY4E7U7ODk7c+4vM4pc74jTuLma+NEM/WawxJfUk2X3hK2oNkGUtX1Q6F2+
nB9R1Ez2b5TtWUsn0GswLJXhZaL1QkOO5I573yA6n1YLC8cLM3o1mmPaOV13yseOy/cEn5cQRsL3
BxGafZN4RGoxIOsSZw1w9bK/2GX2PKvDeg2PO/4sSj68mWagdrQICHumpFcIL2BndCzqkHp/CW9X
W0g3jqcYfEUJXXotFI4ZinKIwzAeaOucvslof2/MpXU+i2APOer3UZJzzMNAB+gKx69ZwCa/6JQG
QX1CcVgISujkj084HuMG+3fI5AuapzbxVhhj4U+INFXUPhL6PzoZPU4fYZEdvUca1WqQBpiOoTKg
j55+sPZp7mhuM4GMi48/90SKzZFX7jWkKl9UHDLvKSrZ0t4gXnc+AEYimyNI1Z6rCqnEiQ1cmTyT
+npEMLaMH/m/4o47831VPLT4jpkegWsqjKVvTrQHaROIFyVtfWBWb4dAGHndqMPsw4wxmwDITWZO
1ZnZcR2tJagAxMIIfPGcA7v5lJT8+l+zMgCeu8LZKNZmV2KMtuQiWbiRHeFmV9+ZmmEru5ar/kCC
w5V3QGuCVEWK74yPcyGeaIxXDu3DUmDimCvrj2NY0HXKzc6BBKe3iTBmFOo2a5vOxb/nCcAMYHgp
KxyO18wZuT4NbFUSnnr/5s8/aphMLi76EjiFhF9IWRVI1939l+rI02UPxXtBVDN+qtuwNXO7fBUS
ddfHDzkJXpMyr7lpfN4ji+ZKscDKC39338UB6N4u3GNYRa+BlVwOw7S5D7rRsco+U/25Kt8zVEM/
23LDzwBmI1QQxnlsRyXhaxZTKIVmBUojUlHECU6/1TnUkGe+9cx2AdrKzApBJLKB1rSXDPPuXYO/
vv5lEyXINvFSlpH9I9CYYfkM4ykIlRfLsplG0x84uchZZ36Wp4yA0bepZBG9XjWbX+XZj15Fhkny
ubP1aah1fmmscOj8qVlk4cl80PQF3VRVcl+93LqczKy7wRyFDa2TTzc77k4hZBgytCEZ4y/h8Rjw
2rHcMYwb8qo2QqHEtJsClWSDWr3UPevClGGeAE32T63uhLvEx6qKPc+Uhceydt6WCFauxhKhcFCN
ayDaM7/raMa5tcbXTcmVB7QNJcprFJf9WOdoB0AUUx/E7Os42rpDZrItCTGNfEx/CYKftBiwf5Sf
efTK0gT1pJMZlqo0xyU17Kc6HZTOYjG9Q02JOdj/9zSEb3YIzP6i2zGwH/qOlXqhJBxdNaXHXy1R
u87tgEV9TPr/W7WgHW8n7G2BUYxGkK+hGAKKAD84YjUOU6S81a+ijVVl0t/QsF/PYkzBG40SrsC9
NpkRE/btO3yXt2TyVmHGY9rWW6IjD/86blf2UBkc8zB0ugX1547kNRKulw9D2l4s1rjOFTnABN0W
X4FRbcaXZgkSBKIfQKWG2ogzEwnUKznE7JP14+HpBOCTG7RUuhmosGngs46dqPaWl4/tLvEn072g
iXCeB2YXooIcKWBXTeJn49bH7S3ELLfymI9n4o2e1kLdpKb4wM4uzZgyTXmVTQULFSVFnXi9GaWb
D20ZEYo0+CQsUkTD4A9rRhHniWWGfJ84A627CwKrG54m9PRoPs0CQp2TcysIA9/CJ+kBSbKfYfln
iqN8eNk+H6iplbEPR7HHOc16zTlEZNNZWH+Htco5Z6hRhfKYP67L2P2vskr1/pqjZjISRgtRQLYl
59kKrYik2ZSoHdNM0fZLkoXzmBzhovm1lz9WYA7JxXO+jaIvEGEj+ubxkQtBtvbPqZKmE9R9GAD+
ysaBz4fRBgzmeBq0nCvxh3f1DNKlUkBcM1DfpzGcJN9yI3yUvgYqF5USMgIdbgyYkBVq40q6ZdRs
m1aigDweNyaA7XMYo3IRJN9pjlZ4lkqKiLoQFiNydRAOV6L+zAPxrYyNUOJa0g7U02Uv4YFoy6Bp
6/fmFn5UMDUlJtlPC/xgeKS8mGpCSyisPUt4AHkluo/BqZUhC+0g7ZFLgcbTSW+d2D1b4r7tqnc/
/jJxSADPKxK8zwr4HsXRr/Vjxhzdl10Vwu1lcGA8W7QfiQed8y0IZBEjAf+atdevGd8vODapJKMI
TsfB9XqYWjfhfAo6w8waFV/50OhK42+MC34fNJA/oXxAlvCl3FlwiVO0cBrw1Eb3xtQIW8LGaB5C
7v3qq2bA72B6RKVqeLovTvyvDkNjUtWaNkKsRKcJmkCUqYJQSXPbE3W2V+rOcIuDH0bYxlCErgbm
NBHfqB50AVBY8+Svf8rvDVLfqUOEuKpPDsnt3bGQjlzbzveQ/Y8Q9a5+7splZl8DdgvQEnePruGW
thkAu6RMAgLl9urWOEYircsiBGNFkFOAZ+MFc+dywEa5lIucqLiZSCQIktupDc6gkpBMA+QNVfSO
TVEeTJk3ugCBbDDWqBnmgEz6GkIwOSTM/S7Io7dcANOgiuPNOtCTGVTCJv+15A4kVXMQa8Ys5dz9
HT+h7IlTe3NVJaFKfe4pBNAzbbwD6hzO8awj6NQp+aQlsyrqWwOt8gdsRWB1ZY5gs065QtqHr6bC
scVR9+e8M3K7ysRjyOj1xGA33r1bQktTep7MrmUX8uX7y23Cs+muwKzR6IZsPM8alyWuBvdM5GXo
aZOQjfh8jcLci0X0Dr94Le6F2bL9Tsfw3/mtrRzDcCj5MtDRyriPLrgzDeCEDqV2taMwCO6sdepH
cnYoYZerRTFF2lkXIn8xczOw18Dfq0aub0YiQ30NY0vHB6PKqjiKO7OrGZTcHytzUN2BR9FdMwfL
QfDbum8NMZbDjv38ZW5OMXKrOp+BHyaDzTeWdCDX3fgjHEU77zNHqZMU9pf1gwwlKC4zIn1suvCJ
5hY5deq6PP9vzn/rlQZOU77X04OJyqScBOKl7llN1eErVI3Pko8f2R+TAB/4LtzcFbrcOASo2R1N
XHQgCTK4nbNnwsZNOBKYjS8HNMSGC1E9rdPRN7SYFtkzVKAAO6PIpLvCVsXsk5TDW91qu++XlzWU
m8izA9qIQNracrOGwwsohCd+elwoq06JV83gDZR2GldLNhsOc/R6N8dC5T+RHNo3DCkd56TvwXCT
2Y0ahDEI2sUu7TI/b4K36vJp9JDYT9CNgqb8SUSufvDMQZAafBGSBokij090vrmPRAbCyIZotNvO
+ilhbSkPUpSww6CkpkvZkHnTG/bVvZkmejXdyFEwTpO5caulhhV9mF5etif+4q342r5PS9bJ8k98
9yekuzM8i2JQ8R18YmF50dpSJ9evyWVBZgPQzd74b5qB7StzsTiod8NY4dDruVC9ddL6hUig/h+6
EI2rRqmfseERZNht3JGQmjlbV/95fKbzG5aDoQ/93fwofdRe/hABUyBwWXmbP05F3ePvCqT7PzOd
2ywv1ZQq6xrnZADgD3DwuEU+Tbdq6k15jPf6xvirfYqOEXOh5tC4TGWh5I5lmVzWXLkTb9WvOCnq
LkC/4OB00cF010v17h3nbOZ4z7ZZBqwgRo1m26apmbooGsvjJFseDXlTqOho2kzJibyyxsCpf6oU
EJMycEZWGJiI1/I/LhE3F0UsZtMNJBqLH+vtTU2UZK9j+6cLznIwRHptbMHdPXNNY6G5zrrA1ulu
6l3ZbRfW/k4sQjk5irCbrIiG2k+GRLiFSrzCkWyS/7bWpVluQXgwiW70QuzFmh3qCia0mvlXa984
pMlGY2Oen9vJCS1dhunTpFJqq6eHcpjMM4UvLhrn9HpXm7diZXuP+niMfo44ZT+MU9CoIgRYtyXw
JOL5x8V+4Q4K07gmNm/205mibNSriRAGCjQYqkvq0CFQvjNT9RaxuE5q+4vqYLcksud2fa7qGp8r
gXpp/tp797oF0Gj4lKONER5c5kNpya1vlpDLXigOqIaTSIoYF065mqmpmHyHonFk+qFKlx0BfkzK
rAtdu44fmTbW0Fyc0dPwsPTCXEyl750x9XeIaiJfMsbVz2GYIOKoHWeLC+Jvr3BSbVaWGW6TTCZl
e18T+8pfgVlQhaUtT3gfRPN4IAB0hYQAeveqA5dxRc5zo+Bofr+p/QfPQcRYqpdirmd3CQf2Aawe
Jrmx3XsClUE7bkyjVnqsFm/lNSfB3n382hMbUomDRAO7v1QIgglcVr+jeawH9RX7CL/lXcqUUS4E
Xh58J6oZSR5Um676YyJMEswiZB5fmEfxf4SOwplShh97khaSIq7rXbIDhIDbQnBn5IURxAsI1r48
bDfJ9/lDIT//LGny9HwUolZo4PQ3LmkqS76WY9Xu+BecoA5zLUjFi+O9YzFd0ZvdFvbiU5WCSicR
HaaxT0EK2aQJU/xNwrjQGSjkAAEdPY6IJSd6BltlxjGgWj5Z4Yla6cLK/WBmuP03s1c3CRSaXU1e
zo3MMkrTb/b4DQajS1BrZ/xXesOnxs63t0/M8IXBT55fwgIq2kOWyJ1en1VeNaPsqJBTZlDWoCtc
gMjq3QJ00kokpa8+2ZwoEJhhIZlphbN/ptVN27nOP409WzDPH0woCOZypN2+XSeXqflJ3D0xi1Yj
8NeNDDHm62gXsnprHlcswwG0xvtgfs2utag9N8+vHMD+sgGcNQrwRJQUJqGILcG9n+kFXTqKdnTc
aTxtmM6sW6WvaebTSWG1Eh/MvkI3MCf3a2SSv8FoXzG3vh9nW8HAIpnlsBJDuETG0Nq6Y4nlLPBZ
+w6rrWIsbTUBbvvMep661f+e8HjcsFgGAb2B6p6TrZIjNDyUILdBF8p0uxtQEPJ3jqRvKl1Yzp7Q
9Nqo8Ll2l0RlK9mUxOIC7hqt49VSxc38Nx4oX4VHgM/XqwlNfqpsXm0yMHLaY2FWxoYYfPkQlu40
+isjJnrGYUpUuNJZldQRe0nPpDXkl39V9kXDo9IuuphzLfYXn2pcU2K4QuzYa8VjuKeOuGWvL2bX
GopJJ9ipC/i+rGodKgJ+HuJCgzhSW/Mb1r8F4+uXcYpFE+3PMHNQBhtjrPv9hfrFnVAHDM/NKwjK
Yp34yE3hcddjEQYHlz6aoNHT1YDtQXZzzOtU+0HoAe01SE8daCTxFd/2cmAQ+Mf2hBT0kPZfHje8
G06ofGo1rGaKXzknmd3QZQtuG4hYD1alOA/ABQVs56L3N88NR2VD0MUFNUb1nyBmnFY4kzmPmoJI
cGde+AM6W/WZH9I+XPQonMD04ckeUb4ciS2bDxlhCSFQCWp3t/MjG8dMbNmSkUrNEZaid93oF6Zd
CDS5IbqRq4v3CkG2ps9oQVsO8eYpV0Uq/YE8M+9KgYKKef1P4b5+QVx5VSvoAdqCSi/YBBipNpgv
IPD2bdNqIQuT08KUOnpt7YyH8+DkwdYT+55V1M/We+zUmPH23rBTL3DtzZZXLH4Uyw/IFRjUTpg6
oVXeaZCNzbPPzCnzjc/NdhNCH0WaAZcdoXd4nntkaH34aT879QoqlKut7WZR0NkyAiv1KYSndqcw
vbz88mZO20bZywNqncWsmpZkQxnD7fYHPABBQwp83Q6yMqCaXhkr0nOgn/7l8CnwdicHHxr9rdw3
bI05dc+Y+wIzL6W+TI91ecExS9+smfATGgHfxsFCWw5C1ufjzIEr8JHTXIv6UTowXO8YbUQBMIt+
KXqQv5EZs+u/pHMd5+usFDMXia+W2YvJ0nicdWpdSZduFjBjqUcsWMalQn0MXcX5td8zxYPT2lIa
axfGR2eBC0BRSz2835gfLWlm0qpWxvAa07ct87ln8Zj4yXUZJXwNZMfqGnLk/otPUPBmS/MP9amb
4Oxy0YjpzPkLXFVuNnARztza7nNVHwhCEuxqyYXrYh8lFhiEgkK9NaghgHkz9qAj4cp4MlQsRNLQ
QyEnJPxq/qrpo8s/XeMWWA1ivAJfcnBP7mfArMFbw+xqbcPezMDIz7k2wmlvCjyWgUU9ZnjQzS91
i4zNTNPanfINAVZM70LZcm8TAz9zS/rWTgUDYsRUvHhlJ6FB2wSQ000JPetFosRscAqcLmsqOLvK
3FmEdWZUZZtPm20H0MpzX2q/z3oyylypLK02cjF4lw2dcFdZsNw/EfIY2t3dyMS5JoNts4QFLmcj
nvfqT8LdOFM96Zl3Pqtel5isLw7yBr9LN8m9kzEj8dciemczKULxl0ovViCMbzpsDGFxD2+quk2x
8ZZT875w4SzD03yOeqdRjCKxaTJPQzEzo5azswarhDgtp9Uv1fyAABkKTnFdee6wXIPvj7LkJ0cC
88/ZlqxjiEm+84/pxhtSNQEMcYnMpXyE4ZRBV+dcyz1Mr6qWDqPIMF8ElBHkEybt0rCwUOnTmHZ8
DhIu7TtPeGqUeGz0ZdYU1K7hsP3gXN8jKFTthAtxnRbrgvRZhFW0WBoZca2y7z7s9BmO5U48F7Tz
x0VlT2cr0fXCYFpbbSB3KdoJWaXMK6aJYrmG8Fs8BOncL6CwS49fV7GJ8czZ/oK6OckVMOCs8IO1
Owm8vQKA6wWCJCPPvNBbYkttYie8V2M4spuhf30p+jZdCO57BVvJYpupWXKY2xDRyNwfaZBJFkni
QGatbVCy0wrpHr57xPjAMcN0ZG5tKf0M4gLebuUIDuhdH78OqhJAa2gtk4Q5QwZW6VG67XAJexEA
F5l/pI50iL3YL7sG5RqBdXM8fawpuZ+bCfF7YZuWe4Bv/IKR0eSal49u2YvTaIMLJR49jaZY/9RL
6BWzlDxITguuk5M7+l6sLtc+y+BxAeKMp4gb+jAYNUCvYtY8McKW9eAd/MDZ+cZkgmB4mueJ+8uA
QUi5hA1jtSXv4yLc/AWtEdHD3nyDH25n8ds8E8lm2hjFypEl2NZpbez9/WBLp8gAsghFxNBzqtk0
NZqnFWYV2DFD+n6WOpRVGrr/Sgk+sIsHTscperRsrYXuItuPuZwOtzKbvLx1a6mmgB+GXNhAV9fL
ThH65yTF6WDlpZJM0zjRtT62QBaxnZEpknOtRi1UHaMVxp657BUg4lGUdcVjIJ24KmUF7H+yI3Od
LcMAsYqYjWiqY6B08LWGg6D1Y7lHU8Dt/JiZAq+Pi9B2paW7ksKuRyDiDJc9o6hIrJACoRXZLfj3
/fywB9GX07GPTmCmF82PFG4nq7TMhQEIHAz6tXur8PK9VsuEtVvVz7B4do/eXLc+Bssx0Q1nIAn1
h/qXd6f4DhjKnhST/6A+cagrMxtAjGHaU+Ir3qLySoEq1rJM/Qm42vpaRWDihIhCqwy7H7ZNwFrn
VlFSrIrscVFaHQKY13ikqcRDhrTe9/w/PNd35L1NcqIAXdc5hei7OPUW8fDLfSkOzVGEDyfwCH2I
MA2JOZ+iqpZ5yd/W0jkQmd0dIHTiDB55z+aQ5ikU3u27xDmPIiBAxNieLgxSuo8wR26o9XyeSmvv
VRe9YqFbDoUeJb1VBxNjJ/FLrZUiNxa17WzQDngO2fUxsHNg79lMTN5dQlVYu5FNHztWtuOCuQmh
PNzmcn9KZ187KW3Pe/5T2dQw/CGNLuI207ylcG7M2LNx1CKZPuHy4t/ktgvMk3PDJBvLabP3vX36
2OD+nWusllVP/Gw9jP+hYWUzCg+g8uh7zEY7kj8iy/GP1hFW04VAO/RuKQ8TMpAUwqcQZFrrMx+W
XobKbiwI1St6fr+at8VI1Co1XrF9AVOfj0cmg+gklkaDgtyUkbhhyYkz6ZxS8WWXbjqm5HL3iB6Z
8TXJNQOareqM3tQJGqJ9F7mC1OMZ5xNxW8LVwCwVypWyJ6mIkFtG5XPc3BtbNvOkXWCkf3gMFonh
09JwAEG6Jad6PjS5wr9CLhBoev7R6xAu5pJWL+j1mEG5BCMAeCYS4Usgl0qUPLi6PgybBtp7N3VJ
RZIDlNHSKt2GyH7i5GNzrUQXRIIWyILznv+ub9rrZkxchDojQb/UU4vevrImtIGhnjPGhN25MsUs
V/vk6nB8END1HDeJPsw+amS9IMB2ETjd4TFj+yNfuzhG3RnpJI3CsBo7esFhoD4fAk5y4UfgJtMc
z/syVGTW1oxCKpDaBplYc0UU0XuIeZmqouXE3wKjMcla9qPi5EaMhyGXEXT0BtHT4CtsKF+YN+lP
3RxWRvLgvnl/6gq1cWRbRwoieEWWo78OFD6FCDctk/u+8xnkNvMm2/v6HG/37QVZLlSujl4IyrkG
wXBFi59BlkWcdxJXuXc7oYgaEcVK/o71IgWjBzRvtAiPiX0OjDNdHvbSjiOyTJ9zZEzkzaILTKhX
os6zebnR5ZQuQ1ckz8DDQP2TWgw3gRQENB1Yubwq3Y3og60V4M89JV8Olp0s/d8Uck3fY/furnbO
t2diIihrtJ8J/Nerv+9LHzGgcuGlAhR2k+PjYyPiJoX7BvSKyDctvE5N9Md86sUH5SDkU090hdJD
FYVSTm46jmDThoyjdIoFejiTHWzUy6Onw9p7+2GjJP3AWuT3SkFc6Zpaz3CJeV2NeQ0dxOF9Ibs1
C/CRgB6mIMIGquJNMuOuspjmjgsv6+Lt42FqoQg7VTjfpOhMGxmoJSK1160Mxka5Rma+O1Gs0dY4
GYxEnUfAYM9TpUWupSTXuj7tMT//DAIzvGqlBo3LtfGrzoV9+sTf5KTyDeLWWyjfJ1vx6/PoNigD
K9ZDmaPK/kcU6bP7sV35BaRfpt9sTZHOIvYAMVHTBgZHXKfUd7NZbwBnzIY5BE11UHZuSH18XBup
E+IgMrHthWpxpzBC2VtlCw5hVLyE9NQm5LWpjyD8F+hEjF73PTxwNTjsXvmJ0fOA+YHnnZ8836We
tqkx9jX8YO0wtTsaVPzbdNVTYzrDvGCKAI9HqPbGxNTYCKf7Ec/x/X1ClLU0u+5dsk0APEHre0bw
pDokIjb/D5mRdEl58/dBwFIKA8pkIKkdI/b7gdqD4YMjRNoMsnT+wJnK6TfijfkPOihvSOAkcXeW
UXP26mBwYUaO1xGHDeiVYNqOY+/7PQQh+ynX0DiQuNDJecCWun9+SMIH5mbifa+2alDXPKwZCv/C
EWeZoRZ1EQ8nbeC/iEgNijKW1+aybnoP/Xkd8IGmaYykKaRrN64LmFwyeXMwg3aaFK1O3+oZA6m+
TZ1L4EClgXNj9K64xExhJxcRnD7B7/ie3ssoUHShIRg4kvRPjna+KivY5M/UXbuVaznq8Drb/PXQ
SbCyE3Wn26HMRP6PyiMOFveLL3dWNDgrcgAsBwxCjJ2Lg/oKpdqxNIR2pEKi/H/83WZjtsOqX5lZ
2liubMDhzAcWYIeA9PibnQ/vis9SdSr1H8LU+I8JEaQCx/m6I+Z+SE+3LVyQHPkBtPyaeDukqm06
wimW6RbAg/OvHPZ6oQszxuBO6aF8aEbyCQNzIpzpm3ENzvxvF0CitkG/evx2p7HLcjJQCbxdUGIE
JPA3WLmpweZbi2fM7BpzNHeQXBlnz9hEbKfPIxxLH6g7X2o6XqpoS52/coqPyvrWP6UeniBIY4ut
HpURRO18KTzpyQy9bHfXYwqkuyzqGWGv7FE1j1PpcqiY82bjW6QIsn/DodBcy81/PLtjGF6JsTn4
vS9Nzo1XKJxpXn9C6OeuF/WPHpe01+vlz3sY4p4XrQD3RImwxuNwoCGqVoTHMEG/e9ZHLhQ5pn6h
DOWUkIiGlLSrgksrm8m/sEbKCsAMZ8aMU0yPh2rKMrFZ78cGTxz/QKWwLv5Los5ELtxFy2rNnBjJ
NZAd8Fc3yqGyRy2k9tWebWxpCNzZnkdaYwqpuAImL2vEpLlKrYlIyNz5SEtZ/IMrFytw2VLddb6R
/XZXTMVkNeSfPGFmhP6sdAL9dmnkCRuum+vBV4XEredyGpFYz03UFTpDRVSV6dBoDEqkd5XYnHTL
qIdDDsQk06XFnFUPfgqShhxXaGhDTQYEXK+QWa7ram3rBD10TdpfcEHcwP2KU2Lc1hSUjDzlzd9q
WPPQLO8vFEqKnRI0Zq2JCeD1LYfr0HHYa4xyWr5NNqhsC5M7Y5kaSRdchfQtM/Tarn1k/pgCxEMy
vZa9lF/0VWbsNMDM72DfTI5POtGczSE57IrLhz9QwxtEH98hlK2/5PM9pRtkCt6Gnavnn5AHjZ+3
0yLwN7/dwdbx/Pk2j1hIbM2xk63RlJQVpSkgZrKZErVw4t7Tvfwi+CsLSfkcspzSRh46PnfZTSbm
DgQeKBC7FxekIamhZ8WbubhYCXd2h1p9ITRJNF5y2SIcKCCGO7zK+J2t6FC3Tz90YgguVKwEsA7I
FK5/OuOSNigNvUXXRXWmtxlu3qdM6FB3S+Gx+4r8qwOliUn9RZEi2YCqjaFADkZtRGfK/gmsdh5J
9P+LiZUOpQ6vSj9uV7bTuHEbAuHmYLhfZKAue2ZVjOpM+3mBQIjAjwnN2E13be/uf43gTdPf1+jC
jEh3vuedrOylGoTapDH1DZkI1uRZBj0wgAtGYTNfVwsiKLvNqTtgVxxR6naGLPbdmsNvFl3vmZhM
TAUBPRqPBIO3DGnCW0Cr+f3UwhzsfESDASdeqwT0URRfn0OK1J98i/fpfIcJ9wXC2CfRmIad5JQ0
NKhvn6xPzl7OiGe/EyLbXOwgItdI2G7dXjH7F9NMUcYLFL4ucJnv7L3KzBJbUnNzm9Ed7A7JVyeM
z8ko4VykpmyRdKeb2ruuYDHM6NKfvLysTob2bgPsuOlWi6wfOpUgmLp3DnuFDXHjOUbnQ18owIh8
UEkfw/kDekdVRxT2HB8pqxFZFi2f9O/G22bziPzXdJPLrhlnoYMSLajuwOq47jexJrBVSXGncdCk
erqH0zd39wuUTB6sXKfRRJ0zW7TqrlQR4qW4WuayCaKZTfZ4g1kGg48J+eUIRXc/IjaXHbfkg3i7
k1AomTB6LQzhrobkPZ2kHZhSM1t3rYef/QGeNVKKeJRkOzrgPkr59k6tPfimMGykgstpfieAKadz
T5oelTInF/qIA+3EQEgKp2RsXpKfKA3AMEuKPOG296ZRFLSKBid60JgqOaSqYR1NDs0n/4wGlA1Z
oEVeoFy+z0yAsIVEmv+MCYSIrt9INr3A5HEsSgBRUWGqsFCX26juoGY5nc4odLBnZH3EtUQgnJ7Z
pE/rHLrhs86UdcsFVFFynxU+iX03pC4Op2LKPnGwGAL95YPEfzb/SryLYv3NL+sKsx/FkD4Vn2yi
d+3mcWdCr1mEDN//RNTCqerkzsygnPnODigYiwynRQcn7id2KV3lPypttXp/8v+z+nABjEywNXwf
3JbWjrQy8g6Bg8jll3VgtQG9tW0r4EBVxPjH1P2MRGIunp/TsWageBxqriwDjW1a4WpNx+j2/KIG
2OmFGDmZobANUub13tP5Z8sEly//pu/Yg5Uq8Kq0pJsZqEwC2l4KkTPM+IFWvmQ2+WRX2VPQXQyu
oDZgDxE1g0Z2uUerhUlOUWaUk/dF/kfTk0B5J5Jn0/Ld/WtqW8jGIDgeLfv1y/z/fpPE+qooN18X
3UzcpI8bzCFKYIsDcOnzKk8pI16EG1nAL+gN8sR5EIAB2Cd5RnPcenU/5Dt7+aYkEKyNPtAm2jlp
DmBexUyHynzzDdaCzmKb6IgH/npm+iBcVQbE7p4iEp3Zr9DHz5tOThod1KqVWcRTUSOF2wkz2hdY
tezvUlH4s1JHXlFB9PtHRQR/lQUnbIxWmhehYT5MVXubhQvYyip0imN4dGll5nOg2OPdiBhp9uvk
GvAtzUa92+YrqkxgHmtu+yC0hPCug2ULUNc4cN9rbKb+g6ub3maP3XpNbxCEadv4LIQ1E7pkVuzB
M7xZRzhje6SE59pGJZTil6UKQtMpRZ427MkU8eKbMGqYQ/fZEloYKpkVNdbBdOR60KCmJOv6v4OJ
a+MrY8n4H6kSm5KKZtFD0ESZlesLOqtBqytiY6BiXCbXVXMT/bBUC7NRIZRA2PBoN1G8kkK/736O
D/nWwnbiu+lEKzdEXOdCcEZmoB4IqRQdfgc6ZnmTWa4rxK7M6l2ynXe/HI95kwBHn4uVgw15WGd2
7qedYIQiXGpsXCZpvolu+BzCYA1AdMbBzWv7IBzW9iN6ZPaH/moVmJekvnm67zUyMx2hzKoLX+Fz
Gsy8ChE4A9sr0nQgcIhKVpWgNh4lO81CIf+Udm9U4RxsZv0ousom/6/HzOMzd0OIBrLPFTN/7Weu
0os8snvjFeh7IUpmphe+uUbv1Ek+gi69akKYUgY3V+nJzs8Bjwv2jDD6sJtOi7W26SXL1sbZsz/W
Tao5udYwHc3pmpWujWsy3mgQp2KNhvFnHUkuOTDbXVPbUCe39NaSpr9IgtVACgNpj3BMu4SydedU
JZeu+nYfSn98M2fcOQHZ2heQpHMiB0StLWyHXF4yPhC6vkxMUY63aidz68f6cmDuFcqo9ZvFLkhl
NeogMn5tF/6eR3ALqNeznSKT+IlIIVHZQK57vhtoMLs0K4S2MJaQoh5PG7ZNu/ZgzmjAAe4Oj5ZG
+KrOLT5i1iJSwj50xKt47TnzAfOhTjOGAEdUbqMTYKaLkrGIiugMM6RyH3h2Gls8LLSQvKHoEkSu
QHJVAWbP/C/MVCvHJIHEsYTRujwI3tI6uNGeceI80LejmbVYa/0BHh1RHP1pQpLPQes41g4sqWRX
wy3zM6EXSRF2ORH3qZi8IgkYQqKMOrJFQkuUukKvOGtRQStwLcs4NrzizSKurb/0GGndDITGILMO
FCN7SDiWgTTOxwBvUupdf+ciQtB1KQNxVLFcRJFrHeLkNYOQnK/d13uiCFU7EXish5iPz/OMfEqd
CnwgetS97tHYp55d+xkY2ri+oNgVOBsUqPBOdjvaI05ogAQllG8eDFHLSNiDRC4baiQEToJEdT6A
r+toiiYA8EIuL/YWUFZjw0gO2+Ue8InVeXTTtzulY58ONRhXBZ4pziTcLSAiUbosHEljHNnGKD6Q
QBBDGNSp4o2dvlARNuUfpzRLTPq5j3RJnQKQrTzNehweGFXrSo6ewhHqpF693EHOnx9Dwgkg1xEY
rvib3IcEBalm1dfHAukIr6RwU9ZyxPR/9tm8c7plxykoAr/3wT3pfpNA3tPFdfo3Pzz6KolaMVGn
6GR8w+9rk7ZyCxVPDUpC9Q1oLZy+62MdOezqzZ0o+MDJ8W+SsppUVSkyO0l4yZYp4HPfyMOKGrBZ
bU8+i/4R0FrW/NcIi9fNrtpMWvR0YPvM53McY9Robv2b2wlQLmpPcG44PkbtqfwJKZ6Q5lSBDxge
zQAXZKfAyMPlUsrPhQ2yXQSHK1CwemtAp/82MaXeemeUIhbaqt08QAKeAU1mbUwTuh5+FogTRwBo
d+ABoL2u7SpX/422i1l09g/cNYvoJF3vLaFWNsq94k1lATYbuJW78hBKxq4vFvuXNTsDi1PR/ZEa
PItxSjh8BY5aN0amZJ3dFH8JBkt4WmY5/A082soVF60lbd020qraxP3pUBp80pgxQhBqWQ3ZjvxW
+YmPgLO/JaAZmhESejIOpO2Qr0vJ6TfCVLzSDJzs6RigDseJ/1HnVqQjGsertOnpZYZKQ5ik1j6O
s8yYc9aONVF2NTnItIxUOSfr7gfCYhvDYSD7+e1YeXItJH2/eXGNlo7ojRNJX2GXbrila29z3PuA
8FqKsDqNinAraGPvIOGPgXNBZka+GvVpu749M59yg1uYAWgV+mZSPssQw+Xe+Ei2iWw3VGmnPmZM
Es1ANrxLWCgP9/VXVmhpOHRGanoOZLTiGoGmYCIuDVdtu1YffDcQIzp8A+diuNgUJmbmhN8c8+fW
4s04RMbV+MIBarF7fbO4gI5oKo5RVVPgkVdxd5IkXuB5mn9hwjgAoda0RbgqUQ9v+uqwgXXuB4yU
oQqfPmD+VTXieAzbdp11yZo4prTAk+f0OKFiKdcfAo0Lhk1JcUNFyy8KCSFZKzxi4D2Q2TusDUxt
AtwsynUYP1jHOYq/85fXsks+/43WrVjyFDxKF/jbrx0XGMGdH1lzjXQVS+GvUNuFN5WpDxS+JC/y
FLfJ9FRWq7wj1x9juEnM/YyFBsXcpiT7fPNOW6Rh4JwuQUPiMg8QAA8j0FK9spl3RoitzRE/AMVX
z4JmeMZa7iOJmyQVvejx1nyb80zBnAOcw1yxFfFxM//COti0NBsN+nbCafQ59s8RNvAXfalbusJd
616N1ov6WDIb25gOLyrGfsxSlZmgi8B1pi3hzDrg1dNB03UeXqrE9KkPxQrH+/ANtg3CQdzmZZHx
KbYnZ7wQ8lgf41oh5sjn8S/Xvgwf/rDS+ANrBQ5gn6Ea/nfxhmQjYSwfh2sSXU5p10MRQ0JyB1Mi
SXqNE4S+X4YjJKZKjIWSfMmvf1XEslcKhifVNvrdQ5KkRMh0wsyUdHUGqIwUdw4JwO3JkPjNf1lh
luKVzBHdKO8e+2cLcTA2nP10qYw/+wHxe7Kak+9ktDDNgaXk30rj64RU0SRYadhUyuUWDCzl/2IY
ehj1md2BhAkYUZZOdsSg49WeCb5/UOv1Hx1HDATuyEM/81p57A+2NTYHjXanVv+sM1ssZist82u9
BpCO+t4srMLihbQUZ6XntG5uf9q/L2ujFdK9BP5tt9i0zAXpIrW9iyN/asasHh/9tHHRBCrvF7R7
Uz9WMma8MZQVothfVJ/pApNpvwkg7ZR1xZ3yx0A0gvG7yExlpARchg65BVbniDyr2GICbimmKLKt
CDO8WIXJaa+BJxnDP5QFAV6QoBJnicx8wT2bfrmzJVwaiO7aYGvTbn0RdA0JlwtBk9ut4lv0EQie
IxbiF39EudbMBkbI4kypDOtMZVNvNCplAJXnTWI++0J1IHbWuC1vHdhfXNc9tlseLUkq0rUJ+vQV
ZLCcHGZfv5Y38hgB6C6z045p9Ehkd+pZff/XJ8h0i3S+wH/g4aJfQkcaGfeqXx0VpTGdcaQU/f/y
PuiWdHubkfNKBUc5MZyjFwCLkyXysMD+WLAZw/Q3PEOTo6Wl+vAkSuQ6+Y/53j3K4RwTKRkKj6Bs
riAwx18c9foa6fXVO8QpvDGN/H1rPQNm+kQR3KZaZDImESgmw/XU4bDee0a3klD/LZSyVSCNt6ao
Qvr5h4fn62KESQodmWxN9UETBHfuV6iPkRI3uSyzz5UVmQ2fiuZSYLSLm4YkLsJm6SMumNe/eoZQ
710/9IMBMKVKCsnSbUUA02EpiG6FO7XYs1DDgs0g7fpaqrPfzVPhrMdIXaEChgtuT7p9D1k2N9xO
K7/RT4/PRewoMGHh9zSLpGQEKZmTDnNJOt6Ae54zlF4/LZSEsGMVf0OQBsZlwRf6GRoNH4b5a+TY
DnOF8hxQD/uUWMmYn1MMyu7F/VlSoMKano0X7B6YvEr+9NE9eIPKIAFkZuGRcYpNar/4HOeobZge
pGM6FCRZBBwIkPhArkXzth7pBlnQ4gJUimaknnsc0jCUc7NLyhd2KRfK+XHaHJDwyOQ4X0eG+WtZ
KbWuSyYmL1ltLs0EXUJmBbArSgxdU9sGxZRvVR1Y7iUt+KKB2Pux8gHPVe3NM4rlGyD5iipkwhsh
ThY3yUEBRhKmJMG4x5VyZn/HjhLQYv51xvePxLJ/8BeXqkAyQktKpK2zDtXDESOUOluvdBQTBb/L
ZDZrpkQ/kG5s9kvDe1v6l9U9UpAykZQGEIVwZJ2cTWweo9gPqaygDEZoMTUfBeVpu2J8PuqsMHJ0
/O1QWyoxBhmFd7MpleJJtRq+dPqCpRVdCSzdVFNHI8Ck7uoP3UBGWJqIiZYjqMeVZjxymAlsgwlI
vMcProyv8X+0xAdHfzSD2mErJbExLEWrBIUL9az5fyvTl+BIo6qpBfbcvY7/8DdC8ilbAhJe1fhm
BiPCpyby3UcQDcGzdAuql4aFi9v1yWS4u76tdgnoB/4BE71b8vpA1fDg13dScauK4ISdc74oNNkN
men2bqpTfpHv4sgTxh3AyNep+iET1Opn6i6w2Iku1fPCUWVDHimvQefPqM9DxbcHN7k8XIDRBKU9
SEHLNjNwLynKmeZVll4NTEBeywCoEllarF6HRgfFw6XXClG+r8UN9iRIK4ozu3JRLfKje+bghoPI
vdt/7XyE+V4BpaxXAXPvpN1EWlhWp5WfZhpgjGU4VHtvDWqfma3ryI1+jbTRYCFKmyMnjvvY1qN8
Ylq/+dQ4oLq7qObIW1hlkYLoOLF57R2IZ9Sc+dqoPv2cN7FFtPNzA2ikfYnTNcwzoOPEf31xSzis
bVRhF9f8GjU6DAUgWrBoCSdR5tPEklX8o3gE4FHlpCDV4odbBqbkd7hq+D24knKAc3n6rAqxKG1M
2l6GulahtQQR1uDTBazOToJAGKAfrZ+0VqaNRIyFwJECD01PRR/oZ+EEPn0k0P4Dyd6a9m9q+Z9w
FXvxRNfiq1zHzPqpYfXSxUOF2xnr+3VjAkXwx3n89faIUkD4w7BovImGXkUgvsKBdFxeJOwJaBzi
ObaxBT9e6cIVzfzAXuOcpi0xdSPcBgc/tRqnE4FVwnkw6r9v93QiO4rNqDP7tAQim+CSILjQzBVU
3GKjXCHUPV41d4JYoIXkcA4xwUhwDx9mKawNrhcvzrwHvxWhKJAj8I07P/yMhHLQhLUM/Iqfaht2
uLClzh+NXNbUVctqTKFAmwc/qd4jJlFU3gwIeAOhh9bcifIWX4H39x3655V0tsOVAdTq94s8OG06
JWVKtA97U+0ZEpiEAoW7wysAx1vA3O3JfrMM+usOYv2XV/8A3q9N2GKyqcBwvq8x6Qcu9d+DcVkj
TRE3pIn2C1eI4kkmdk6G5aaybV7bYTGc36v/OkL/arb7UfnKFMhyHD4El5cu/nVco+EwFVeAUJ2d
bP02wfoj/eXGjHlN32aSeiyrA1V0x1g6L9L/WggPVrqfqZKN36sjj1ffsH5eUxusI80psbEGKVLl
lh0rk/kwZ1x6QoAKzLHKutJwiJj74AeEdeZnCF3lWM7cylA7g0vpCUmG5dAD7htXMUb1n/Tdz/OL
BuEH68ok2eQetNBrosoPWjFsq71DauDlV6Dusli/51IZp8uclfQGSj970RhdXpZijpC/RiAe1ToY
yewcHtkwFA7qGOcgIysdCTLrApfcL3PVij5wXh+14fo/TB/9OvE615AAZnXdgo5rykBVppZBNj/f
DQxu8wt+eSHnMsLHK4uHnCOd0ZLaoPIgIlxbwPooJ2wVOXV24C08Hm8OKSiMe3MuiVgvTAhG66X0
nC+CtAa3mUnnWWnUPNBdDR0m8hGPYQtOoJSMDtyAyfT4rwj+0+R8o45Jw2BCpgizZg/Go9UKyv4y
IarlsdZ9GV++3Ln39M+Ycy1zNv2ZACmti3vZpbz0gALJhVXaQkDgsdo24B88Kikzy2eW3If9+SzI
lX18HZI00HWGDfkCZIfKupSy5lshVQ31BhIKm4LYywVDHqc/c+JEzir1Edfle5IqnKhGreM2b03H
KAIXdATatdCmh1zGZ4di2qGtKBOcYmnyqMPVKd0jN6HZ01i7phVaqiLHfpAQVhxhQAMqlrs6EwaH
NFhSueJXm7sQg/iOMy29zq9kV4Wj4mAhJ49l/zInIaddzbDepeHrBS7Q7TNeic8ZKCOz24P6U+4u
hxexE0C5f15qCSAoUQwf9iDvJUK9y9RybHr7FnAAfn7RNpTVk71oodRwOkOae1QBR3akk+HFcIIM
2njEiF4ox6Rge139xN68MMrWKRZxcgai01n5T4tPb/MPncfQY0x2EhkcjhC3+b1knnRNk7lEr5D9
D2dLFvQH1XOQb4wfEe+jx8CwG9YmAq7PAo7aG5MR/J3Yy9V/VWDw6P1G60N3rOu1ISdldQ8pYfaG
yhi63r0Hu+PEQP/2NUk+YErf+JOZWj93ReM+Zgs0aws7LDkOFofVkYWD7n3N/5/UOtNMGSl3zbeK
/Bz9Rfwy50qhO2JNRYgu1QmCK10f175fWKYIO1CCKfePKkANvPcdZzN4ZvZA07Wxnzd5fQ2yLHqi
eyJHGoz1anx/bS2OpYqEDOneBl16eIdpKO9LS44Hits7kHZUyE0+HFnz2+lFTSO12z0pP6/bcEtp
6h7+XBVGqfDT4BLICb0a8kwazdmeYeAJybvMr++yXvPmzt7CeAlicC09fLNwUC8ndkKFrkbPTnya
pLyYY7iIWzhNJ/nJT8u75oMdPSyL3Z76vFIi+wcO7W11ScfFZGrQMYBfPr8tQbcJAOs576K6s7yR
m1Xf+gMUIMDKQWvzXG48+dtgDPHEklrMN39Y6HObLZhxshiIpAYHS99p10pkw6Bh84VhD5HYU3dH
RaJZkBRImBK7Bx7ElSpFQypXl2XRic2VhGwfe0FTFkJIulJgP5Kr+vpCZ4CEJo90uojmED/ksJCU
gXTVIdp3SczEwlzrz8lKEfnkP8tGrj8mbdHnW8E9AYLfRW+su6WIbO3RPuR/9xo4V8F0fm7MMpkn
GRBoHTvxEATxV1xsHa0vJDMqWHaMZHhQfoGWABArE0jfEJkxoUngYVD8B3uokVuAjcfZ/6sUvgfT
mV/rVP88BEdoIWjcMPpfQqjCv/Iro5NRGHTlHL2Y8bu7E4oikomuwK3FpnqrtcBeuXSC1jslpwWz
TFO/bpH8d6wBvKQk7mOVP/IYYXwuRhEfIMb/a2NYLMPIhBNetlM+D6HafjcBHHfp26f9oqikKhtt
NhbeBSSwSPlfP4b7cp+avtD+2OJvijfBn8B1wYDYF6khjAApYTD6j4Kv3VPzvjl3aa/5b1LJmgOz
ShYzuhwZ7343iQQhDiu4/GIspytm18XKvdcW6Q9xRladcFCsoEE9OC1LPaAd8ErT7e21sQYGY0mk
V94Z/5hU3unCRpbxR6MwRjkIyNp/5WYHtg98W2c3GFu0bfBrTwVvhrDnCCMPY+/C+bd+9lftlmxM
TnFmNode8+p/K5VmCAGiE2ykT4ZjWcpF0TEPnz0iTA0W2HwCcb2tfdqYovtwk2JBHXmrm3DEgYTy
VPD+rrjmMMnTMOO9MZb3+nBp6xPi5eCUOdhHzuncOuI7YR0mqpr118OjS5XcZ/EArK2ExF8SGWM/
HEYVeFmTUSlgJPI8y5UtN0BoWuuFt+1zBzBerduOIF1H3g189j7xe3jVxg9I1jfhiTwOlizLVG0F
dQQlkGKk60XV30f2hxZ3Gnc0EQmjadWaQdxuXgkLJs/5mss2Uu+FwTDnq+lT1kCRLxmuY9jtsrT9
8iBbDlvDvl2j0JnhDVYFROLFuNgVTpQXlk1v6IHxrUU0p6TUvGgEwOKvIdsjWv0a+lVfh9S5DQse
FQrm5pebGbnYoyld5f6ee44cPjbVhbWP9DEDyYqPoy+d8tDt6NWPfLmCu/USEAztsNXZTbOnImWH
rPLSyRxS6xd2g0oEiB7ErCT+x8352rwZTqPVcjSTpiC09cnj/apsz+ztnON0URpoBRqPWAGJDELr
vBy951texwmtm2++U4Wg428c/wMjWWK0Vh1SyCtNO4aTK1rodNIHdqUoaD1U4/ub41aLdD5bz02z
jiGOw60I5lmwKeRe7QoroUnlG8ZWYyEYUvopxkspQ2NYk3KhOkm47sd8kwqA+9mA2iAxQ4VEBkBc
HYZfCiN9vcz1wmukq3GbK2Q+ZayPDRnYn7jw7nmGNATQtBAUksNx9XO5v+Fr6hoK3sEbPmE9bluj
AAidC2p5BbZ+bVMLgePdxAkpR1bR92K2a3Dl9tV/IrU1gxCpm/k1tULNSIhRtyjOZ/j5hff3ioEk
+N5LcwZGozr779lmxdmWpegi7CwSwSuicb4sBmspJgUt/UbwUiktuVnF91MNsil5BTtQ/P0yKQOV
xi1GmkiqjL7zKYRh2dki50LucABK4Mr4a7T2O0wiC/Ov5v3zy6EP7uUzsoYDwuaUHC1GKNX6JENE
6WvFKgcbAWQqdNkQUvNoWDf2h5E7pEr9Wbbc5xsS+9ai7viLVPZ8cQF6OHOsimXBfwG1Hn8V7TJz
N2jpAdq9IYWtuwa4bnj5/5ZdQuTrEeDxPDpVl9YeAotAVsRtWl3rpoMJBT0Buamw/P+q6Cdv3IsA
Bsyi+EtOhACN6lWHFzZLKRUwYmy4w1jukuy1EjR3V0cd9yoz5tBoS7mKPEgK9qbsERX0VdvnDTyW
TRY7+r0U+YgVNv3P5hwTs2vErhNYUfbXEgBc/DG+8HHkO8Z3n65/GMo10hpJremffxzeYrdZ1ZGB
NY7HSIQiCkKD/d8HUba9CFqa6xmFRd8p6nOHM6eJJHHIEidRHfGkN9Rg1hHuOZGUoogZY1MrrnLY
340iAgRQJvvNchd2dM2muEmnxS13Wr48hwMroby7qHy5XBOhi7ftkKkKkkmVhSAxqOm6Nhi5fZe4
KdaA4vjt6fSs2qm8sAqRu2f0fAr6h2mkpfHSmrXFx77WlxgsQVXGn1G1J4CNJztNNdEtUZHt7BJO
svidrG5n3c9Z9GHEXAASvhTzbjbZZnbJ2ZwlVZwnYzSSdcnzTLLb1wTr+12j4LqWzBpksIgGM32B
enl7wNCIrNPO357XwTdM8g2vWq5Ds6zM6LPZktjc9YiRQKYS5Jro9f8P89aSvfbGA5TQTRxNNIqK
3zFO5Q6Dcl1x4evcQP/0lnMmKPSKxj6y+dnXuTjn7KTYV0Lq2yHwwgOOmRrGWN0+zQwDYs3Cl9dp
0im9uMpI+JUwFDOYAa4HmlN3EzKwYrJf1oxoIRyiDLyxlVxVIyicmHuHcA+2zBIjWuLsdpfRXpL2
c9zNQLSAYqIUSbA44suQDcbyRkgdrp6XImx5/GrAPQ2HiEEHvoq8RwAq5yV61tl6cCpj1yEAqh/Q
XJ1WqAb5T+SkD8F/6zHFGfGeQ0DSM7Bf6tKErs00VjZEC04zkSQPeb00P2eYDM6PMLXY30EJRSd0
Gat+sPwPVIWwpZOWkIFyVHwKfy4pRwJHIr3kHFiiU0suYDcPac0O+YNRQSlO+xRQbmJC8mNNBg4j
URS6AWfCcLgY3mdysd/ULlrUY2Lav0O7fkhV6wegsvS6FrznokkgswPHhcztpKqqy20YA1+/C4io
3nL60KMrmjnwaVyEbWXxrajPTtSEn+XEpsmh8bPiT8/9rgblUn5EWleoJvEd+LZUU+mcpCa5yWJ5
2iNBNUcgFC0ikI18pADX/yO6mZpdoUkOXyR6Z+56zwIJBCTBS3lvTdzBwE5xdH/Rq0po4DpEf7Eq
PUO0iYexsJlC3oGah5Fdlr8jBXBURHZiozfxkNXpg11/YLNltp4bE0y2P0I8q/8HtnBL/QoAsKmL
dg0ITkVnDbuPQivwM+xqxoWe69a9KC2sBRU4Op33Xa31LYdp4nWH+4KLEM7p4gxWO3yYQlhu7iTs
qy3yrZImKO+2+K1VZFrvoDkoZuUArUMnjzeKrSsvX6Uz5IwFn8FHvhX6nHoGayuhwrmId3zijamW
udnTV2cnDPrDTc2icBCMQ5SlbGqT+VdncFMNwKMUzwP+onC6Q9ivaSruwuz49nJ9GXQM24er3sN6
FI4xQ6vKOJh5sSdktqCMa1YeMZ5PU9yGFGUuUI6jbz26YF60LzgJDbwSU8fySVhuox7XrdZWpgtG
/mGN8mBgMXHwxlsDCJyTC3A+BMalWdmYpwnoMLFiRfUc4SLssUyDE9Zb8jJoMMe5Q3XTFrLHPOOW
u0FMtyGTSoIl3eopbQpIDEMEwjpteeKfGu6lAKVEzR6OhvY/T1/GAzy+2gMkoxOFi2+DJmAhXFrZ
ZLOr4gqrMp8R45mtrzwlWE+j6bwJVh+X7as/vq699nrFAKjtr9k4Rgc5cQ79h2Awwt6YNHG/RWyV
MxcN34izeoFZ03MEG5Y5eapUz8R1niWTrJ8ZaD1DdW/aiGR6pBMoAwKhF3v55cNOSd1wwO+Cqnti
zoekZwOl2SiHydEBSizHcOK4ZFblpJVzs/fzgMwLQt0CGafBwXUMWkvIscAGYxrZn3OQzLqGHfoG
LN/9ORSXNps7+JmIKK8aiEjuOlGccu3Eys61jxcTacioLaQfarPGvZwtqpkz+6WQ7hZjDsu/rck0
IASa82Po3tKqVJG2vF2AF3PKshMlWOlNdsSEG0DFHD7InHod8zbVZv674mEGufDm8t5ePZzcdd9Z
d/+kmrel1eTQP9S5RA+Jhc6a7JwtX4fciQsF0jJ+byniWuLWf0JSAuxec+xRxsAKh7yg1ytlPBcX
pxkduLEvrGYj1fScjEImJlMsvXGqTkxKPcKBiCpS/74iT7ZY9aW/PHPkQtxlH/ouhiFlEpp/LsUb
1oo4KJ3Jfi5F+5PD1IRtP+/JPc9V4ThGsJxM0HHxFd9nBdHqzdF13jRof9V3b3XutODwAuEOmpgW
n+0VFb3kjEyvtk1NXsXfNRyXnRj6ThZ3bO8p1nJXAWJfDa5Cx3/RqdTyy2bF+DIU6LZO5B3cWLLn
105/y3S6ZEKJEqlcu7KbC4NOOGZpZnovpgXDW9IhucPlR/YWQQKBgqzBFnlUeSLSAIxssjXfOMzH
phQaGi9YsjbGcIOE+VXdTspieHE4x3s7aDdVdFa8EDwmXUKOkffby1mNFoNSdMQUMgWkHP3rjCcY
XbhA9hgexzOkj4Hd57Rtwm1TS4EhiMsT2h83BG8AfHbBI1sT5LU5IOoKu/jOTy04FsnGcGacju5Q
1xjL8k6gLx+ckBF0iCDPjO17r2cjR3e7bPvy4TRu2qglfnSQIXDvhNgC81VLoClZ7B2Ynk3vc0G4
NbtC0F0H3CJLqh+eEF39+8g4QT+yfj7Fm9zkAnHKFFWWNJ0FzIXwW7foDAUjeDU2ikIm+lff6RIj
wwHeovntb5IVMQEj7n/Pyc5M5oerk2GCVqb71tisy1AzUWOd3V1ZlqeJQTCz0ulw/rOpu3ZWMZC5
qiK8OuXNjZ65wxR6ZU2ZAj/ik6JHwNqfG2ISRP8OEcUNG34saJFc9wlgpJFot1l77lBbD93wUVZb
0SWNbfvZ3rpqLjcPprjuq6cVW/3dfI7SOhY9skM9PAkiX9ViPNzhYj9ABiE6953ozMLC0x5PS7Gf
4O0aNYPvyXg6kobrDTGx95Bdk5tsJn8UM7gjnv+qz69G6VVz9oNFxNXXhU1t3VXyMiuY1k1b9x17
r/T9mxsgps7KEFAtmaIZmKVbX/Yt5jy5t2IhXcgI/u4HYzxAt39OEgybhLF+ppR4tY7b24CXRjFg
Lz7JVeId7b4ObDa2gUmR2/MvV0FGn98s0HfTQ55Br10z8ekIAnCK13IzyD0/8Vh0sMmXd0wLxJRi
tLMnUZnc6e6NPtQysaceKmCXuRxJeqH2JB1vonbhsqMSHnusHgN3XKIMKNGN0Z6V6O8kp2d87JZZ
HF+J70R1mPHBuzfec9KzLeTgbrKkltcs7S7aJHjLj50tOTzPbs84DJGVu7mKeRBOymoDVM1aCWrU
uyQD3uzvmY/2nQwaanAIJJbgjp3KcZiRsjxRur0maY3iXwPKZUOcH0kjdT61XhGoNOnpoQS0Hxl4
bUZzhT3w7hsSSjpqpBG4folxNxAkMCyzaiE9JBBwANtfs1S4QgcqCmVH1wTYMTfcrlEW6D0GV2Yu
3C1A5w7Up0kTr8BiBRm9aZIcJzM5lVPt7m0QSkE9y1SrQoxnmcUF+OFxmeXgew9RdNwKY1Y/d13W
9oiHDNrMfjpaX4fn3oMIKMJk5X2Av9h77XyQsidCLM3WNYyT3rvjLoL3U9DPonYZKg3RLQ6PgTNs
oIXJyVArFFr0Q2YtUbLixtSgjmxcm75ALo3s5v/ESTbJAqtMwvdjQ34nG1j6ARQZ3qSP03QkeluW
U29/XCJXEu81DXfgGFZntI7wYS6zk0VNeF0u8JeNezuerm79hB44VYN8qeaPfmYKe9Fd/u0ejB0g
dZ3pQ1Kp5aptdSGmnflWu+ixZNDHK4PxXok/JgNYxF7PEOuNDxCNyFuydWSIvqDUMai3yM0IGji4
o4CD2rWu7qWd0GncGP3E8jcYy0WtHxHm3T4GYfjRazZwKC1sadr4d0OrAkX2dBv7X4EbBJXgUrZl
Rs0IsPZNcLN7QUpBv9bNWT7pyhYQqpYDxBYQBvPT61c6aQmdpCkqv5jto3jjq58ohsBxY39j0or/
nCwhuLUt6Gk90N/PZhsg4n2nJwVzLnI0ypxcuXCesrvQiHY0u3QxJJVB3CneymBzY/wUs/IvJXu7
vWu8RdSU/GYNvunRiGLRiokBNbkzIV1UOOfAhX2+8r2pwWAlIW7gSm0nN5sLiIwIjis8n4p1vQwC
NtNQkjSXke07fjTqh2NboCXgzT5Hb1fh6bP9Q75cP0qwpsU8EnU8o+lb6OrlTDwqx1eWN2N5YwdB
dT5eUBf39EzosaKSN0TD6aiRBb2VXgGrTvi3IqSdAozDojb12NBLaQe914jSF+sqLNfIWJr3YzGT
SBQQkaVAojXiesj2hzmosI79Km5uZQVr25UqyeKb7iwYxPdddLl5TijC8m+RCNl5dJpnRBu2tqhx
Usv+ZhV/QxFbzHQgrLwxJPo8SeWX34wJn0pRGq5jJF9ytdBsMSx7sqOc3J2od0md/VXrsO/payCW
jMsq7jWQTyg9F9cHyHPIQCpBreMCDRXZcGpm/ChRYdHHEgZq/c1xA4mfJUi7r0+nr6j7cvv/j/Gg
OIJUVWDXYeX2PkpzpWaN2pUZsiTvGJYm5I/QgGDDjugxNUkB7gF27avyUH3IP6P+zci6LPBpbL0V
TgS1gb0Tq5sPw4nPaTZ66QJAAGGgC27K82jJg7EyueIyAFLoKobnc7pP3vYyBjucNPK3s8RNakqS
Z0KSQauyBUcJF9cvT32SAdjqhHl1p2L1UW3zylZuzgHKrfBaCY2CTuIYDEMS1jxwycv2RGq3gEqC
JMliUUTYwTv5gIengwKJR/kjwO5R5+PA0nVBZXMf348S46nRVn9KK9nAtXhzo1E0SFU9K/PNmgRL
i55lQAJL1WQSllVRQ1Lnxfr25WgcYttQMLpMiX56yeUVT0pH7tn7v0VXMJzLBdmLcj9jfxuxjKaT
UTTzdA+7+YpiGz1sqzIvBsIrYkDNVqLXaxIqkCL04qnRwlV2Hst6SpqiWiS5IJW52oYoGOhHT6tE
FZZT98CR6d30jbjsYVupiSJEIAxBTQKdxDiB+vws2V7mm5Ps1hf+t40tgkaMRF1t85XjhdhM5fBU
eNLVDJMwPr5kg01CTzIaDPCk6SbRTfN88C/Wl230WWvJHK87P6ZoSVJQ3/+7tEh4F+qC/yNgz0bY
nKw8uj1RcCgSbVDOb9K2KQo6fREa+vy110+ILdueaT4Lhdj0BXVQ2p1mv3/l/kdz1xxZnddXL4D3
sSvNRjxGJeyH+utzBTyInSkgbHK/yBhedpsEsxyf9LalMvUTTPemithYXzDiEdb9NsdU2aoA7oxX
oF6fnfwxTPoW3KB5YtE3VsubxNRfBD9rI/xBg4CKzYDPWdEpn/oWD/cAw7rdPHZEHu/wiy8FtiFD
dNLGG1rEIidCgNyCuA8YNHvX9nzc2XGRCUO7R7nHMMusoa4jQ8mkeOy3/13BkONv8P17KdZvG72N
CdpxoMJx1Vi0/2aEHNpgrDT6mD99RLVBmZEhtk+yeQpmAq7H9QyBw0+iL1vAAt/8KIe0V69Y6Bc5
vHVPrlphUCFsagpajnyoF1QTtImFQh93U2QYlUU5/7RZlPtmzFP6gwW4p3v+rI2QjM0oweDhB/OD
FaY1euA51YjdqJ959apmP7YPgwTaTBUu1AsRRMvBnl+1iXnUj5DIepQSNQ7Fz3xnCZicGvogdQ/J
fcaOOmXLYVsB3vpLdowBXCQtq1SWvPShHoBXEOrqZgwMmhxiBxiU2n215CSKXBGnGTW9fVzNvP9I
eYqTFZBAeX6atnK8hOtsPSJUeuVZt8KyxTsYq/Zo4RPoxA2vWDQ6T9nm5CCQB2tPPhROb/NdlRJH
40iDrZuCCaxigcJOMHWdHP5siS/Kofxo6mNm5ZzfgtD99fMNtVvbhVXqywG119LiBkk5K504Lw7E
HDi5UYdJjsK0HvMjawGAP7CCIob3N36EtcSarXX0PtkDLYl9v5Egm7ZGsQBwRXLWc60VbILyT6gV
/ZawQxP23mbutiOolWXRW70v5gZVKku+RoPn+f8Zii5wIvH7bCQZHr37CcZ5EUpf5IJ7m/PvGuKG
g9In5hvY7K3tMRG2EGJX7bczoitwcId8Pyi9Q8b9Z2nFdn0MmgQ83Zs9auO8R/vyJrK0Bhb+hykK
emGuMJxRjZz2utqwvJqO1AdOuOSc+ydVqtO6pweLOw56heUkS2S1BaOMtYhcpPgl6o46+wdY5KsM
ssXuMmiW4TTcfC2azjzopRY9QX+Z3Mi03/RyAj3F3WiBweEnU92QKOSYJqsTyuAMkwhYyuBNbWVL
sUALiAfdhACfVpr1snLvvKncTDRVnHUyIqwBubkVjDJ9QORmrNQ4F1ym+uXOonlWxRpvuVTGF24K
SUNcudbiJrnK+CHRPFfZ/Gx8anTYW0ZQQCLVkLiGBQjoRAAQuZHY+aFi7rNv7q4j+IgxCxRwroYO
afpwf/l/HBHA6rLK7hDeyXK3ltGxNT4LnweDkuuF6lEL6K92roWoTyQ4HXsqNMQxO2Q/oVSIDm01
vNJwBzdfO9pDD1RJ6UMp8x6K8RfJGpfZ5FEUfWD2GsxGEn4X+ax7GkxmMp2xmqwhea3yxm2VGH01
yHLHOAHcG9exWKKKJMEZTiZUhCbbCBZ/qHaoxpwii+nRJdMKLr0UkRRu9ozEBD0iEh75fbnR+SkI
GpC9Ko+gVh8hkBDLVlMIv/x5YBZhdBMr9NJi66Q973CrKozOiy8TDuKKEGzG2k8ZtBznHoRb+ySx
oO6yvmgYBDqsFChCD5/SV9TqVEJ4PBy0PeuHfv7s3aHtVLUEDpMJD/XjqJxnzdHfN8yPfUyBbuKX
/FeETKqEsRkgn9YsHDq0ZuoxtUrrLIiSBaxflX4oO1GTn3u7RIcXMFneqloVjxxCsxdH2bL1aa5n
sEiWnsQKnNYElsCXtoNfW+/1+ekRlMEt50Wm5VGqUppeajRxLRNb9E0PeLMlrzUISNNT3iHHeDsa
78J6iI62W3ZtWI8bHSPRJ99XbuwykSt53OEgA4p14eKg8AJYkTfBwIZyvHL4wSTe2Xp5/nr8AQub
BeblytsdKnGy1/LbWXlJsVCIMx40Lx/0ed3RoIV32k8LGm+zOMS1ShRAf7lGwdSbF+xC4f09nJ88
mkabmNGMQ1INSTcqFLH5x+gk+vEYgYFJ5mJdXKNhaO3JFxvUIISP2teoxmhATMNoTRFwJFvNBQaR
bHjZLFa8ezJiYmozwO/M3tyg9WZh8Sj3ywtPWRNFta+WSrekTUv/DMFS09fU38PVegX6Z4/tnOiC
EPjgeOaEI+vSvq+zOGaB0tD2jJdSFHHZ97py231zjMw+isPz7dVOp7FhOF/yjRUGVpwsgLQASQPj
hEOt/sR8eqz3FuxDE+Csl/VhLPeHxpb1dGGtqpxsJC2Q9kXMVyRcBovwtJsEZuDyMZM+NDHt0IUP
r91H4Bji6WoX3iGxM87fxLCWxKLf494WSMHsZPpi8y5rt7iUWXbHwGSp4HvwWT6TOSUCQVhD0dR1
3vzb+T+aRvP5a8ZYe2deMvqGFZVcHnump7/2NJLGx/1n8akAC9x0MrZTbyzZuES5DDF/hq3mnp7E
cunb2ZIZZQgKUfZwRB6M9G/I9HsElaSLkLz4T/z4Vog5QYuPf+CRVidqEn/zuQIPKFZddgOgBV7G
X5/awibH3dmuR6FMXWjlkUA7Fqj3w6a7FQ9yPTp3VJpwdq+WGsvyGUyq/SlEnrRxRB3LXeUCkxsN
vyv8PDNpd7YW8D0/2u4KZH/2H586zCqRxNoZflkgFTf6lsVUQCp60AhcMfMbaJVnlXUHivQsihOo
YXyKdHsXO6m7k1GBIS0rUQNjABB0JbEM5U01JkYynzfyw+YCacWcX3R/XzIi6OU2YTAk8kiKIeNj
P20UFLMP8v+v/xtofj1mRiTDsVmm/EuuqMaaruMZMo14YUZSjETFBmKmOOWMeVCwu2t0Hz7RfcsJ
RH4UDiKpGOTNVtA8mP+AxIH66+cV6weYFoZoKISg9nZUTKs4uQaeWczIM+swXittXRvgOTSGOc64
IiqqAc1vN4r7yKkzkK5k402gb6cwUgbvGmeQ8aSUyvzutQSVD1nhWsZlUUb0TMzlQM98T8spkMnJ
aSGw1xd1pLclcKLNasJm/kEomcu/tCguUeXESF3ePJvVHxFuhTjkRwoWW7co5EQoYb6TkEnd0HQH
fn0olsGcOOvm4R15DNqtWcqhYRYLKnbBNq8EBgJgT8YJTm0I8fgK/unywVN8dc64R/h2vdemHHWU
qYv15uit0mwgifUS1FR31jlzAQBgowJIiHSxBmvVmzi4V5VFm//fj33X0GGWwEeSp1x0nFpwNJcB
PgsxA59nTWp6R/jZZyYApLJZFcNMJHP/pgRPIDTia6My/M5e/aJ3vS+eGmNVL7nNk23c28Y1kH29
2xc94nDnbFu8F8VCIWMjOELm+cNOuPBLVTjh6lZkr5xvUfbpaxhUQCMNi42syidfDW2LAw6qbf8S
O7mnff/UT06bNM+ejZBT87vMtbjLKKTzI8FZNKZvvFiXiqrID6jp3w9loOPZyEC4aif7XVNdaa9y
RLJe8ncnZopZD0RA0NQXoGlJT/QRhj2b9YpAAFLRWhaZ6uyU40MPg5di6mIGAs4WVctpBrz+hke5
vvZlxNuVTrQIUYHa2MHJwfPzpipYUW8XTzx96qdH37cV0NN5y4F+1FvVkFgx4w5EiAMCFvO6L7aF
bimGwuGdEjkTFkIkjNDTb1VwIr5rYOCM/mhOv4lHz6EVz685QIg6H/pL5fcQDefo7IXa/3LPeO7y
X6nyrL30HfAcNJ++1VplCKlYI1fbHyvyIeMf5DXGDbedel0VuGX3FfcfP+BSatX5zshkN8beFMN7
cHFe8mnAPwLuAstaACfN9hzpuF2nqgLfy1mEUIIvszNLwz17b0j04Lx6apfN/z/3i9ry/IZvyHaE
KuE/ZqjuJ6UqrfzQwG8P14eS/7XvWFgoLHwVr5ROtDvLzdFzgWKHKiD10n4f3SoyXFf/VKmsHFt+
GrcM/UvuAXN/ok0hilM1EHeBszpw43mp29J5LDDiC9tNa4DYLap+oDtu9uJ2krBxj5GZuhB+RGdD
GgLAk+V3XmV+CXW/8gTMjwSmM1flxG5S8JJkPLPw4/YCyLMwrgNzYtAFYahEvqvOXuQlpH6cgp1d
+XWYb7JeM8iqkQE9a/QxUSTKzMml5MU9mIG372BgTB8KN64ks+F98Km5qXQTJQxam2f0YyU9B93s
CHMI6tBDQeWzDvnXMnbrx5Z4JUQoRHjRZz561CkxyT8/Z43roKXDnqxL2URKjZo7XVR4YESvoLYw
0NkYX+gqTdqHaPh7iSJ5Dtn6KgNMqLr50Rc12wPo+22iozDtt3oz7UuUoBLQYlhQxK3ZoH/Zyv0v
QVGbXcri2VuNDqntDFbsjpxLj62NBgJS/lbCVKD5i56sFndcQdWeEOnIjrtDmpvZ92qz+3hyBPsr
P67wb7Mw4ZvfdboH8/OM7sAkrqygYZBeIqJ3TlVww/tn5Jb7n1tQ2FUnS2vOscO1I6tRFlkQWR+i
k5yXBM/Qrueyf4ETJeFRGqxELW4NeEen0jMA4dQVyEmdH7tOVL5HQgGClyxArv6EUFmLy682DaOh
mauNA+vS7E3ANZTNEx51hFB6naHM50RwWAVtlDdissX7n62vIz6WDTW1nLI9AfZD7X9Q1XEXLIfV
OXQf3BOoxvtyIKD6OVsZICxzbG79BcE+ylYg+0Rk+Dt/PZg9t940+z3lKzFibbbWQYAKz3NdHmfR
vLvj+Fxtm3SechkgJqx9Cq4O77ZTExFwo7tQaMtxNKjkeqIR9Q4XZ3IWVC0RY42qwWv56FCcv06w
81/Cy255d8EhPOCFuDcvn1J+nhYI/VzSs29yCUpHggtXDXmOM6ZpYzcCrvLNPeLz1V9mLfdnsocr
cLWe/lWcccYYnbNr1QlvJ+6YGJ+nvZPhHZ3V3VBtcvk2NBGQrTh7YXKWgkExgNfFQRjgMdJWnzv1
rsC+jt7yg/T9Yhj6Te7Lt2FAsfP/ayuIH+FLjqkINKworyjoge7K/bMAsLM4XHCRtCzvQJUR6Qzg
RJXGxrdPiyti1AFcSazAiQaCAOklvsTcEOeJtdiAr1ZTi6+AUd3APFUN+WbJ2Am9GK6Q42URtOI6
OViS278FA1pWgD6O4fCuW0LRpZdiExtpmE3haPXVm+NIU1FfV3IkejSDMzHdlTBgOAnrFAd/EOfo
s12bVk++2io0jmGGYfi7ZopjhEgkPJhUEmsXj5fJtltYXEvKJzKXIiTiAaZrI+7+OwbQB71cLQHY
/3K4Ur4xpJhv65MHojcG0nTxmgl2enMlcLoSXw8CwbZXxicB2EHTzuuLItW4E5fZ50B3buzCO25o
QyduYafFxdbDEc9uMTrmf8JWitmZUnUIUEnrjyN3LSV4QYmNZa4dleVsEmlfIkhXxhHUlvrGe2hR
ULHrWhH1HDfeZvJXjISWHYzXvibzFyu0Vql/HQeuMYhlKKIChxwLE7maDP43dPhBL0saNjFu4XiB
yYaWBtKctFjoWwNTSPY+I+6IIpgalubVcUf1H5BjI9f4pgdsTlXfDS4NMImDot//fEJnsaDv38br
EmrnurKyLwwZ9J1WbHp3OhpkW5p8qdurD4y7mOXXJXZcnfRieYPrWNPaEBvElI/+OGDaCT0DwuBH
tGKu1nIG/8zJfCW/MU9bDtPxqsi5rR5As1qryvLUjahJ67q3oPqc/9vtuf+dCZKxdhdHjQH4hOWw
MRi5dIPHYpp4uncwiWVhD79Utzr/uzQacEzWkw1f3ykfyoVKZNm6fhnb18Pkg2POFHoN0C+nuMFC
Uze38bC9IyAmXIheRTJwRznGEVACi81+nFxTOBr+qSE8CoK1+y74MF+WwvB4Aj8527aw3VhX2G+Z
1XKfozBHS0Rxh3iFV9RPh9lM1lR2VkkhIWiqRblXtZv3JLjIwD4yO3y2BRCvnLwy2Lq0av7yAzif
OFIjPb9DNjeNIjZqKZr6yudXT7PiFC9c5mfphCCZKv0gUc5EC8NFolMtAZjP8vWq4AG3YTZpS1Jb
L99kuu5HUHPj2J817QO/lSjYUNp4hlsWZgMhhTPCQcfk5ufyWgEa0lUwc5jyHL0pFrgpDEXS5GW6
R3mn3pWn/paB4TxRweo4Uh++b+1jORwNpv5hJEIsVOCjuJEST61JbJ5MAqFCw3+sNvdaOwWXxfep
kWYMs49n5xFBT0RHPf1XGj/asykPMqvGC844imMoI8qGwnMwr1AN62+JKADsiFR92er5zDr7FTZE
cyvaQ7UOAN+EEdvizuldRpVSduM1tP3mtJY8JJqVCnEp4h7RsAw/92AJEb427w8RNg28l1OlLVKj
i7jo4OBaDvHB5anYeQ+FPz7VCFBQmicoF8kC0DNrSdMeZRTFaq9MzlSmoIWntBbCHMMpgKCongN5
TGoq9teFtFNp4UqCnGastNAjvCPyz2AiFSF0a8+BczPYXxhpLOADR02vuhF5ebvGl6cGICGDSSjM
dxREzYkgEIn08Jcvry+n3ir+RVDdLnwXLRPk/+euJC3QkX1bZ+U87yBBJwOlSeHt2p1SCq0EKUD1
ZRh9n/uZRBGdp0gFLHCGSjOozGNnGJyYqut36l7hX0bQ0dGQUzO66CJUUSvaA3DeoLXcKYGr7gQu
kE1qkxZD+oqvkYQYrJ5FIV/mtPtuStlvKev6j5kyFqDCDotLmhYCL3ZzQo33tNG0AOfHOehJH2D1
HKNG64z9LhuST4SzZbVzTZtlyR1KdP/nm/LhW7rUi69eK5iLwcX46IrpANDLS4nSGlxXBoPvTOBw
EjKO1MNjlSK3+KMmcIYM2pXyc1N6zcDdiENQkrdAcYkVi10zB/C+6O2OfH+lrlrX+WDmNkFjTVDT
zbeQbF8X9/x1wDLGbG0dpiu9FEDynjmD6H5QlqVO6vjWu5ioDndlwbb0MW6E5en2FoaSpLrTzoHz
dnCghs7ejDDYzGFJ2vzsZET/rrzjHaM/i7w6gGV0XDdYvWdWmlFAPpfohJKtUtIvtCISB6Txqr9R
0stc6x+LAJVdq7Gory4f0xxlij2M+uDa/ACB+JhbHMSfMS7BcbgjggC9Hm/ZfKyTgr35bOkjVZYI
mvWjkTp4LD6qodFJG5V7Bx3gQVnKGdWemvOa9d1c4rFxEpF7Ee6KZN4plSkdgwjZvx9tJ4miceak
JBcvi6zX5fRUpVRwEssJUr6z9qR78rnMFQ39qlm5FP0qjHFxqJtF4bKFn4EQCKR4xxdQUM1pBgGM
sURrM1g8O+zlW2ol+xctPtQBubJmIpnY2jH9aP6gXcoP49bbKjYDf8s7bn4AatjMOn1hmmpH9EXj
UgV44clgDoSkevoaA7lKBnwSV344oduMiqdjoDsNuVeR0psefqyUpSunsYjkCZKaxwIgwcS0nB5h
VD+bKKyg53WSG8tzbOcDNBriSZalWKH/YalvhEEDM3zhcQ/d1v11Meakvmvq6rAFzQhQUOLUjKvP
RsMKBb3rXj9G+zUzm2TvqNYE98EWICpEQS323eBhBUtYCebFe8EH6+WVOVDg2ueNiR1q26rI46kZ
UeJ0yiQTPMK7DA62YbIvMwFxqIo8es7NKi9eBzjfaIGEvCcrahlFpyETbVgh0+i4UPe5RloFumgT
vaTzUeuicXnlw1culbbOJvfnhJzH0Jv+CQChc1zdgrGkXIMrWvp5OwFCo0YHf4fXmEqJ4t4NYRAC
hiVq2CG5u1kZ8cdkNF2yQ97JdxH4nozmsTSSWFGqojO1+gfhjjRJOyjIer/yzNov7QOv94AC3obC
o91WYMjxDA7842hlS6J6Z5QaYCLgc0YVFOJ7YLFwqVv4by7zD2Mgc5WjniHTcRkvHmuz6ssE4CBd
RUafQUN8izsgvXcv3Va8+a6/CUbc0+4TLPbjezRKYW9zL/63mXpx07XKOv9cdfE+pihja9VNFag1
YWZGuRsfoOTy4Ok3IVyRHsWeqG+L+2KjEF0sW44jRESoQbwGvh1KhK+OMGywN5xMEyXO+yQmFk/I
Z6dUwrlOnLMOqcnZGZG8Whsqlb0tX+c+T7+8a/86px1ZvmISXrs0M1cr9aOOIZlmVaHBxIoBw1jy
3Ok91T5hfwWk6RLYmiByo5QFokq+iaSKiKJoNrjT4afZuWlIz8j9KgdhW5cf0y4oGLOdD4O7s/IH
2wFKAClyoo6KW5P2lBMLE/ipJbKeLHCenYOH9lh8vf2Ms6FkPaFbFMiGPUY7/22tLOgIscE6io4l
/NihxsFDoH7PjJ7AsZ+IF3dvw8VRa8RtVpOYlwwEik4RRv9y2BItfOVfKLCX9mpXrgLMYT8653a/
OQUGxVLPbJGhfU1Un08HEK/2j7zea/g5FklkVt+B6yO7uJyMTmicAho0SI98y0UpAL1zMfwgVJ67
53yK5R3L6CLeFNY/pa3qye6/O9XA0ng6uDkRqX5sUuP4Y5DCvlwbqYltFkf8q4NRQHWCZdqfnJHx
HbTze495UhK2ULaPbkklYrsLmk+R9unrHn8svWIO3ae+ukhj/oaDWEEnqsQhnWW9Hb7DPVX9+05K
vjxZf26OCMOFQFOxG2r86Du4TR6GiuNhMNbXMLs1sdXt852HLFv9jVIHupuvH3muWFcYDphhHcsa
ZmrGceTym84A3I15HbwVj8C00Ff2H8cvv71KivM4S05ZWGdes/0zmUKZzTCuQloqiN4z7onEhEHm
i5ML/ZuYGyzkdLSGN/a1gUGUYuOr6LwNpwcL60Qvu9JJNWxVTFHEWG12mKfJMnYQ4DWo25DMkJuO
IBft0LQIM496HRd4Q1VGydm1ufxEBOmXHuBzwP59GrO9groUEFNHqeqdMxBxoaKEYjD4mKhnh2ag
9ZW0r3pjZ/wPC9r10ZwI+9W1eoV9Td5NUiizzocVxAGYypz4RdczFZDS066itCuqgGP1wzx3mqwK
57KpsiE04nrG5mNMjtRJm48Opq9l7tHwr/xDcoVv2LqI6X7UIB+8alp7OD3oXnTJkZOuCetLpJ2j
wW4axYtlUcMLnpX/J8RmyEvdEaOqkMXDew8Vlcs6zACHknWlpM+eo1WSeEEXIn6Y7Ch9yRb+RfEg
U70ay9KFXytrWjNW91b4mvX3DXXM0j++i9Jk91q6Grs37oVOl1Ov0Ap196P8zX1sEIXOVLPS8Nxy
py+qVYTS+fGvwAt1vClDi6EE96S2okX3KRFhpEz1Rwiqi8aDjzlqdKmTIPNsFEvxYbvsoyB0+cdq
AJL8Hmh/Ph99hnZt+VhJ5m5q3PFoCilRIPJVSRePJDOPMcgLSG+558DD044PCUNVwPWXr59Clvv5
M2yMLzWVoahPw1HlFqNYbYDvtqRT2j3DDk6It9AtiVekmuBNLtAePhHFzh7eSygEx3OVTFHU+DsX
YFmqRFpUVE8H4NIvEtew8p7pUUSQ0lc7liUL7TUuVvhFS1fEIFLcSZatqhhzkYtzw1v0JOGFTgUj
5CBhYJN8qLxZ7v64ayHQAUN1nnCYe3StBg2aZETLrlb6H9WY69PAeos2e4hnc1/dpKkJG4fzPJNo
Mek8aHPk1d2BTQ9IhtSOnKMfkmwDDr6DNQ5X3je7qagR6V+yj5t3YbpSlLDcDTJgaPYdO24qs5KL
PSMAaCtk1D/GYe4XhDqkDLVi3sPwLJD0l1qKCBzPyHxTswywUjKOS3tZy5klvN0Oo6Go7oAoAQub
2gf43EwqiaqY111o4bH25pSh6E0JGHhcHZOHdO+5uew8wIKnH2Ynoc87nXYQ7lvU0IBe9StmxO1t
Sqc3mAM0uXXrw9nDCbM+LNjBcFZCcXePd7ZLu69UlPfJqTKFo4Jze3ePbtDfFP5v6379dQrPFlTh
/4X7WFNFNcViIViK5MXNVV8+hsY/2yuCH0+i3Bbm2A8A1BYyIseCkGVzgiviTAvvi46m/Sxe9KJY
wAsp0oaNJJ/BO2zLD1qQw+RRhp0IcwjyelI8A4/CVZV/0T+bN4yCo0NqN4POybksrE/GVaIvqbAn
COycqoZVmXsuugfwdX36BozoVj/EmfBTQErzrYJ7Iqd3pmTv/+8Z3VGPmG25OY/mdSGeg1rtspty
RRhipZXf+usZ0ndkmRtNfiE9bGivrvkZY5ZvxANqWfBsddHPgeeq2g57liwTmFZYxrxuG3bAIPWS
1B8WyQ/MKws16iXM217DS+Tn4Ip8q7cXLzNAOD/jrGiwZD885wPhwgur5DFdjlEjYScCCIpmEJFW
orKrKz2wCF8zB/RE4Zb/OgA6hGWzdzUWseMaRlwV7J0GCu3bwWSYQ1g1HCGswaiicv5Nc4LjRpgF
BZKOpkR3Kh/D1Vd9snOsI1YFh9qBjWa5hGALZuFHDx519Je2ECo/NvF0L8dX9Di1ncQS2/kN92oe
CpHD+s4gT/top609VbxIIRlOzhU7gHjy8dgrEbDCtJrXxrQ49GAXABmJDZQVLUGLTjev13fCFcXq
7SUGKoF2wqpamldyjJDICCMGf8rJT05herYeqI1m8MDpQG5qBnZ1JlXh0WbcwXlY8Jrt4TdmAtUa
H6SajbRg10eIs5WNQAZioHeJMJhmzGTKaALBnSwMbkEK9QgMNX4amml6Xthxp3GxbRuILhXk168R
QcA+TLLzGW6TIN6tic3GTjeHG35l+utfJcsNO5bXdn3i4vnGeEsfEKQ8qKo5wxbd6MlNFWuj6Rgm
wFmeIOf3qJ9vti8UW9RuK14fsDGIPJGyornXR6e5FzSkWGBKarZeojjg/svS5THte+dW52Bruw9d
zpTefleo9fiQQGS0dnuvOoWFlJrY7DtZmpfVTMY/S+I5h05iLzOxL+YwLzbuu9MeEKj/s1jXKRWZ
57iOUtMqAG9TevJ/NN6ZhqVwUOd9bC+4Qjg+PdwQv61uR7r9V5V12F+pQnHhcBz2EpWSxPDUY1wx
fYGLyrMGOV6sKdW3OPVSAATPnqR2dPLnT0FJafHEs9FRf7HowrLmVJ2YmRlvQmhVNTBS3MsG+uEd
87GAPtcg04L0Zha4N7Hoj9PFMZ4Lghs2Pt2NwEfyDP8vU0A3QDaLKRyBvgutKbwqQpqIVkO/7gmY
u/u7lVsyRUnXmzG1uT3YJ6CR31QPHYq4lUkstuLmK6fRYgVMPbFyQYLorKxOHksdecMBkyAs/dZ+
IOqICgoCjhRk+2PgSehfOnF0QhdJyEnPi8vEb5e4XN9pHx2U7157tSWwkl7QhyghRCi/Scf/vzuC
dq0v7OyjJU4DoyRUhZLJhjTC47dhtiG47sJd0zrkXcg0Jbqnwnqr6JNfDeEAdyQOxGn8HMPkd+KW
CwQ7q52tkKjW5NI05B+D0962qNxuBof3R2/Rs3ozTAL4IM0Ry7pW34hWvZEos0CDi0pS89ITByjF
b8kJyXo6m9m3u3YHUU6HnQH8A9+zsK0Wg7UXVkmHRiHTHzSCBLHSr9X8CYfZRUy8Af+nXy6e520z
bAi8g4Pin56m/B56Qj1QMWVeXGzeiL6xTo/6jut9nq9eISumnN8WyJjLMSn2ThSznS9i+qXoxqxx
n71vuw+rtu80Y0dkJSouVXo6h6xpO60wBJPkgeElv+mhJr9VyiHvUGHKjNxBcWDpHVztjL2mxMB3
pOALev5Cl3rTOahWnDa5iIDf0FqE5jsrOMFT0Ef8aLYJA13UnPud2x1GCxByaoT0EN8jkjLhqkmV
qrzAh5znRFXi6GV5LI7mI4P6eRQuzve01pUJsQMIPTaI2hKelCEl/w5LTL5aMamGIvKw/woQJT/R
mSvnU/au4MP5vxRpmoDnJUu1sz9+qCYPMTr+CES8uIQLEa5XFMt3vgAyt2bZbfSLzTqW9bKw1Kby
wy8Mll6VjCNgVqwHp39fArONm2xg7A8XlrU/u0xnThxOek4nkdN0xfZoLQVouJlUV2qDQbmhfTV9
ZGtJFZfqPmhbnHa9QtmMRIe3R5BRCSCd6tilJ6d28OPRoJAZd2Jg2q1Xtzu091e3uA//bI8IMJoK
DTYHyHuyIgX4lNJnZuX30eQZuVTG/GkCx0YXIY/+L0Gy63xyYa/tTNBZoL+OAglDFPk4UayN6GFm
nrC9MCY3CqVwjRRWypDg4BA1C3jv2Vc194GO2T5OIe5UXlUdl2gNmxUbS/WTG525wbdC3qS/BIiN
yNNVGu96Dj2mQNzoTMCOwWDmJ9W5F+JnEAPpc+4z7AQGPEodhhT5TH4uopGcmzUFSUxQtR+LwVo8
bj0tTLTmUJ53zCLRbVdzC+No+LG97YIpMLfo5ueayYsC55tYoSSxi+Ew3/Dz6aMSCGilK7sF/cwj
7A7+np/F2TuSf0ZKfTUtI+++El1Ub/biNr1cdDavAVYrSGYLNPqWZcfqRvgDiBbfmkRDR1Uv63kr
08NbGKlO4qtBDcX4gd3UFQ7e4IPHL/n07iAdb/25uEUq5fBzRBoMnDosQawhwjy8u7wFckNsXvEn
A4w17MhdXrQUcLoveZ8y6Un3r6WIFknCjEB5Azk/xfbgl8XYjsH1tiGCIZiYLIOVc9wo45EdgNOl
SjBPkREGmOhQQfX52gENKDgCzB7PNXCnrwk3ldBjnmZcF/tm6V8SnbX/LhvnY9hPnXX0IcYEX6tE
JzT/O6SwUI8kMwwwVfxakQQ/2PSz3yQtIsgsnPlCx53XpWaUxpCaz1MPfNxNnqTePk6vvTMepciJ
gjlvY02DgBDOmPqoATwy3GSb9ku8WiNpB+9AZYXnjtJ/BXam97iJlAv93udmMg9c6/S0IRvSX/PM
j+uHGFTQp4SVbfNjzXHjA4U7ywekSYFJ6T44vul/GkPxKAUu+8i+D4U6qlITYca72ueZn/CBtIOo
h4kAk7L4K8GvMmVUFBEwoLnEwmzwL0ZaHYyaWEnUCVEpbSdtWe7GBQLt4DkC+GLZgTizlu9VHowk
I2+eIcrE81V/YDK57eUPP3sKGiiddDg3swxzkSAFKBGOZAZwUCpePK4fc0ot78vfVe3tSyeYMre6
xge2z62xXVpQTzvj5TdlFEG8MShCrzHArtDH5pGKRAp+Ta5WBb2DyA6ObJ3CyWYNthXJMAu6kxGU
/YTVHtRFmVAwDtBUDH0IwXva51SGji+Ry13FrZMXoGdT8pTfMLUzFMSu1Il3+yFIqKrjEgrfHL4q
muCKwp/3oj/0NqHQc7Fs5nv0HLxvux8wjpZOXSULOq7qMNz5/SMvjZS/7BNzw/VOHiCQzbPtAB9x
Bm+jrAavn55pXS8HxsxFpnqfTPH3/U40JiMIJQ9STHu6USdh8X8o/Bt0zUM8YrBQGZNGQGnKhj5k
+mz8XzY6B9gDeBE0y+Rk/1i18FIGD8jRMgAH2W5/eiCs9FFq8zKmSHsYo9NbDmwW9elyGR8bbv/N
BGP/ulSz/6spMeL4nCpyDxeAYGK1h4m9qUflV+h5tvwBuqbLnJIucrjt8zs7AXpd4RLeQI4vYUU7
iEOVQre5rNGdgv7AOxPrLsELHv2ZLIU/tzlzbb6NnBPNWu4n1rGAov96flSTzng8z6DcbT09yUcF
C+NyLtfGYDACA7v2VhFoIMcCX8m/sW2qJ1pt4tfh5cX8E1e8hdzfnm5ikY4XLoFrGPW2NH/7yPx6
XRyPqET0YEMBoj4tsejvgU13XPLbydiGTHqEj2h4mOMeKkqz4JRxUyxJaG9essBR0/BJiE8CFXO4
nxUTL2erISmAsKQhrLNuwdtpTF5KhjZVfMIEi649hGyQX7gBBQTH+rpxZ7bTIs9oyOPOFtWRDim0
6VPr3x1Y8WzNxnFyTBlqkFoTzT0Ks3LR40uvQnXanx8Vml5NZd6xt4qxo0WcXSTyA5RXfcSS3akH
aatpyoVIsM6ZmhoFlq78bLa+VCthrIl7n/sO+Zy2y6VlYR8VhcN6aQSmc13okGlx8Cvli+BL5E6R
Um8bHuhohUgSrqMpco4X7PPkod1CLlOgQkATNXJ//y3WNh7M35sooF3t2erG9U6YGSZy/izczNje
PblEx+IPRpdb9/tAzYSdSoWwPNPjaS9aOHWxU3yU8KHhZscs89407L1gWpk96TK0QYcPUlYPN7fW
nhla8bZDwGI0LNGSdha6jb18FTMF0y0a19wJ3X8Mqg4tIcK3ez3p1AjQ3TorOFoWuCor/Y3Z8rcN
j0xyL8VQHIjcJHViK3OfFm7zXau5jsWvkkZgEZ3rEK+7R2HkKSeTlSZXeDNFgQRTAmO6j/h4MUyr
UlfmhO6GWdPeKbbYr1P1uHrV0zII8D61F+42Ey9HT+S6tuaFKgU81YAk4ibrB8bkXOzzGcgqidDY
qITrehS7+uHLI9TUGrynUGKgrzBR439MFtZZ36ttQjjFLW4Uzhaz05a4l2L1aUFABm0SLrVu5mCf
2fk+xwJk2mbztZDR6JID+kp5HiEf8XTmuckJ0mnRWywP7tBDEqCMm68PGdoJMvfFcjsUmP7C/jhx
8VV0n2d6M5cpAlgTRcrGPcGPxPUuyFsFUtiUdZyOspoPSHexDj8qx6ZQbggJwY0w/6Mh3F4qNPdQ
xiJfjfyibseY8Vt0+6xfx8aAf7Q6sw/SG18Z5Tg89RGjYAnBkRPOhJUu8b29gImj2eTuZGbVd1Di
zBhacX8ROMI8zQNf1Siw+bWEVYgz3W3ujcMWIHA5qIHxr6Y4hl1r8hBJbmkcU7j50V2sgnH5xbRK
HZ5s6rpx3Zc+SaA5TeOO7iRhGd5CYe5p4ONqHlBS2bqPMyhckGzJa78MOHg5EdVHp9yaizCrKBMZ
FuwvVM3kEOa1vVG49qJDb1rvaEstc3ranaly6xyp15sUel4S2g1I+k2DkCFXhmHhOTEOZ+2a4jgU
imYW42FsM3BM2HwCIj4HLkowT++bKJNp+G11Iujv1TFMTqIdn8zMeR+LaVS4NF71Dw2/zhRN3ovi
SkwAdrOOtz0vvROh+ujMa2hwdpp93dqBA9G766DshmL8R61n8q90EkSMa5HR6yAXQdBeEGhyBxVY
Fb8Qs4xQkDOmvI+IXFe3+QNT5mxV1dlnXJcQtvS8PshQLi4YwY8HhOSJI38MmPihIzP5UNTOnt1V
HCrGRzBJr4fAckjO+MQKjSdm8IuuIjDygaw+3hvltpPYt+djWniXIsSpR++AMC9LUXfq/w+oYgVj
m/dK8SD29xEnbLX20xgC7xGFD9uO7AbfghVxv14D9GZXzF3TNBiepFReAoutnWLna/qpgw4zEbm9
kpY34oebwUcZ3fpKWfbXIy/SmuyF6XlKUZh3moAQvpJMZgkejpx+HNGO59uKWdK5kxW0GCN5ri7m
legay4Vdo/6As8RJadGCvY5j7L6/WxmdQqyW6OHcfSrX1Bjs9uek3yfzhCcHd8DArhMpCvKSbR+y
xuIosdv0m7enMklUDKElA4n7DxaoWsidP+qpMA+l0eeSYem+ZXGbf7hIACgqzBRh42m2EfmOz9kO
KMBtz2X+aFUgKK1lukatV3qydz8wt3Vg+Bh18wqqQSE7PwRCtJe7+RKXS1yJyZAyrdANdMjmA++2
Ej7Q6qF/As7Z2KDnPQazX79T1oshl/fYCTLtOVMLkrAsA8Qr6ymLAqzRdAqzruvjKpFoSDbfRoYz
5soZr3z89tlj2q/O+KORUNmuiwmAgajkPAlmny/B60dCqjP2BSo0NRP72WAgKEmVJEGKohLdreDv
Jeb5Zxx5lbYBCqmEQbzlHbINO/juh4aflCf6QpRRHGPLo8ods+iKI7A3ghjbug5alS7UeBlrdt+e
yCbVXsqv/MYinRnJXBZf+c5cEMZ2ciRVmpOZ1hVTz2n6Xm9Q49u43JPhT1mnF+kyC0IR2y/R2Mzd
jYeKPn8yhsjp+yCYss3EBQbaeH9jXjmA2YlKHUdc9+zl/SiYaHi9bQ8aytJiNHA1bKCj+/n+xJMB
YTv/kwNFS9udhxaGMqutB/wTxZblPKXhW9c/svTZFHoz5zy4ogTBnPgzvSt5jzrQyyEnUpCkZF/e
58ycifLwOSyf2ls6qWMBRIqT2E6mvRwPbyTekba+gDvCKjBDZHwU36glsihOFsUfeHPZzjsWx/vc
Rj1at19oAndX8P2ETs8ihbyhCqx0suaqXS1r50LLMHxiLbG+uqlxBxHZ9dKGNZ0RRKXOYvlEov/N
Y2IeWfDSf3Rj4zNvdma3dS+KbyP5mRv27Cn6KvDP5NK1hDHIOjgfGmOFME/FNboNuZ4hV08SFSnw
Krn9+GcH+memt6AY+JxJ/IBYAqPHFxfcsQEwzAWI96/c2yiwp1lknO2oFHmZddvgUjVs4+UKxgsY
oxHLwxMZ7sLvGlhzg+yljtssVm48Q8EaZ4W4SiZv/sk/NRhBjUUSqIZuH34rzJdu6cQmNwN5zzie
4Abq3LGG0xSmYjsZo5g78vnXX2qOldmo460moCFlhvjcaXaOp3H/yhO1I49L0tJz3bjc1S3DDKBg
qgNRRUZahUqmlr6sHBzxh8lLlvwL6JfD8jzdYDxFLkbJwmWpk1lpSd4ZUJ3cEO+UdC2y/yHKGUQc
jrArkmfBxyMWutyrrhDMyKp7sdrUrwDVbxYV2aj8JRF29FlvO4xDRHFtcilE485PtRtVTYXI0nhR
ovXOhyY264Tl9d95TqlxxtJfZmQ9rxJvG4jruZhWEAK2xEMgap3ZCBBQgRQtn2Az0nURiiNTGUkS
lNXqK/4/5Cv1nnDDFO7HaQZn4SXl1YRs7eVCj2V6klGmnymZOVzkd2jjMFjtUzZGGgpoAmPEYdUN
9eS2mnTavPunJap8z+pvsfNsG3v0aMachLFb+BL5p3tVUn9DOOw5OaOI1sHlsp2vWjpR02suXkFJ
qpvL8r81RUCuo7StNIJHxpVOlMFZ9eSvqBtRZ9o9AFWGUIr5uuraUlr9fO2YtOYLivld4//Oam9m
fE9uLGaM+NqAvbb3Qygw4K6DzqxHV5/q/FblZhHU2f9BEm66nvjvw0yYTXFc95Y0LGq4asTDbsE6
agFUcm0Uz2O5i9gy7YkZzTLDsKknn5eUcplXpLnLpOwuGUlsQPqCnKuLdANG71mMlHMJc+BxyfOg
ar+TG+bq/Ms9wSGckBOsg/2m8R8Rp+ogiibKII/FzPcz8BRpnFEKJFG0eCB1bGId/H2ky33OvFcD
e4ymCyiTUYrxwzM7mwkwQHhgvVEFSP+t7jvRfmELzQ8RGE4vKwUuUw9EYSZR0cuN9+xKItrqW/X0
5GFgcAm0JHyD0pLtE8/5cc2DGYDx8Ii2cRnvIXKFf66ex3xrRX4GNYbp+qU+jRqMj/EtGydooP/4
xbn62kLNskKq1z+clK5hwGDjum15cmh4tS/cuFBiiFTtWVC0fSsZ30ftENzQqxd0CuKkGjdf8w9V
S+w4fUK45/Htgu5d3v+jJujzo5nd2HMkUR9a3V2aRgFeeud4gzdisqOHnRXAhGVbQyBpTv8pa/gu
q2X1bH/u57lLbsHWcDTmftcqak3OKt9hcScwznyszU5QlGrfEk0Hh2kJhC9CtX3gWOEJRQfLsufS
UdJsNy96CMB+S4CL7IcMXJKf4M0CarzkJd9yetZIDzdCC27HcQw1kqAhFvaX6itg+dY2hhQN0c3M
Sgsz2gCTEebsKPGBhbLjEsrLLiUGBsYSB48xGts/vj9psqc0O6mGr12kIqPWfADzDOeOmQQQTCiE
YVRYcE/He8GqqAp3+pDQs0Se1jjjQhpzbnRFBbpw9vlchuay4KcR7kcAUUeh1+J1ULTHUqInrbEC
lkXaoUXPc/KDfta5T2dHT93B9mC2z6Al/hEeFVKc7zBEEsq+MihRgwd60PM5+jJHOPdSYfC2nqpq
TFp9i29Yjs3Nr498NO/0u0RQvRQXkkrzROvJgMDRS76H6hCMRUYtiBHBygUzQLqHVRpv5DmE/fB6
M6brK1llnZ7PRhFjj0wWaTt8CWXA0FWDRcf5wwV9uB7JHMOF09ctNevR+UtEDmC21msgOcqyGuaJ
dWVys5CGqqEZoDtWZxg8feQO6OycUPlIviZk0VvIvbRHw2oclh8MZ7olDWDQ0f8n+WlJAPpDBxRy
JIOlDt0ugEKKi4WIx+vmBOrzrcLYNalXRRDh5mRVvARzlzyihd+iqfVo9tm56AMvWNSfVu9RQ9XQ
UlX41M7+tDBJwF77NcXzCzlLZkCQoGCjouwNqy1eC9G6rY45K62uRfP45SA/AvfQ5cz8kX0mhrw7
1ZNLp/eqQxC+5nrUOaS0FOd60u+MWkMBXB9vsyIzNrEDyOPS/HFSuwdkzWNvCq4M6db73s2WoeZr
Ime4QLfj8KaoU/eYIhFHKJdvkqn3vgAhv3oyO+59kaoKkiKVrjuJtAzD/yeRUoi4Swk7rH2CHeHa
JyDYeoBQ4Iqf0E+0WxrOCtuY4osNaNPfN9V5siIl9Ev6r/4CB5SvZXm93O+Ynq2WP9DnAoon0ZEJ
kyd7YczMBYEBicBigRhIxC1nQoFWKMYrqg6XXxIaXZ266u2t4nA6Q+cd75segfH9YRDaGzOdXcu9
EQ35Horh/EhWQtJ5WTsCzsqqpXmhy68eTjkjIpJM53Z2klwyeMfE+fBoFALgC8eAHSjOu5Fowt1C
YHX0Mbyblz2NveAt/EdFm5Mj9CREPRNzWLe934XRqFblhNg1JfpUx/8+nB+TwFRJRwcBgN7gFTsK
ZVJeEUbXPlhYJTk2eEp9pSyZ6ZMqxy+03M6Qkb4fMAG+Lpg3eq2Q378CzPn9Bx+cjzElQyUTB+r+
AJe/+1R+wcogoTtUvKOR2f8wdXgtgyx7M46cj3TNVcvmqVuKzxVe+3KY3Fj0jsDDvnLTknSz46r3
k3uYkWuT5yoWwo48TiSF2O4nxK5ndWmCh2j4TCTN3aOPqUmdnmruQIqW7+VgiICE7HyB8TZXyeFt
QWcQnQ+nHCPL5rLO3CFclWhhG40iibcZKazae+xoJkBixNOSH6ObyH2I+YfQPul9sIjoILYLvu4C
dYKOga7GGSlSayVEnt+11zlk0OosoWshq1CgM3qwiMVWiLxEnmKOSeKlkWRqGR9gVVtlvI+IP69z
YvNmltb17NnbubVWTlOiKAXc6rharK6IK1dWWh41WyDwcDJdMeNnw1EQvsuzxMT4AMUPOzG887zU
C5EspVoWXVI1h+QBCmvUkm7alKOiCH+mlPtVtxwHjbBvT9mQ7AKl/2oOP4/aOCyoaDZIzE/Q4jtT
idzMxbG+5dYxA7k0Z5f/Qx8HCovE0cCM3LZ1tSKf5s7uegXYSLFUATHRb7XLq2F793UU4Ynjq+gx
Sx+g/yNJ1eaV9D0PlZsyR1khFehmMKyOJ4B2uARxgUBkjMggVuTRzEQeaxtIq/D3utfI3prktWpw
XeaHUzig3I4LDAC3JEVYbhxk/BgTFeZNA5zEkh0I/dmucEXr33s1nmM+lagvJs8eS8j7dTeAMrkQ
8IP4rKe2gIGsIhy+Rb8Wj2U7ut98ouchfQ96PHQMiVwbpJ0TODWVFRLJ+8liW//81+X8GCp3ziYE
4/+7BcvIxpxD6ClaMXrA33NKn07/stwPY7m293yUuGYDonmHAkuEBT8M3hx/pMrfLH6mv3UJqS6y
9PpgD73eO4Uo8tri70s3HW83NpZp4wPYKyjG/sELV+60ZHH62cLmh2Jn2EQ54NAyunblsIAXyGvp
QgLUiCqJabAHFjbXLUB4IqRuMwLor/aJ0v7u9fXDkMyjsMMCxprSScSNFBKDDTPei5zUOs5AZ63c
1GT4tENnOimu8pAk94NqYDrOo7u5y+IftkVVOhNbzUAXbW7Lx8PHrvJ6V/Pn21ArEI4QKKZwNj9O
D6hQhufx4cqCBHaZewKHJRuoI6Oaj9/+WSJDChCt7vwbuVhimiQagcf/tOhdixluaUPYaXCvXBQD
ya8DUo5jwpIbASbIYhxXtjr4rtDsdZvIj+CMjupMT53okYB22WscOLsJ4QpLV1r/as7GsFmim0nu
QKCQ5BNz+rPJsu+kLva4ij/ljVt8XGaUViTghs7QuSe3KdkSIyfxs1nab/8eER/0aR5p1DV/lJDF
9V1v7e/nds6v+a7kijr/YSz+EQWezzQaLAfZCQSUc/I2bJP6EnIlwD75R1jIJ+/QpVHbqbk/9CZr
uDN1mdnUIgW0qB64tp1jgjrCObouXpmW45KvDLHuxnOtNp3W+m+k3iEUudZ/BV1vAVZjq6B1ms+h
7RiUo8GxO2NK5AUONISvhWC+gDpJasP0myri6Kl/A8mAOGkKRvrr7ac9sbNjcVEXRxoU2jLmLbNk
CxuBsKmgkwbD7QH7gP+xohQ0Ia0446tNwYrJvPeueXTKQSqSOPAznfB8V92ep1h0Awo2+yI0sjZC
KJJJO83vUZNR2UzqWI14rkC08vc0sQgTs07YVN6ogbGFRLk5MfL0zEPl9bSc/T0T4MgXdjxfUY1n
o/dpzN5tJltrItDk8dR74pl7Z8B7E6N/5LZAj0za9k+5QRH7Yal86SIWyHfiZtIASiHZNJ1EYQO+
Wkf/kj8q9+/okW1VrWwViaHpxOfRxiQyERy3OVvSfWO9gI3SBnpK935rJg7ngLaMocHj9kWo1v73
Sx6PjBc2bvxXt0pDNvGwZ836hRTMgFZ76p8ediHItX3CIsMll34I2aN9Psk6YeDFG1LYYWpFseRe
Rgd9S15hhNwxWzG9aKlvAXeyfC7BdiPcYL/va5jnKJw/uhA0d0vZSDZIfLY8aYDjEn1VVW5ZjtgQ
fBEjL40zBR4yU6qztKUgyWGvF/UWFxBk1L8HtxV33upwB737QWpbVjcong8lhS+52LaxchGlEel6
QsLdxmbKLFwMFRQqsTAMB/TWvmXdbLyCTYJU1AhR42OwG7w0qqNlhQeVyLmDBEQuqjJDkqRme975
f+rLSboiooOrXcqcLcNmYLNnwRn7uYOV+uK8ZMX5pvS+SgC+ekXj8XGIwi8FjCyRq0MGNavjU0iW
u9r9qmPzUAdJXTa8So1LZ+/aZV6JbRTF7hJ2Bzbrm1Kn/+/NYAWEYaxn6zgWG6Fcjk06PCjr2YAM
Hc+waUMjjxmob9dwvJdEn5+gDEqL5myNcwkXAwbZc8J/vwtJRTIPqJriESBZUM37EXGtJRjlV34E
ipMyvfRSeYdXfBLfSueUlo5p3USUE+fPuiCGCfzjbFPfjVmZiAuJa23Pl+nSUyBhBswxDaugSxvE
uDV+TiaNflmTDu60fVDD/3jx3kUqspPBSbYbYs46gsadLXYPFFdT30ajyGhtqTIC0+OxZ5MbonJv
We4+mE3+SrJGyKK/d6aYydP/6ojHwq12KoDPJeW6ij6s9lA9dLVp531WhcbVxauCWyCF8uWcaB6v
jH0tUOXXCTW2+3GR5yhjvewI4UE4PvZSAZ0LjJYaZeq61h3zbLOdIi2skCHg/hWNYc2YyTis6M3W
4eZvARNnkSzV5lz9Ds4IJyEJvxQeRss5P2YpM8ZUNBoiiH9iKgmqUYAi12NYuzOVMgNNH/YzmwfT
yeLxhTmKsGRkzo+QpAA2WzfCTdTI2rPIipNZ1mILByVC4x8qvOlKIDb4C2ttt87PenaDF9+yWRAV
B5sIafBPr8Or9lMhpTuSsokEcd1Qtbm6HvCikaBSQXLR1OoULkzdWYphu/6s6Ds6UHMgfCYbp5S1
PEdhbB3f4BhlD9Qftvvi5Kh5ghH3uMzPnju5nZSEAzV1k+qlwk0Vb8rhSDuAX0ImJXmraMgdBneT
VqcJC6Ts6Q9cOIcMnmQVVqsB08wK2SLzQr1lQf9//mbLQyjmQg03JBo6u7HV4Rqxilw8DifSjbQg
FlS5wAZ8sCXUBHLNO7c2Ld0h9uKIOmzIFg9xhM0OPnXc32Sv8YjFFYlXVoblePwtsoe/plSuiQ2G
b8vyHrdW8MjO8QNyX+QxGqR2hNNvNtZUA5LQ9LVphY8xn3FQAs0Q65LL7q7daw9/KepLPbub5JfS
cHim2htvwKirz4R3RGdIi8kHorvseohUVPuYmLsm/FRMjSAGhVB3xTL3fySQBoQGdZ9iMhAHmevL
5pSa+AKrXC5RkEk3fohRog7wSvvaRjOSQQD2PPbLUMTs/5ByPC6UyWZ4T/oIw3EFPkCCdlIaFJ1o
LcF37k4mKWBvfnGoXs+RXkzxZEpgGwmFkTeDAMk1hPERusi5tWpjO07sR5suD2mN2ieHSuoK6hVy
aUolFfYXZ8efY2TnpWqtDGr9rlE27s7hCZ3BaY4WJ+8h5UgaXWJI1kZ/rCqF1JBto+7VDZxSHjyP
/RcdNKbIs//hp43bca8fEOFeeo9EX/K0bqOICQ2Rjtd6S0QqFgeEKxMgRWiw2G2lHeamsHDujwNY
PzHPDwMdoagDK1bnavQwRuA9LA7ERdW0/qMRmxCqKMroUKZ2OCbWRstR+aZHKMQ19VNiKFZpg1dh
+8qA+BxHHJtEa42W9/gbs1yEdMQYQIpqiaeIfRiio66a579u55v9j0apGUTMFfaTNgjlN3gsi3Qh
MaozgOmfMt9jkHgMkvNDAdSRtuk0jBCqmS64E1PVLwF1WDOA524L0+bon1J/OcxJEifIeaiWA611
9NVhd08Q8Flf8gtx98Qu7do0fsnWQCrUO56pmoM10IOKflRVgn6IFPeCw/PBQejWfXvMOyOP4fCX
51SO9DGFukx7xGWqIeunvxwFHb0FineTOM/RYXsi2gk6k6ipOVHyZiyGQHuFAoqeLPosGXb2Eke0
I7o4OWJM1P1xVIq2d998E6c0O5XwUSibwEIlSa0kLzbV16Sd4Ay1kO8kaFVVxZsysx73AqmoMzym
bptSx6nBekfEUv+KxyWVXLHT6d6+z73XnxSCmbQOK09djcnPBLfTwxoZAgc+hUzTmKNzmyptr9z9
I8V0aILO5DQD2s/TepofCbbsdy2l8AoFgIls5rteG5b0dLVGTaxTcUN5N6slY+m+oFOUYUQi6k/q
ncu2bzRhJQcL8bA0CcxHkCDEFQda9QAIc+p/8xcwurrKZ/8jM2mAi/lZ9bgduPMkZSRrF8nzTwSE
l1CoaqL424r+3De0OZeTAWqDfIaIcZSFoc9Sv1ovxMXoz7cPsn8r5WMVj5e/AqMhk4g3u35FXjw7
CXdgJtBtx+YSo3funbXMNze3dlMpDxcctgZr4I/piHPOfd7UleNiYI5m7hvb8/NjFJF086AOqQ51
SMQd+6d0tor/jJ33KYU3/SrcHGLMgf/2ZSGbTtCS2sSCeRddsIJrfI+iJ1NgZCNyb7BUfsbX/PHM
yRkjpb0HA34eozOQyO5dseanBZIFvQq84PRy/PMyzfWhHwOZPzScfWjxjQIe7WQnzA7jHz2txiQs
ZmzVSQ9eKgbTvtsI7kjnrsUaUpYFfF2SQ/F6eYssEYZ1WbLe+LHPY6tonWCa3FbFa+rKuu8g/9Tw
uV6djc2OqrqkRAti/Kpj4/Yux09WMfixfFIg57UlhuAYcQoZJICd1E5vC58m+dDzIvieDiMMAMeK
e/Bacy/909bcQxAOJi+AU8kwUtzxYkeycYn3pC03qKVpcwMM1SLI9+BVWECPcO4u5eYAQAY5fSBB
Uv3Wtw22wgqGPqzJ2XnMsxMp4fRfUhiHQoq3EUyIzWB0gqKMOvhbkQghl8rjRdWF6jBRePgG7hEZ
c4r0VvfriUqUVUbd17kKGEXDfXfboOSBN6naeXbtP/hE/N1Cech6nSv77j1q3Spu7j86YZlqg296
0xIi03gGAJQ54fL1+gVxNZMGum773C+fW5lKVUlU1BqbLZbh2RS9DXOY7R3dNlUsARwXif1rf2/T
tVakkP+ui89a0URCDSTbp9NbwP+NLBxn6aOHK7YXt1dzF3OkbfVdeRHrs4D9vffS0EnDTrSxBeaa
lzzbacFsnUn/DIUEXykpLvVFxEPydbGaZP5ibiAf4a/o6da4Ssiv+eacYo6Xdo0bk8GPZYmh2AOS
77OCDxx1Sum5ZGLPZnC3IPvmnmJhmbDU0LYWUcfnhHY6+ebZI71PPjieqSw1jh7YZ/k56Z4BRe1r
/K16vLWmNCqGFe7/Zl7AJMRVRQKfN6Fxi64bxn5lUoZGqvHe7/9QUK9edXjBOQKWcW639vl/sgC+
+OzWzw++Ru1DL3qjUAMEFyczI38UdnIfRy3r85D636YmneNM/FUUHnKw4CkBDgvA2PQwMZ0pE7Up
n61qt+sEaWqgUa3nymZeWq9dWpAeBypIToBdxYMVGITKYYMDNtG13CJKT6ClN7gCtkBP8zGWaxMl
K4dzd/1Ts3N2pjeIp/1mWOROXO4wKYr+zFjFB5GwBe+m82lCkABBk1LBCt013r6tAxVa/qAJZbxi
/xYWh/qlCnGt7FpeXIKfMp6ZgauoyQ/zl1oaR2bOlFIERMWqIhYi6CjCQdRIi8FoEMxLsLgO9/sO
b9szmHbZPTcDVtwnCV1ok2sShr5f5CHd+gSg9cNOL8F1XlGXPHunLn0pSmhdJ3JZa2nrHXhikUjT
gLhMIAdO0tHx0e9lPtHVZSVOjVxT1RWwoxSTOJrVr3ME5tbEGdx+K5xf/NtSdtC/pPKofrJ9IWk+
rCkUyDuAOHMFjf4rNji9gbX+hJLtlXuA7XGZxpDISLY97VEuXRKpmC5dWg8SbfgWc0J3Sahhq6jX
96OufhfY+Rqv5xdloFdQYZx34SmX95nFdLR4RBJ/OAdj6jZY1DmoAlu6YSAF8GsOtgC+4zbuUwSy
KHKMTo3/3anbFhmGPm8GcGflppaPGVsJVQALdIf12BcaELqj334R3US0chuE1mQjbHgRg6W7aJ7j
scINHde0tUemV5rf7rLTbE65H8kcsZqGl+z/5bvIohFP8I+RxnF0H9UHM2QL5E0UuUgZS4pfx4gb
CdvEr3JDbOyYyHAjZfIVEVp4gUPdOAViBJ5kpzPsTKxRM7M9poz/5B++JxfvFu79Yoz7oMD1v0IY
of4zQMtBgxnIhnCNqxOxMd1GGdWEB/9mu/uJJHr1jXJ71mLMUHYNn93HAE383RnfkF2bGkmMAqXq
UPoz7j+veNHK2V1m1yyFjjirwc2KTheuEi/fg3OdPyymWgkD+yOwFdDE6PxBvQTgdJ2Ci3GsAu27
Qk9cMksoIzHaJNLgbAMdf/9LW5lwSHedVrnAQGTPUd3Et1F0IPcjp6F/c5kCMYnzmg4zESA2kd+/
+h/CwLQmaMJvE1IQjKGAyrTyxorArQKVZfUMyknZOVnQO5npeS3qo/JRtEakkTlLg0nnIXfDjg6h
U3J/GMST+Oy7KbTYnVOBoPEjv6DcRzc3n6Zb8qRDRt6crF/23gixRIEVDO6a/22GTEe0BliBblw5
2G+JF7KJ3g+FVbmcHuin03rSjXOQpixvIEWc33MtcEPE7KtVu1T6nFrmAxIqrx8Aq5Ee0kH2DRAr
1pDGADu2znvFMyblKKS2X5+D3GXqceRnrgd35dMHy/jcmIE77AmXqVzyVvoJD+9QkdeuXD/zJe+k
UPUSbQZTEb+qvgXEehbvYy59Jqoq7T03UeQkOFDjRgpG/Y/CJ90bUSDKXfhGr2O/vhriZQNySooz
dLIC9+5yvVUR36UeBczTHr0WiUrAfZCLcJg0J4Jei1EMnJK97yP9hIQ6AHsmIxXZUhAU7HJYrE9m
KDt0OYOU8WFltaL9mMik7MOJeXYgHwoamOUXND8T20TyfaTyqXtDehzH4aQADsewzTpcWez1tDk4
MIzu2IyokdY/fQTHmomL9+41oK74NgBW6Ogz9Qr4LS3nIDSOd7Ms7zbRWwBdzJzIObMHwGW94Sc9
dNhO6BHNw7tpUpkljUZ7Vp7dErHSEGS07ndENGjTVaMdrG0Y1fi5m98lgTS63KN1io+r2rC/YoG0
qAMwyJ1FLr6lPmzrawBLFgFuTueBfJWja3/EhzrHP7/hZ2MLGs9cUN+cnJ4lHQbXIsTUEkHjrpxS
xv5o6fJwboIirsuHT0iQ5oh7gqg1iIvWHCZRLA8lBuJu+/OlKoJDzqAdzSBtQRKo2HsuygdiR3q8
NRs5Yxq0nj31b2Hvh0NkryYgqEhD1YTSZ5RjVvPf5wfKfLfddhtPwymK3DRug3Q9YIUFs1iXXsNh
rybmAOof/v/JZ63yR8QATYir5s3sBqC3JkPujUVroZ4AW4tAyNYoK942yP2NLenA4y8J/99pr387
mdJRNPV2I3Y6oBm+Gb9f0+j2ALT7u9fRujBK6TTO+e3pcJe/GigEtmTSX1JJruazcpZPC46OjaA0
o/UKR3amhIw2nefr2VNNvNptNoGAiK+0vzAS8WTw8JnrlUgpF5dy8GM9eGqSHgTk3uywY3TXiA3v
RrbSk2sxjPLWoyYBDfIcFNnRcK65L8lJ04FVoOmqZzbSWYPh2WagmN2H9Wk234W3YWzXx2FlZYFb
MEJWCam964CvH5CejsFm+2T41WEh/nrawZon4IKF1GEJY+Zffc05zif1Wrv+DvM0CLhhuuXORaVB
9jpk7J32/maQmvecu4KwAy9/E+OFFh9HFRos2bVjML+cqgFMHqew7101vmK6qiGH3ahe3EdC7/fQ
EslWq131wx8Nk1MG8jReEnyMCVxrq9psCJw4jXDTvgfumGYFv/ufDkwRgzHh0SGJk+6X9UM9EfjH
3AIxEXz9HBXylEaosUxX9rCIpB6+u2b7Aub96b3Qaxreza0JebhmNO0pqHECAiPDQXuRcSzeQD8w
RC5n9mrgHDvjwHx6/fZPlKuQ2rLp8JZC2M5vJEB1Gjun0QBJv0jwUjOhQR7/2hY7OYEijGRVVVBH
inaOS5DvxeVqSKeKfzd3dyZX1aiyjlBDyMz0kNMQCyzXAv57tE3AA6qbqQcqt1HlSzLeFTAgu0Oq
se7xT/S9AhEP83DQ8cueKZn4r4xaUQjm/BJd8jDRBG4hD143e8ZEYfIo9xJuV5aRPv0Q7kBV/9cP
W6YRq0ssT7bFen2SHMPmWMbOore7b4+J5u04jBaqBSVX/EGtd26F4ff5jNzBU0z11vV+rKnwma/g
jwR9jThfa2tUHMZQtRF4c2kiDIdcFvYuqstCbL3+b7EIiRzq6FRjPZC7imd6zPLqTnMWMRhgaYUa
YeN7LvUXmFInVgew+QvoBZWsF+tJlsKGHz75EqKKBKibrZIWu6ARd1FmaOYQ5E+tx4m5XP97yLLd
ZwT5OLqCWVzPQZuUt+d/zsjJ1J5oA5IU2O+RraOkiCg/t4n8AymgdimipHuRCRutuEttVK/hLYaZ
8qumQu8Kd5y4rW3Li46jTXg+GEMqYAONpqzpGSMStgorDaCKUu9RiSOP3HkSStJoGYSbThN9jt8k
gRvf7K1f1wh0VA+XLb9SXWz+AnFniy9k98bqkWwyLQQV7TRkisyefWxrPK/u6RpaOtmD5+3v1oFI
t3UwvRkc8WNWHrOjlUuV9hBMxvQnyWk2Ai60KHH3dLA/urrqiKnBb9L3C9D5gWaLg/f98Tbv2eDi
hp4pLNhMzlDBy5SQ8NyrIiSpAm+f8C9WVcC7KM/ZlwvMWOLD7RymPEky2VSJ2bJa/HgfNbcUjXb+
5B8EBq1tMzQ9Gyek40RcivfN8T3bkI4TvheBb8puDDhE3F/+JGwNXcex1IOUofDi3RejviM3zy3z
PmymN0P7+NVRbbkiuxBzV+5xuSf/BOLEPbCxbNUm0XE/slXQSllpfvlvZAkCPG2U37tblkUoKn1J
YRhAEAj6hVWBtNMDcnACFPdNxIuxqy/UbspFQZCDco8pp2xomugARqFrV/pKMBtDMn1iNiP94T7X
TGDIviCf/GGxbyqyS7BrTWoxk5ZEcA3gMgczt5NQm8OUjVhXeL5/2CRRuIbhWStA31BMIYxmX5kZ
zgAcOWjxZiqgmHpjdSBJFan3jL7xcJPmLDKD49SVI3sntPFddbmj9QieGokSPMViHWhzru9DQEAA
xwLakhmw0yFpiVf7nOgHFrUol8w22EGcLUgajz0ExUSlYsFBZE+CG5CXVHKPJphE0jFx04FNv1uh
JnIbpTCQWQ9Bh/lhdn2WtwJZQ3/Awz6y8M7pJRQP+tjtXa2+A/cqCNn1m6/5xvjKLkJZf/5Xm/wV
g+/FUtzijEwnuDru2mkh/evt2sUuwTPgxtMuRJO9tzbM2Rh42U05yoz+/8zrrHnvHIdlmt0jOLms
zmOf0o9+y9ShkS6KoRss8r9IFiEx5zcgedtzaCfguAjqBJ3DJWLYcS+vY4G8oLuAqHMuXP2ol3ao
7S4ah87Oo9GmW7qzttZuy4mJQNTEFw6yaaDduK8Cee8mtewYL42D51KGuVU/LNKXh0lYooo2dW5l
40+Rb0e97416RTqnFRVSH+oYBwoQLu0oaGb+xXMFqR8w3hUguIY8DExvFRCDQ3Q6X93iy7YTdi4c
Os3bmpaY+XE0URJMe6wyn0cOEsn4GrhiHPLiSirL5h8XBhNQYUiU9TrA1Psx95Ga/kAlxUoMhcPF
MHLV37mw9XbqbZBVW0JwDGhE6XCLoAArkl2Pz+GXWAXPXSPspcUqVW5bXPrv3xZGoHvHhXjuY9ui
wKXnK2p1gdZmR1J1ti+rfchGQYOeX8pMkYVGuL3uDpjzxxocHI8NbDIS2DIFKnUOnEL6lTqtWIZJ
662SPShHsRGAGz7sBP/v8nRLIeZ7pmwdRmj8iRjajlKjNoBVRbhA3WO7yVxa+2oPltgAPkR3T8QQ
SYGjD+FGWsjOW8vwpGMKBr3cVOZAmLEOt1fTOL7nWd3lThjvnk1XS7tUREvwvjvoUyszOKxPBIZL
c4s0ioP35u/BUETOxrPdVMOmyZa2BAetLElSZkCF1HV6nnynYSpb4A9cB64l/WL5YoYDil3N/ILc
fc6GjxwH43tDW9neSG2oa0jt/vf8cUtqZMyK5rKTZwLu2XckSMUHgnxXsTtEn5lngTzDPR8koj39
Ikq37GoQp5zmGQIs13VkiLKv+pd+ABpNHj7fQ1pMe7Bdmrqh5a28510+rkHy9YJ0vFX5c3TvxK7h
wT0Kx4Gi3zVYkdHz4gzGoZB+rU92GaAjra9ZBvM21FN8SbrPFhfSm7loRaMMHZfzp5grFy1jnAjP
lSIDYUrAMXfQGY5QkF1Z49hGUh76K7MGdAkUTLhn+qVfZDzT772Idl4yq5BdF5oQfFujFl1g5K7Z
odFb4Agl3oWB2vf5TV0QOUpZ33lNa7KELwQUoUFuYqZirtv2HTR1j5XQxbblnoIyEnIjIeKhY4A7
0ydIt6TIxP8ojWsgtJXjzLi33x/+FdIO85MWgyM6qhJkA7a6uUYgP/Y9ISb5qL79cCNUdrnV8UoR
FbzH4gJtwooTO9HFZCFMEgvRDp+nQk3yNELd4VG/GVvdysIF/9XFcLNnCFvM9sWEG5mMtnHuOFI3
WLjvbyb/qFgR21j/tSMSNgPvoYrd/GISh5sTg4HLxxcRn5utyyiFIa5MxmhDykvqP3IISfTEvnfm
eU8RDVAUbi/fzveBlrGVCTE+hZ7tnGQ9vTavgA4pqWxMI7bNt7cxZqW9duq5mTXXX+LjG5AAEkvi
agWgvslDHCjWT386D3SC4jIO8DWZAHLyLNqNiDVETml5NmxTWOv00A12wD5oVtWnvG2J6A4XWRKF
Nwp3aATgVojB32TfUCFrkON7+QjK9mfLITQqDPaRb6UqO7tGW+v17zp0lxlPteLeQXDouS28eb8j
sh8zmjRpoqHKS+dC/FZXRxlCv35GPcZcSUBrBPl5EDogUOscDLyyKdU6QZlI/w9nwOHFuXdAvalN
bRHXDRyCiuZIOdDCD5a72xZT44poTpPmfCUuRBNRrzV/BrkBxZCgPmFvSXEuZO722l1Dpj/RbRVq
juvvm0TeMo6HHfcVc8E+0kCcFKDwgbkpFXAk6yej9qW0IyzFe4YLFflKcaqoT94/e1Lp8nEBWL9o
HW5loYU9G3C/UnIAHkCMNVYrSO84PKv2IJYoQ2iKgagI+Qt4mQaaEkVd/MVkK42rhpb8y8oUNtD0
YOcErPHctzarJ1Hx3wYCrupliIG0UzlKjzEqEvTd0puA3T4b1Yo5BM7WgfEq6oDGYK9Jz5jXuYLU
onMTTsj39Wzca66lWd30v1++AAAiT7ZfMWHW9leS+ZqWN+hVYdBDijcUSmR8OMELbdjAjpd4dwOj
pyShAlK0YbQXyjxHg15boEaAFMZgZOw9eFExiLe8fs0PgK/zDRh04yHUFm9kyXDDXQB9zhtT9wQT
5b+ywdZFlsFf84qY0TZlTMd/INVgTklQkoTyyQlKDUTe/8bE/EOgjB2p+qVjkg6KJG6w46uxbRD/
2Fk8SxePglVUYWROX+OiEcHQYzlRB498aSjCoBOMXJ4nfm3Vzi4DXZUQk2D1K77TH+WtvX11l6V9
5gBAjsVTHytN+gT6SLBpOdICrQJHz6YiUUk5SWRn30PhG5YnsUoVqCcI/ufqKaRiN6bGSZDfUNpt
UKpAJTo/aZT3LSEsHNlenuobraqS325zVUyZJu/ROJj50iFG4pASG3Q7q6wCFbqueDYjhoCggPxN
5Y2kgvbnxZ/boaajU5p7/tGrCEZUdmcvO4/i0X1X03q+DQE4oWFrAh0/q2E7EkgI3o8l3wUuaQIs
Q/+sKKNRENoPsKPbRsloffVYFBS+Oi0m4e+wl16gYkY4mFPQuMt85Q2m6PNKJPu7ErkeScLjKeqH
PmAQTK4OqOmCkI4qFJ/8BTJi97DpNDT8Vd+9FEEgIhf8T4viJ8b93p0DLfgin5lpHE0bbQVrVIo3
vxEiMcojmcN3V+D2ggv4x3MTQDnVEauxAqmtkAeFsxdEaxiu2WKVNxZy8I7r4iFfta8dKo6Utt6l
fCQVXm0OpUHcRymtZyF41IJB69798+Uqen119maOFF8PQwOysmr9eaSDIQljEa/WvzDSUsXEQ92/
pYAUjyTInAIvVLvgEVtdF9vb1g2LiVO7UPHD/o/uiPRfgO8RewHdICApQryQX6xpRLgOwuHjJ6k2
WiWyNMYcbFK45eQxNfU8Y0iXArpbzgWWhClF1P4RDR/nd41D3gujfqwWRamltWTp3HmGuKlRmBa4
WOJKbm6pZqGtpCVZvD7mCLfFgYa1v9kiQ1FWVi621hYydtIS1Lk7gNKLfel1GYT+v8aU7tssYpq2
hJMSkaDnLYsc+ccIFd2/e9Q5oEzadQ6iWM86E32exzvFmuZJOV7bLODmMfv2PWf50Vbh6ZqRwB36
wCzF9a2sjqJaQfEiCghn9DR5WGbl65MBnCKRuGHySi+jfdyDZiyZ+IDsZXDaa0yV4hPes3kTEkeo
x+RPW7uGU3wclFw6loO5rmerIHZ2xYFvlSMYlwK8MK14KNZqRN5V1GyrW2DiHfMURW9kcu+Flw5M
zNDMNAD4VUrs5K0lyCqbrRq6YOtiHkh3HYw9v6VH3+RfLm2PZsESmsqL9Mq4VzvLKQaUAuXsqSZz
dOSAWtBKtNpiH3ouAa8OWYBqnFDjruio8C7Qwvbu9yKXyrEWRM2E1tJJip4Mh58h48WtrLhTlmjZ
2PdYqhIlHZueM8j0FyZzquL9zAk01O+OXqn0CZ8doFqUq90JYKjQEA9UIGmRauAL+KpOdFVMvaIF
qKOGi/+J4pVZ99fCGKleroCiqqAEwvrZqqdrRIvF3lGRGi1q9JJbIcE09FSJfouOsKdjr50MVGlb
9H0mCN0JtyK1dpdwYTd5mf0oBBN01BGqiuPJ7RvWjIqZDJrXiFlPMC2WF8z0SEKEtl0NzSo73uBg
jiAN1VdSD57QAKxj4TsIyf6lUoxsZ8rCXj2NBiVY65P3q6sPcX4hAWpHULK60jarPfyh1AzCNKQJ
xBPu8fjukYgWm8ARWu0YveP5sfCGwSOGK2hE5DZfQ0LBhROxW9Sj4//G7Dx3vr3XfFjImhOKFZYH
FGy7QFcL539OzsJqoWsudWjzpG4toEYNI6tFjTQYtKfCk0I955jrHHcyGxUCQLJpP9QVrzjF4v/+
nyzd6x37Lb40/3sSfAWJr/vQ1tRVvF0Qe8L0656eb5TrPcJAsJoJeGAXFuPn5RgJOA6mfcYmb9gf
HYvapWKq2oy8pqGgoYXy13F6Q5rzifxR5wYxS4B2g9aO6RUOze2BjKmUo49c3GktmeIkXqz4Co/r
0wMeu2QOCegQKknvmcCGbWTY/K27Vbflo9MbuUwJaC210VxCu3mz/oVS2QfbY1bU7sd3dyc+/ncm
+2HNHmRZDKq9GZjzREFwqWyUi1aLYPbG5fILn+YljLy8J/cnG6Ke/MdVzoC2BX7VgnYv+qE/Ni68
kpuSh+RPgvwswmWqAZvVjCXlNcl3o7V0V5ypngLo0Jji8OWQ9tKmztIRtgBTEnkgDyodt3NttxfY
/Vb31bKi//JfW3b21QLx3KqsrSnEDAAkWkIXTRmfyNUFaEZtKeiez+RLBsJqnQUvHKkytnO/HzvD
yuU+1uDN1Y02oKrkIXz5qk/rYONM/euFAbuWWm8rlSRbJHiU+2oS2TorC+o53Y7Q4DNJeDwn/LTs
wuL3gXcGN41fjrBKUyXmoWQ3+uThVsTOIAORzqfFLqgZlxDcY/Y/ayPgITtQvB5DYxIV7ysOKkb3
4MuiIT0NX4q2HuUa7/pSCET/9aSQirktD6segpqG3uaME7qDBmETffCmuo8Sef+oomFs3yVLuiJm
42PgO8JQxrmFIPuDGfMEs8u30stIbx+SwZdUvSH8mO0wMSchisBVwDW85oQEoTEq6ADC3PFEu2l3
EpqkuxmXmieAx1POkRmiai8hcSUAdcB3EqO+UfTwxn0QayeOixjdFfvo0OiYuqAmuTtZwk24uzh5
LaV1b2Q+VSLvHBsLD0z7UzEwQ8adOJDBolaqe3beUnAU5B5XqCJhDIxw4G4QS8UYE3KsLZV1ny9t
uI8MVWPGHmA2F3UYPtafz3nLfXNfNq/9KvX6FZEJnH8As1OUywg9fituvjCoIhGV+27xjtndYGDp
naq54+qAC4l9CLUuit22Q2lXI6wssI4skmI8AvK1nEeeLkkIsc1klaXkl8rJ+1OWGV3KL8YfWPvb
1lcBkP5ieD3tiewcZdONbnUhMkM9CD7xlNEc15bS+EiV+aGXQH8eA3k3haPTMlmrkPPeM2plRAML
5/2IdbtNkO05zIKC3oxKdF0cOw3A56NoYz0YCjAul84cpPqq87v1rcd13zoUnCpTLqgUEV61ezy6
1hIVNonicTbyMrzx8CtGUdDUvA4XOpKAaMoDkTzQKcWs/rPduso2bwAUqHbKUXGRCHjn7vHA/Rh7
cyO/QLxlOYIPancGeomY8OmL+qZZtmt7RwmkrBFEN5XOExQbVQwpTCKWpq3SJPP7rX5d6/NrruBC
icq3AzoVnoL7Ajb2VS9VBOrSwTInyS3i4JSK+tnz7/LNpnj6IqVIi/KlmyC0kSaUQLJRyH8SLYNZ
Xfiu9Ev83loLCEngrz2rY9no5/GqRuw7OEazxQUX4yr7e9mcE/WPmyCLVQlSOSOQkXtBB1gynvj2
uM5TduXeOSe81wZe2CsAT6lLyhYa9ptwdzhTllR7Id1R/PQuRyj8clJL0Osk+Mtwv4WaRtiisYaH
4RuqgpAJBrSgD0Isb74IdsteRGpXvCmO9/NCufmw1bjSKFJIVsdn4SObXg9BIDV57Qg5Xk+QJ6hj
StB/Dd58R1fY7m9cypD6CKsyqVxxG2hfSmlv2Hjb6a2WRF9bq97dXRmcIGef1A+bdYpkTvrqmJE0
BSM97pyF5wxsuWRCNkc4SCQUoyGoweTBMIP7CjLKE0t8aNtidTN0okCL1deJAjoIJfB7n817YWSX
YncEDUL81YoJOsUPI54q25O9PwT4YvfEG0qh2BIzCB5PkLSfVgZGbuPemy2gx+mtsfpJ1CF9EhEC
Hmgv9jipvlfnJgvvbACe/t3Rpd7r4cmNzGJce60eXMZdfqYg8M2nr1Qzci3nmyjveoqFAoZn8ow1
1qi3n817NizAE3S7Us6klULWNkUB/lnkH3ZPhgfQ/qYId0ayntDVdPhcc5O4g/Jkah81bKM9y9uN
DL7YwDhSI8sBewPpNsFiOWLnDsl3QfstTMsmM7b3CAbbiojRh9lF0pU4T2dH7jO9idvXk8thaOp/
p6K4gpJgd4FiAAlpBrY94xFa4M3GYRgtkp03eaeFQbj/xGXl8a6vUvZmq+1XicryB78PNmNhBQFR
zEFAYaKZ1NIS3I+RfVvaPJgR6K0iAxUfOM/Wy6bZul5rUUtCS1dOCeG/aKSQHZOX1yyWnxRN6g9M
loUK+zvSMqhKz1GxDiztoFvTeLSY7v+wQ7oHzR1b3Yi5aASi/lBFxYs/JtmjKzJ94rmvTcctdaRt
CMZBftul5pEaTTt6MDnZ8pc2LfcYNbAkT1x/aqnaw8/suQt3k+c156zKRj9DSGtDnytZdNG2s/Ef
0JeNSyRlmSLVB9X5a25zkRs574xIKfaobd+0u0QjA9EMhz8ihK6/hJ+np138kfB91LvutfjtyCcs
g/IuG6dmf+EtptBqYFgtT9zfVA0y2/WAAuImmSkvAiXsj8jE7Et17nbvgto3RiH9AQaA4F/39xp/
2ZRqS/sD75p85vnMr9yN1ghPe290NhbYvIKrJ2dlN9FRB1fKwa7hd0KfjoebLkunkyg1Nqx6ppoy
As0MaIOKDryRnVfZnk2nj/pxOGv//UBasfOHqFJO25HBj1vzAO+7s9SSP3h3vJ9nUHq06YBmTqSR
i7wNTCBcX29JoC1rLzGif3EiP/u7t4J1aHNn2ecMhPwLQMzbFVR91/f47TWm2bRZTTYgt/pnyIkT
LTg2m88nA50uAZ/iyIkR7vFmdpO+Y60cqW+uwjaimgC6f++UlcG5wzmsyY3rDw2MARdlobtS2Q/Z
MMA7eyIKCgMn53M3LMtjfb70gDWYWZpWO+XEmm86F+ceA8QSqak4X+p5B4sSylBG/2OTwCfa3j5C
1Vpvt7BVKFELoX9FT7P6+G4Uy8+MY0+diibuGubOjtWBvCaH4rpTe2v1eEsulnH0o+aJ4mfZyR8a
sEsvy44sRYC9XccwAGAlrfazW0Dj9jH8jSorDNVnHHgDqmChETq5HT8BillROqlAcwM1yYYYe5Zh
X9zaoJarZLMQVeNIvqFH9ZX3Px3lGPmoquNl4IHNYaFsuxrNuMgUBZM3kM4/YyBW8k7W/xatKpp5
BeVwETGKbzZsy3qhHh7tT+F9z+M2TVc7R5sq7dekzin5yGNsknwRDQnKh2cAfrQPLMF0Ubal4KW7
reJ7KzSUEi6tadKsayTCS9XNVV+uCbI6TiWYWOQtaEy7bfRNSmxqsv5XqN6WPvTnt6pR/EParidE
UUq5f3C2ipEIlP8qXCEI6FofME2Ed9VXImX/M4+jQH1mzgI1WK1X3vBIz3cDDhzTzwo5fr6DyA5g
rX1NxAImgd0vV3QI1UJzBn2ZEhBGhmLDv4LPh2sLaW+Yej95G2UM3NeA2DpqoFHJObEDH/tABlRg
YUlabN9LGGOFRaHTFBw0+H4Rqf/w/xgiMpJH2DjndW/ZGvzhQv4ylI68pudUTqEPrvDguTYcmMaq
T3qDzRzCA3pZ+pfgSxeXH3lbuOJ9mGQrn+GrXMNHhywFyS9rEZUh/65yYnpeg8/kyGs7cdgPh2ma
kNbEOpXfvkuuWZEbRJwh23fxOOJLVNVAryV0HANIrR4KUDz0xCRbTSIewnP9wQiPaKGMi9CwB+fe
opaj26+e9mFpA9+QDf8Ms0YTDtjDwHkF7XSYethbfaclJEodo/kam0lUrsl2/pW8MD9Bbvogv6Sa
O/KQdLaYcHqtWQq6ePcooEYlShvncDAlwi3MPrfdVthiPk1owcxfUNxFM42ucgOcX9oC2JL6EwcM
OW3glvlOyL+Y+fKQL+uNtknpdCvBKqeW46pQ2aPzNYRZslE8ddBdx40IR4cg56hsiWKksNpVQqCP
fs6KndT7TVgdZ5KTxpJA2p/SXlO8Y9bptO9ccOmwQ844wryLiRP0kC5FwkHuR7cJ/ZAnVU98f+im
LCZwQaqWzthTQkgohITgsb9Xyc6b9xE3qyTEp7/1iB2KfmyPMm6WOqoQ7dkti3OTYuLLuwTp6NhU
zFvP/EcaYIgl6WMyXOd6SPzim6uX9hKuGmyoo86DKYXUjyyn6sllDorvb93MLu0n1WPLzLu0BPIm
TNrIpIVmiAGIPc+24hsKzyhpQ6mmID3vH+JLdMB49ojM0n3a4SXgLkGOPswKLlJiUx+n+xsmWKVn
WnJa3YJsU71pY39FRY2g1SVW172pGdKNw4N5utxRtAF/QmpaS9ld/f3n0T2Mpwa3pTFeAjNnQCE0
CL6KRJ+KIwVwyuXaYtKFiFUuOlNf7hLlSqIYJLs09BfDJJX9fcvlZMNZ7xFBIWNxOJ56ettJMEWA
i2B2eldLRBOu3VU63DYe6m0wzZGn5QyghTUCsEps6tpOTyAs4gn1AfJhBVonuCcGUXD6yQV6xG8u
wxiskvCD/wnEjrriw2JuZRM6PjR85uNOdBk0L3jHM4lD3LrxQeUDKPCH2mpBSYxrIiktXjfIQc0i
uZ9eRLTXIPnwNFUypNnSLcS5cTdNkJVcirbPNwsh8ilzibbD4H0x4w53hM+BDTRK5GGqio4eNiPW
v1/8mOjn41FQIN+4xCwrvV+MhKSl6ySPFSP2+1jttSNdR3RUEr0GwPSa26xjbyQD7NsPYfOMWLVl
UeZYmLtE/Xs9ktq/1SkB/N3joaNGjB/jrbWflPYUdG6Rc67lBMkjpjehW6NqLfox+uMSTn9ZmUOI
VLnWXTK7TKR6nS4KIoO8xeCa/ryvvl7TCFLZs6sfO3Dig7Fre8Yy3SFbj3WYjPcDuqzPHXemCP/Q
IqRCBFXT7xoZFff5kNkuPTtAo9UGIw2T809C+O54vx+jczSjZRIp+5fgKjKUlnSmEiC4UyrfQ0Ep
2ekEb4cyC7Ad1YtjSoN5EBAX75FCCzH6XsXu+/UC39O9VL3NT5MHiAr9+Iwva/m9hlIRxzAGfFPQ
5EiFH19k5nXYHA57rymOEeqJ7bTllfPzo6FuPAYbvv3r6e2MZ8U42mdKzlpRtP5M8J+EZcs2DrRP
7pQXuvgEWZ9E+WBY6a2oDCWxUrz3AEngXfiBd5xu5tQKDlxQNHEOERmZ+JwY4ZE04axuqS+9ZDxO
XYYum4WiIdz35Cw2VbGMiarfBGx0URp4j5+PlFu3CGj+2vkmH7K9VmJ6K3C5dINK4tgPxMcoU5+B
i3S0nYwQmm3+ESVAMNB5kJLzDXWGh0SNl80X5FIy/aT8Dhzmpry0V70mxTBqCKvjmfWchMXzfoQo
ehumoEPR4pcuw5rfsRky54jYHP9LuphvjlgFBb4dq+R7BosigDZ6DVW/yy2oQAnN2tpGSh3aKzmD
ECPlxlqHYK/uSnrXbF2XEW/4QAYLyJkiMho+6+WsChx6zcRFIYpQGjAuOcHntWzftvy6a+rDVDkB
QWYmtl45FngY2va1MIOx5+5rdsfXS7BUdpuzp3u2zqDgF6aYsGNC0voW6Q4n25jFWyNhQsBDWBuY
r1qrdpLzFfZj27+DWwJ8JGJchCJN0V7UOz1C7kFm0TghnROgLoHx4VxfNtalD+PgZr9+88qT01t+
FeACjIjWznhya+Sp8o38H2VMWhWjWEPmuOFlbxoGT/By3aQQHD0ubuOTDL7Z6US0qOD8SN4SFLfF
CNWpClhGS7vm561ZDetWqsh5ZymnIl2yK7Cpc6UAB3HmQ/OWwZimak5iaVtILICaybNPgrF4LQTq
d+mxLLQOjg/7GJL1B4PEIx+VM+EHhKZzE4I3ZXQD2DlK5K/6pvqeRPP6F+gU0Uw0mzytitKtq6Jc
/UNUS09MfWiYH3upAFuZeNPXIE2UZwt+iao1vQiCYF5ltBw+uFfzK9vSgpxlEzashmc9tFem64c3
/A1qkMIPX1umAkUrMZOYytKceWfxjfBAennA7OuFvHF/YeoLCFQRETqy4HA9obVM7GVewqjP3+gp
rq34EbN7TlAENbI0vnf5PgOtNwMiW99tpZ4a4Cx3hyMKlulDYrV7d30R90Iw+7iJsf5aK+EIGcCR
t2NkN893BE7Xhwqmi0YKMRTqEyBx3pi2ay0JFgR/60xvsQkZfq2zZhnn6smDfbfDG5ApwCHgSuXC
ooNIVPG9dUN7wvcsfABw2SIAOE1JqrE0cVXK59ISCMddVvuF3Otdq1cfz5IZ6eUmm77na8rs3B+P
5RFgL0viXU/X9Uk/2CbBOrlWtLlrv8efjkihrdwkgSTuAhUh/IHjRUY51abImqLlJCKyZXuI3bg5
Pgm/MfqN1+0IINwPdLgJvLst9UqJbp7GrvUaxhZAcOEdg+K1LR2im6G288qeKfK84uxHWeMvh48+
CgI2AAA+gC1ud6WRaHhr4u0mXJCJuoSCXrfoO0LWfQkH8322RI6fXeiOTZTVOItJVmRbeh6kJlGB
5sn/rrWb/s8WSPlq+KB4TswdEFRd2WXGyJJhGmjCMgFkPBV57/ZQnCrkMG0R1OBHduX6nZg7F8wy
xf9COqWEvpwLpjBRcPJdl1ZbpZ3+uUGfMgPN/FLdBH1ybg3YNoFuwMIyIEA0Hrjl4u8n1fkjeZNO
hBLYCWhtEA9c6NngIM0+b7YCHEvMOG0FNYk9wtqmEXciWBw+OuDckCCj6CYPv7Ad35IJc7oKu6lf
iXgodTLwLOgTB/bP6zsm1IuplP0ZwyjzHpujaRoqcKm/wTRUMIy16DpLITWXfhYZmJuZ3qx1mA/M
kT/kfQlNnRajbyP8NF1rZf2Zy24A/tjSLeQsMypb+iXKKywxhRNgeUU+pv/QttMLKsRinK+ePGAv
UGhWK0SEFW4BN1SjwPE4WoWqdeSEZMTRl7/Zobd/d/+18sj8GkbQp8Njy8LoVuRc0t1eKXG8c6WR
bAkecN0zqcs7LMCoQ9KoDYlK8OHIV8doLxeY8xTMTcfWcmkZyX9rzCujxoCA8W3eMqYrgo6LkwVn
Llz1tldA/2vXdFc+HQ0AmIMaOtZoZvtPbkRbIHfaPPK8cCKIY+BGZeP9UaWgi1SdRm/Fr1g5AaQy
aYRRQpWoE1yW7CwTlTZTNR4GdX2IfonSjj+GooHO94QUM8ZFk7VVPdoVJN/h9mwwgB9MmDyBhFKd
y83faEpAJlMUEEz68BXyL2NNnmDvO2jc/7Fq6OmQVNJ0x3GA0UzjfLuziKQYM+WVY3B9I6v113Mx
GMfjuU/42/dyXz88dHTeG3m0Bkkj4OC/bHhaHx7AK1948TQAI+iEFu6VOz5tlmZSsJjemI9nwl7w
0y0ROZcfte6CRFIuAOA42wIPLJebx1wxwT3f6W/3Up3LOeNGvE2RAMatXSp2tdVneTglQfRIahVH
XjfX3HbEHucqSUuVw3gw8VwtAQMfjruVKXQrHoA1mHMCsA2Wo4vgdwzhxonCMzJTnzFfqAh1y/ii
RORFkOc2MkniKtoKG4eg9nHzVIhAzqb8BPP3OgYZyeLPjhPBR60nshD9e7bO3LWNBX1IB6WS7sDX
tgpLXz7jQaY7HbnGGYC6azlIuxvj/krc6xQn9Pqn7m33wrB5o7sUqS5X1HDhBYCPW8BGVkodzvJA
zRVtoVCLVVM/ipnKNGtn6BSRJgVM05x6tgg7AaaKtC5JbmGfv7TGfOjRugZryDWIguxhAMCVJxo8
tYRLDZAg5EK8TgrkBVH0J7PaGcgbPKnkjqBIv3SML2JhOjgWUpZ8kiZ8z8Idz5ReqyDVSZ95Kf3k
H2XSpIEGGYVqosPIQvXHzg1EkbBCXHOwnsERw5EeXdxUcrMG3oPDvXm6o1e86/f4LOqNNgV0hnp3
6CzwUeRetwJJw0jKEHRmc9nEOxdYOQDxaRq6o6Mb+6xX1bUGQgymiXtCW3/KzDShNHiUc9qmjN9G
20jgSUiMMstUZLtuxGugv7r32Xa02OR6qdZnDP0EbLNnm9J86kGZEhnMEqvxiixhOZ54UjxJ5ZYa
y1sVieB1uYgr2RdVUPlY251H+NTRiMKwbSL/wGrfxwZbatL5jPUGcMs1tS7TJQJwxwrBuHhcqC0A
F3FuA3kSVknqEp/dIzY8EDMj7TH6JX66J+sTuQBHgD3u4oBSRujrT0Bu8ybpM2uZ4NPv7NB1wkuk
XgbzUHD0N8lL7scum6xMxcXQvzH6rccSbjIy8HINrN7X2YXqjuW0OgbfHZmAib4NezdMR8UMVXHY
MG3lrBlC5SWNk6fpCWTiCakwRUuQiAjcrKtaV8e8aQtODOTL7O4AlCCiSu4QH+GvqkfaGFN84uYc
HudulOpfgJT9O6rPp7TzQcU8HVji890SIvmquCSVihvgSPOjcsAWwVCmxNgSAVoUUxPBp4+QtLKy
tUwqI97Vqlt+I8C8rVh5IZ4aGD1ElIqGkzTHyL2HXj0LwZjkkonEamzHpcSqQRc0mMNiR76QuvHM
VcYR4MJNCeAqgApJJ0OT8ZukJZPCeM9pyG0/WHEpZHICOav1GAxnjyoyGuG2sPbIFzt7WoVgVRfG
yUcGfCmoMSiB7LvFXtDnsiqpvpoGCXB0kVVP5FhaVD43s9ZItiiRzm21gXldP/AQZUwC5hyiQcB9
Q1/KqPJvcajMkxpjh+1/eqMhOHUmD12D6JAUly9JEm5uzYzCZ38W1HliSEoxQAi1llf28660aah0
5xzgghwukpPPOV8nqB1edEbH++6MfRKK2K6AUA6bND34nRTel2jN++N6jspUjieqzqIhHR0DUGi7
/N9isjJag72wWHvBtXKLCl9HNtTfJ2ZHmaojB+DtqwRUcWTc/4+f+HwX/iHoDhAbwSjY2TLjjSob
JhnMb1pywiF9AG4uHK5XMN4AFVqE3YBGvmUCZ8039wdNFh18xDj0mBtDXWz5FPXDcwewlGtIQg7w
3zY91uJ6mJeNtcAxFswqBtNRP1YHswS+JGpIsZHWeXw25nXeqkxMLkIiIhehL4IRvbQ+kYdvJKtm
/YmLzKqJSKfFMHMvWtQFePITEHP5bCCAjqTaJ5ScYBUnxqGRWaU4Nz+VNCKjXqnYVzT3ZIo0N7Wa
hNnqfwhkf/Mergg2iD5Y+TVRbIP6yAgbvuJyrCTtHSdsAcvW+LaOLC3mcc9oRaJJVfKb2aryJcyX
NvKv2byIpGZfEf3GKod58phlHYLbtq+kDF8ATKEcBYxSYsaFHAj7OAHLDik0jGnjS0oDtpOFJ2h1
kIhBDzbJdyMoM37CCXlHywygEybZP6I+kmczMpts9+JS+LdysyXtlcPaG/y8KVsm/b+bJqsUSpRz
R1EDL0/Kfu8vfznroz/qzspc12SNDUsNIojvoG1nEEDf3jFMBp0p0HVN20n7isil0lI+fVAJQ8u5
CHbgRggyJfQK4c4nnsF4Ru6L25Z+0+rR8Hem0w3ta66rKzccDXZ1x4l16gxyxlNffFeZWdIkX/4G
e7Kew1XKeAtHN//XgzMkM/XFU+hMFctXKXD5fAl9MwvHVeK5Ltxd5bK4r4iT0AE+WdSQ736YgNHO
cKK1zVUzepSeXULjp8VxSpWKz4VfoMqwIkyOrP7KUXMa9vyh5pgJQf8EswSb5hod1ZCXUWiicGqa
Ulwfhb4d3bmUMWBvXaNJWtkWnjuUJPQ67XKBfgyD0kSof8gJ4OIXuYTYS51UDuPsKeto/SpF+sLO
NB6zpXQapJiQV0SSfcz2Xvc347PZS2zGmM9lmO7VglVYh4SOcEA3mgndhT3KPMXiY0JoGbIk1PjE
KCyek3IaXgAWaslsPd1mRFIKPYCbajKF/iHz782Nyf3cvPB8db4L5kMxkJvhA7LbfCh9V7X8iMLy
y1mwtErHzzGgfb0NcUqv4qjNu/KsuQtnMbDK6Fis57rQ+HsGEufOFjYwJ3SDBbZERTLWHfAThOa/
dWFtJeB14sRpJOo9gZc4qjXpwjM4w8u+7ToSkw6gQJDEgkt1eUSGHAeuEy5BG7oerXB/UDbQ7Tc7
enrcqy0gJMlezh3MhcpFA/YLaHctHqGG/+SINOnjyTw94GbZIhgGLX3/jBmM114Rza+rWjnFPIt5
FaBhOERyOdzszxqCgcz8dAe8fXaY368P4FOvMYS/KbZwcwd6qb7cOlsmflMbP8RpbYA0VC/TZAhj
KDL90ZU7qA8xe2SnrP4b3qV0IPFvod/0uGQ8dHcb9tp8OytUOZedHqvkFsfjBPu2JcQeAEUEf0P2
x5Hf/Lljw+Wx1SHXf3nc+fDB7Si4YIxasAOJTasCJ5E1SMCBo/9zx0Yndqpap7AAYERWWLR1YssM
IfU7TdwgXOf/UmIHzJfaVVeSBppUlCtti/SQnyeBel7taozTwLTKG14j7kJQ0bEySJAY07ZSvEPb
bmksfLmZXlnVKycj36NteL48HLALp8rFS3jVJtcynrm/JYsZHpB5cl1HDJpPGXUIz9hnPfumcEct
a68o03gPTqn5kCsG75hSQeIureZSSTzujFjLuYqPDpX090f5MZsqjODijA+bwSFTtdJ37Y/jUmy+
B815ajZWUS9xGpt7AomEQakxvx6jiEjWdD/dpo5XmqnxLXRn7N38wCt6rWoj1WxQlWx3aikv0DBN
aWgHy09QHrlUDpbvZ0Kh/OMvS3pd3DCN5PBfjCPWl5z06VZT/dzRhUYYvqsyCzBANgWIXYTmfGXG
cwrSgKAv48PYC3xmxhbU5OQTLL4goTBB6NL/1SLIoDcN9aVIkiVUgNoaX9AtiT7Ll2eGHcVnRTlu
6UOu6SyfQiK9uzkvOCbiYZe1fhyOiupmYq2BuS8PD57nDzoIG+ertbTpmEUc81dhfkjvmmu4/XY7
4EJIDUZSGxKQKlP14jhIHxs1F7wfi3LA5HOhnnII/vdoT0ZMgt5+ZlbAVzYN7wgNDD7TwDT+4cul
fDfmcSffqgMXD1B/bQLbOycEe4jenCOWxYjX8oRt0PsQVr2RhCQ5UcbEpmdbAI/pFOxnf86YjONy
z4X+Yl5kE9YKTggMjPwHwGdOtoNc1KMLQbxTxRnkF1oewyYhCZtt03Gn77c8pFWJHw8iOjHpk1Rd
TaDKyogueydK959X8QBo0OJt5lwOC8ukdNW/347XROZSK7EToebr8WfIvf/ewEyniRk80rERu3zB
gvOi8m3LaJnbYF0512ZNGLxYyunmB3LtdRb7Lq7xUz1ouesDyGT7zr6tHTe2Za7QSiBMBk8Mvlit
X5M30hN0g4SZvZB+yVHEvMXk5goI/+EEwgizzihbAbJIFLMXkuynVi3d/1o7xs6DsG50CFhS4P2A
jHFQjaUlZ450coV5CtE8emA6QzUhE0iaEMt/dlSgx1L06qXr1gJaCtJSsHVFdsV2fy4hk22NmoHr
EGPDdAxs+QUiyBcFascXiZ8jvo+TI6kiR/vhzyE00LWNGXcx8fi+KOs4WHooTMTftuSTBlt+GMvD
rZmmz/e3/qkE/1FL7xPgaNiZue/+xzEMu3M0pRqwMJHTt5rZWNnvwvfcGP6VRhQrhi8Q1gRS/eGv
3CibMbnThcsk+XRGc2vdaJVp66I0z3RandPH/V/OtHyPAOr8cdI/GOqkR3g8B21vd2P8lpt2FZXq
DbMv1D5X442Gnxrq1cpq/kztcLe1EeeyhgHF8fK+lhunTEbfOtbuPREFV6OUT4WBxlghq56XyahS
TuRK+iqpoDqeJt5EuNIaX5Ehy/OZJvUEGr4gJ7KyDJ15JgCpx2F3usB40cPWQT/rIyFjD3w/I5zE
keuyIeCtsybOQLrm/4k+yBD4yPmi3UtcncZKAkvfyPvMVVLIR/OgReW3t8ZkgDWEQqu5NVG0PyjU
svncsEGwOi7g0CoMl7BH4O/uQIWI4oSSpWiEQMLBwd6UFXnztVb+pGodK3Gw8h2JPLXV/8YE7YT2
vrbrftYKjsDc/uaqVJXikSQYys2PQBVgRoUhO8/iwYpZROp3nizvB3PGUFFbobs4W2TnndOcBq7K
pHHbu7usZeBlvmmWBjMyKgseksMzTW0x7oKB7MxpZWV1j4CC8EiQD5jOe54hw4XGv0zr3ibw8bBd
ur6gauO9JAkXru78k7Pk8OVnvv8Kuta7zBEl8t76qlfMRlAS0PzuM/55xCC399T1vR85UySSGTJD
drMAdKrAdKWhEVmLitNEymDKtMZ9+OSKa4pg7+p/5iXjIZWH/Eog3zsmLLO+14REk1xL7X0c1Ji8
cl+IwUGHYGpp8PDNRdfv8BnN3WWGjkHAWTud2jk5S2uUWVlZu9Cn2QU9iNeuZ+yLAuOzQr9eRCRn
fRgdLg8bVtMLjQ3YOSqeE443ScDy+cpUKLGQ+rWP5XsW4wQMq7CoWPoIcXKsxwJJCaB24o1gv7cq
rb0nR3HX+eCj+jZKp138w+TP1aM77HOJuI7qulgsECd8hsDQ+irNGmKKOasR7evDDEoBobubmDis
rv8gJ7Leov23M/XgOyIwEiAbbFvFvLgbHI4tqtSAMgSrULQlZ4BpDXWsbY8uE9LDS3V29E7r5euL
CbYZCGgyoKqunKeTAXg2gwugr4diLchrmbwbNe88opmZ0XQkq1hlt7aTY5J2hM7TGCw7xsiFniRR
FAYj8IOP8GU6ungzIu/wQC/f/0U4TbzQWNLVbxnPyUw16Th+SE4zS/NyLP7y7t3CIla3DP0sdyVv
pHCjOsraXzsWjK27GbXI8v+WBBylAPP6yA4D4cW4Frk/rhOMUtZHP51aWPy884K+7eJ30Z6Xasoz
fSd08s3xLO9MxPuJ2oh5Trj14gKPiqAMYPu7K2PJyELWa2j6CPq/bqcbK29d/xZANbIg+QbH3BvP
pj+nB5dWIm3Q8GKPFcgdIrrPolf2QIzVeCJzK0OmE4gnE/YYFcN1lpVf3I9XwPexEcAWAsqAj1aP
M33rid8raWGwk6aaJdVyifQJXiT7AowWX51f5oJjNlFgeqTkKcMM2dLOFbguKpnU/ExnA3v1WE/5
GDqTR75v/m8ryfYrc7CSKVBfpKAAcg1plEW05sVrGk0S/NX3W7lunAa3OLANDdB3v9US/r6i8Fbw
gdUS9o8nEbXqGIw4FY6WXsq/wzGQ5FoFkIor39kEVwNy9w0fB3RQJ6rj1f9OPEw3s71IipXi8MuH
HRAWOOJ5aZw48Hj0e0gGWHT2XBxwKJYyV1X+KCnkqlYJeSrGbVTtW/N7DBIr2PcOj7jkOde0vrGw
MbZh/Ul0Sf9CeuTLtCFsaKKifXuRb9xCbyX4iFnLZ6DPS2CtFztYUdYcFQ9BmMXNt8eQvBZGDMTa
sUA4vryK6xEl0YTXC4ywyLNbY/vBqG7j/sq/2YgmXhALZxfBJ6xbYGRbyEeb2keuxuDIyg+QJdUq
DPcf93J8IVDOQJozXzxxMSSGZjWKT9ArPkwHWQLF6c+L1T6MsnVHgPfzFmWV9NAg1UlpZZIbVOx8
4nF828NH9JJIW7JnAHtwZ9rzt9Ki1S+E9KdaKMS8bSuklklHKLrBWBPloMT78bgP/W/a8+6VSITx
ZQa2ZoIZnmMjPrEVLNWeR833Pk1rMMcD68wZIF5I+h6JmWv0cQemrWubK39CWDgS55/TE4OsdPPD
psXPWhaaRAAj1VtU6Y2eIGkUXYqxqjLZkuzRcrbw/IQw82PRaPA8NoIEsCO1Y156MD/4GW3vuFBF
MTMOuM4hpUKQLrHHDD+4Q+Sbdkg+B7M2Cy2VA5dSs0+/iBhaupMDFrobC7S/mbpx0dVchZvYMaHM
Sl0OXq3M047lrlABKPEGY80qSxQQmD0+CNQkdL+sbZpQD/AXZxP5nB29oFShkf3DzOT1UMX0mhmc
PFBtXTaqGArM7371NFxsvSmf9gZKlqlHwckCgipS1OKVICXkywLee3SElaxDw/bzypbjvi0WxNSB
EBYj7Y90k8F5+tZy8URcPvG1ptEVXFduO1DDQwn3Nm9r0Etd2PFA1F3seO3VzQ7zRHskCgZE4/Cq
GTBb8S31khMh0vag0A4w8qknDBc6wuam+Z7G9vUTfKjg2itRrwmWew18B7pSch81N2ri+Ef4FMTO
vBGkPiBWvoPRvTdxKkLcb9BnA/5kjyKxDdHr6bLxMXLWyvCfcMgqz5Ga+FTUUcmIzoy62uujklEu
ShMDzEqGWPw2y4Mq+IVwZjdCyhxsQYnduJ96JWEgHtJKs4RCLYXKw0YwQDpViga133RI0zo32pjt
CaGNJAQimu5wN+byJWQUuxVR14NzqK3rDUswOQRqa47pNhITknBKGJ75rD5rOQh7FGeNFi8IWXM1
XbFsN/fV4Hx4wwcytDMZpAJtH3nOJghVuuEPOgPXEpNhh7UGjNTjtTWhQuldAZe9VaLcvFgv4DMl
cYnwyBqQsc0onXqSWp45/WoHIL1Y+5dcFHh/G3GrBTG36JTBwkE2qZ75ka2E7RgIx9urAz5KHw0K
3ruz0fStRk7+H/51wj/b5/WO4IRxoJifNpAqst54rJg0kdNhwl/ZkzrwlSYnYb47m73m4KXQSZRn
C8bpX+S9RG392szYIXsBIwKxZMP/jL2eKZdUXohUxg63WQr5xEdUFtt0EF4r02NY+3uUzn9/K0rx
PbeNxL5Ebqq66Y85ZO0UGuyfN3/sLJeJZm1KDyBnM6hKDGdT75V7UOecbcFqZH86ohVsUExavtuy
GO8OUTxVGMWgQVvqGhmImH2k5uuXXm89vlmNgvK1xJMitEqmWhUyImP4D0jkXRuEZ3lLlafvSmuy
EyiGmJNeZ3E8VscmVnfBygr+gjImJcyiVYY2sZy3y2zdno53fFEuybtAonUpy2enB/QSX6FHwtld
WD5x5TRzADnTGReIyBK6bw6xi+OT02n9rH9PZ8CODi7Qoz/zNcDoX3dxKxS5y4RYY1GTGG2TlYNa
RscEA4HmRWgPNSq9cf5Byfga0gbshBqcVA/W9YbIuEs1wh1ELw8x2xxjl2Umbib8UJ9ckSpLsEbl
AcKpa0AywAmuqNAF54XjnNNfssQSEV5NDnHlUfZJzHfNIrC82r2FIgDOcFjbIZaQEyB9+60N7O6f
aUpmSvx6nZQ26lXeF33D/nH5iq15WfTFUwHY6IYXXHJsnHzixUyFEu3D1sF1NQcQOhYcIJ9vjST+
rQ0zPT64LJxJ0l2Yj5jHbYGmp87GZvyohGCt7+DvKuOGo+pG79uzmJZw6FHRUIb+0qJcfdE1o2Op
qpCOH7PP9OxKCQYJbqmhHlvWLVFmyuoaJ3xQNnErsRjZYWwKDHDRBWsMJ4p0RmP81Izhm//Jd6Y6
1QLO3wqqZKWoBfnKAA04A35jMt2/UasEgkTuWX96R6AE+AX/vc/FwaOKCnjjRfzHif0fd0P6/Ikt
GXEX2pQiLYUlwZSS6YDyfdL6CNCLEMbHbceXdgiZ1iV9APhV0R7mzhOkzAXJUIDUJubtE5yjVWst
m0DNbk3z+K1rwGgFiwrgb3y/BQrCbDX9xWWuXrvm6y+aHu1fo5POU+luoTzweY7F1RXyOGZSrY2q
696x7QQ0SyDRJSURiNL6Wn+ThGghIzFLGYWnV4Z+R7rBo4XIyVTwxHUVHzV7txsrri/ru7uuWDqD
BE7kM0R5C8ZNQQRNrmqWN3QCYNVLp6qJqHmCNnQU6o1XJxTF7EhehqRAiEAzcoxDIwboofny4t+/
hofYe1dYDLUXVksyz9zMUOD9HSHxR9PmKO1079QAhFrnN/CMguPNiIXPwFEQCbucr+q/4dcGwTuN
tSaR9CwyQUHtue2/UtiNFSAFfV1dUHaeMnTMmYl8x4EwBMj5OdH0T3y4Ve24xbmBBhdmBNSV7q58
POsPYIDL2ZS9z420+31Dkl5nhb9oVjAzee7p+eX8PdeE3ItrHBHUOes0sqlIgxaldVZE8FPeWBWJ
DV4evi024xXbQszJDT8sqFW0WY4+ANyHW5gMqpOFGhdPKXp9r8ofSeqsq5CE2DFQbOXb5rX/dNqi
x5F7fNQ49TFEffoNlDWiPmqyUNf+/r1du+GEsLEypCfvmeby2tCiJtUd5WwVmAr3e9JAL+qvLCEB
+m6cyGgFknrWRkrNfbrbE7XMwVFuQDr37DOPZ2ItpX4mcpBkd1izdzhy+B+vNdyjlVzDsmcFH1eF
M8fY8E0+rXIAO/lxSCEcx7y2rmAgKBxVZZWFy1DmOPfpCPTHrbOTvKDyFgpO6Z5/E6O7Q5Nfknvk
27QcwHyL9xsN2b+NkHz3LHHR91d+5bvw2BewVuvmwYL3z0ma3Gbf3yJMrknCTjhyhEp7+L0D/0nz
jvDnO2b/63qFusesahnVpcQVbSCImfGdeKKgXvtrIutF4j0Zek5xlSxqss8mLAZtcQf8/iiHsK5u
gXaBHD4Ftcy6cv/fjn9v9jxorLh/2jxm0Hl4dzaOCdEd1QXrVQ9Q+YmQ8NT50USfdifIPOUct3w+
uPUC6LFzRnvupF0xcxwqlR+RrYzsb3RRDfuRxXoFFTaeQm8svpqqWswRFYfUMj7qifywVpJKaf+4
nFXyHhvKdRYumRWGtjZk/ZPvtQNAeNjsRRH/ymAfXCScHMNZRB+bIl5KGA27gbOA0mHJw3sVJ0xw
CaKVwyAdollwYBLP8QM9yLoy7XJ8twqGg+73ZO+iCnQVyrBZrZsbHLtmkkMaGON2/LbGnpbeyfrP
R3JPWFXvqq8UrhwIt+gSRWBs/yIoIQpBi9EkS5dS1AISeBlrK7ggJ1eEdmjK9eiIxxR1zNlIqBif
E4JbRNARpWRxWRLugALAJJ3/dprw0CevlmdfFRwicPbsmwLOEwNPH3vuIK3VW7s1NEUVItUpkrLW
JmlMf9pT+X3yEsCA6etFwfcUbyDVsnysNn1EaBzN2Lpus0m7gJJ3SSaTG2dlA9IlosgIquxJ7itw
v5Bq5uGxJqxh3n9wYyMnP7VW2ZJlVM5p5iRLFWCxcux/jk0meeJ45oaQRQ2MAulIPIvzdBpV+08I
3BxTeymaKZ8jaobw60/UL3LDJMTODDgj34Nf0+YAJgX+3g511OsE/N51C7jQOO2RysjxCL8Ahe1T
Gt2sxXto0d/vQlMAJR2Fs0qYppTBjEe6ZDDgYFNZ7tqRL4KLs0kGqbDa7LEGYm0MlV4OeQTYSldD
Apop2xOL+347I+A4h6vQo2PG0ZYuRQ93lm2FNY56tBp8QPwAbzlL4LZwr71OOBwIdWF2nat/tF38
febwnu9MLEsgF5U2lDx219xooFdftC4LBsZbj43WhXBaRtQsjWbJM0oNS7i/lbe3onc+qCCrzwOc
iivDwGSjmFBD3M2/LeKVKoJ9jPk59iCadrSHFCh8aVMHYaEqiw96RPLAhHdiwWWjdZru5n+V6iH5
PpV/B6TtT16zv92BXUYGL5XlVZXRv3YivUlt52KIpuTrh4gNngQxxNACotY39v+y6PLpNEGQJ87+
HMbhXqZ13k13D5VN+AugXnBSd8Ku3QqmKVaxMIiMyJemrKv2XwiufSM86FlPGB+mZSU1sQxQIl0L
Y24Row0k4qhNZEoEZVXvT67kDDhBVdHcVwxMQi8in3QmTT2SjZauHYy+c1ErDEGtCv/1CBVluESS
ThxVNl2uRajIJ89FsXWP864YQH9hF6lZd+GCdpQT6aHigKUCPkL+w5AQQegjq/bL8vaWkLQCeV2A
aLCFFTCyccylin8iqY+YrnaJMcotCzAVPVm4XKe6fvQT7zXDcMpnd+XQGrZomMK6x6VpB4ieqVGr
MJ/ePL/AU+CaPJn1aO9I3wQtlD6WqE4SDPWOMs2e2U4ZonKzyu3duX02ocu7t4fe9QKIMGnVV/ko
MTH+PJPqGivSHTpPfQpCvQcFdTpDTA5Svox/Nph+VLnfIcQjotM5/kc7AXo0fY4HIILQ3RqDu4cr
sii4V7a5qt1uDFbvgiOa2JvwMj66w/NJKdYbFVG4Bm5LVapvSvUCxzojze91MPW9KEF39QIPc8iB
abZ68m6OheYaqC7ezEk2DliognAJezJ8Y4BW4IOk29xlO+RVZQJ5mIzed2rUmGJx9Y3iH9MZ26bL
ifeaz+F6NA0+f39vcyxDjL+jnebZehuSLCqk6lajYM11dhvgGMBEMxoDX5fTtw3+pArc7r9h3faR
GLbC2OmuX3AtBcIt4WJ74eCT4mvTRriVab94zQEs/A0eotNzH/8RUKtcJYvtz1gYOdEq4zFiKtJw
wYaPWY+KizdImtYVz24gugQsveCvDde9dNaUVgP3gfHrKvxrdXI+vnR1Rwp39no37QKSRpyEiYHZ
ErF9VR706Ynl2HIYZqfduKM9JrxYgnGCgUvwZ7f8sxA6RTapXUMSFQ9u/5GTFaRpzRkj5/u+DQdv
sx4CioQDe1ecf0WPgXjaTIA9oxdAtgf4o9qhQruSVLXilmwtIFpPr6P9F6kqk85mXEiojEtt5scd
Ikogrtc0/Cmdb6wozH8ERZ+2/GS2TK1ODOZWTr0FQnlz84rZdrLr6JGkanLAAdbCZJL9422xgEoV
BhqFRlzTw0NVAlUkPVlVIZhpBPhTF8stRtKfKbrowXas5SB1JaQJUqTe4OgnwUggqEV2vsZ+6QD4
5/xsL4dBjw0e31YffJKK6knmYtKpCp7BI65zWjVjcztLY/RJO9Z8eKTQFGpoWmgFyDnFlMPq+7Ll
wxu/yO5VuUduzK3d/1bR/3KdCbQEs0OC+NPhPi3NUvTj4+CKPc0Qn17MBLALBTh/E1Pe2Bkj6fiE
wGGUzaMk5OLNezmoc8BCL8tMYXXo1IiQl2tEuNXHTrawWscMgHKvjiqxJnLPUl7oKijiD6Sk5wgo
7Irv7qCzfqHJMjFG+C4ESEMBkYK94IFD06oJwL8DhhceByn6dfKqukmswj0PMFdVO1IzWnOtKCZ8
hVziAfsdqQnkA7QgeMJTKzFUmy7eT5hI1q4eAMjrgRZvOntPei3dfZXftJW59hmpB76yVC3p/okk
frIySMBQKRWoUcR6hupaZ608HIUG9CZbRIEAfNkQWqlfV9pIViFQDPVi0R/G2lyhY0y/gQImO0OH
0J01yvu29ODKjD8ICM8nejtrD2LCsOlagOvCXBptFs8rpU3cCoIxLwDbjS+TN1OuruaMqLvaUTOB
OEKKUooV8gDje+DKLDblYne1mODKhhCHyI1vDus+u7hC8Liz5IXgeklFyMSodiWpA0XF7GXztOos
7fUMq73zRJ1fZHnrJzmfgZm0WAl+4mVLJVA2N1ouF365zDqbXTjSuWPSdv55JWjyZCIJ8mRsoxH5
aZ96KgDNmAqs6QRUIGS87aGoAsdYpqnNRS/PYcduz8liWc5bMMLlMiznJ6UAMMiNM94pbOpZ+d0Z
xXooQDZ2ntDbGcGXuOLRFhmqMPX/E/ejVpMTPaMUm2qgOKXYJf+JrUibI3m3uXpemNatl47a7VwT
4HxzyUjLw91RTPPJPGTVXtJmcw+t5LMVzhF6EjhrHH6XLxm44HYAX/yF/XguQYm8xY8uJQJfxut5
ADCkffyBzOnyYzvok8NREhcAS+AGD1zYF5T/4IM5jbM9Qe0ln/dORdXNiv4xb5roz6C284r2Nd7a
mcyn3dUoTmyketddLoYPKbTeGZuidJSmnJcx6bRyPLCepiRa0COE4q86LxaIgjDDBdg+O5JxDAmT
4uBOL3T4oWTADG+DNwRQTpmvZnk8hZZRyLjwK/F3R3PWGU0H5qHLXE6bXKd/3heOCVVpluCgLQ+1
abquyGi+t3t8Fhfuop97K9LwzsYsv/+Uea1lGeaFVzzX6BQwpHel7a3b6g3lmA9/IKS4W4/d3a6m
A/eOhOohtbuRaDIRUocLufVl1FCfua20+zj56/Agg5AiiGB2PIW4dMo4UUnbrIrCDnGWuEBB2WLz
ceq16JBdtOyZVPfXmkqDIRzUc6XIhGMAEyQFFKiwZQvmqNJ7xQ57M0DRnz/8PLWn3PqMmaZKPCbJ
IC0kNHZxKZ7N7GwroEuRSfyBWVrQKXHqxeEOh+MsN+aHpVxu/E6jRvXSFTch0EhpjaE+/FnTuhVC
+f5JUE/TWVpLJfvuiEtQJNMmfkDzjiV7U7u1XR+PobAwTeT6kSq4e7NErNo/LAIioonR+Gv2UZCP
O7S/6jrvzzhFWvADHmvXcQgD5bwOiRWlgqjCTAN9dBJxYmhg9/5PkNwRaHVMrLNVtwvyu2SZoKSI
7ADvIYSkqI91C9K+v6KXHjMyaQFH06HxCIoah7lrvHXSIu3QOHJ/jNavn0+D1aeNyQFW/kbydJsT
8yC/dIquJX2+LLnffq2AjjZz25DLz1k6oIsnnvTmV+5LaGdOytI2egq8NYft0eGq2YQkpEckpUpM
/tOEqlh0oZKp5b3cNLL/6S5sJ/CieOF6indoDgrQhJRtYSqC+xFRkddB07PrfiEbIrM8i8A9j5PE
sDk6jmCvBtQTn2GhDX4yo/mnIdTGN+PKQHYCwEJc+cJlHsEnG/cf3HtX7f0MTdJ4W9up++K5kX5X
V9m0Z0/PLlPEC56QkPd5ZzCsaocUZSG/0msRc7wIo4RgC87geEw6+oJ1IEJZ7esvjTzsU6sWUN42
zbmvxbeIqlReMXg71zIO5SnTdskZEUmJBi4hZ+Tv7Q2SGuiL0WnhROovZoEJNvLt6S8uxMrd9YeL
521SUKW310cuo3DrmhTi1A5cZanPCSRcT03aS6zdVDvP2lCPokeU/Lhf5WFO2xnFrWOR44myLMEB
yvMMLHiMjBFg4gqLep4usegpK/tO1nea6tKjoxXRhvIwDKtgmbY5ibN1irtsiWt+ogvOXhS6J7Ws
nLOp8oosx32A31CR85Eq/5VMMaErYy16MBzbtNxGO+zwxXBWgDO8jFi1sOuijjxCDlP5pjChkrPS
zB9aLiNHrz8MnEJ8k2cuiL4qbvfUnhm24h0ppNXpkNWGogiDMuuxnVLX7k13rh5NDFCFZcvlnv+t
vN2NSJqPfF0SmkW/pzCpVP8TKAc9zywKKSdqWOMN2WFY5na/gfVP3LmL3gu6H/Jm/GDKEmOe3enM
IJvx7TrQaE2tw1cKO+7owFWsQLqMizX/FxbOGPzdRibX4tnKpUYsSjONGsdfYgob4ob9jBlDSEXC
Go9DikkexmzDZckz6U/CRIEHk1JHycVzxqBBZMZY/14YxUdC4aIbF1lhAP4z3hN3XZgkSSHbU7BI
izM4B33Bv2JOAsYgVqYUz1xtvS9vIqcMv178lCLghUwyHNuRbSrPpTor5hTYa1QGnqHrrMYFUGzM
hbOLXodogtIpf29G64URx6zdxdw5D52Kw6sOC6f6k5EUlvLmZCCH+NKctWly5mqWFZo8+/Swn/M0
iTInrjsWZSRAi5+bMRDMMMERaAi2QkeX4Iof9lPM0DTBDdfmxLMEZEWKCszlttZgfMiybaluowQ8
ALL1IG9FpBdSXzBhKv4PNUifkjn1ts+IRL/qOw1gopHNvTXcr/UFjT2+HMjeCOjAP42Anh+pBBpV
6Dm3jnpNgEWlwEGYGx53UQycd7nE930e5QPZ9LWPs8Qn3ih2Y3nu/l/LMkNpp+BkdJJMv5ZWyIrw
yEqcvWwv+jmwwB8dFxEo6nohCbe0F4jADrV9e9mfSk1shrOWhJb1P6+AVX72splQsBKlMZQRr3E3
2L7sJcWj308YQV67ZlDlEx2uFl4cdYXe3GhCx7mlEG0bHOn6ZckL8u6qfhQK2x7A3rll8mvzZxpp
jGg8/qjMQ3FjdmdR38OsbYWjAWxRtqY7aibv3rdgg6Z5C0MBvbwMw2JZErKtxqkGfd3JX5QFgpB6
Yq0qcBWNqGMsMntwplJyY+lDapwiTzIlv+o6TlYaPl/34v/9VHBHsAVLLdJZMRxTgrK7jslIEFdz
3finJ3Np+7pyMra1BO/afe5774Ka7Fl0kTd+Z0iK+rdUbX3kgoE/SQTmDSH4HMUVzcGr5eLl5CpH
ZiGiMYC/p9MK1stnWU1qeQXHTLqCvtH6Ax9oJLfyBDa6feS2Xz3ZbGhJ6WkKee8kxwxThCMulXvi
mLObHOxAnYy+/2fCDJTGxNK0ty7a2j5QhAcBfdmcR0x9t4Gc5M61x1C2fvNi+ZjD510m9+BoPCGr
T5o1HbKrjIDJ4EuzD0JYbCDUPlMNc8MxSgRtxZC7loucAb2xjsJA1cLpTRJlCEjPW7gijXYa8/Rr
5Zc23JIwDoCz+2Dy51Kt4FzcScOKWcJME83FXInTExfImF0aSwxSzQj1GugDkJDubIWXyvVFsTJu
Sc4yLeOecBi3BHqdzROg2lGXatXC9LhA3OV4OJaP8QDLzc0u1WwdTsxeMJ5Dpd722UUrrtV6VzNA
PIQ3TRqZny4mFodbwtyOahvjTvLnHnL+sMHMlUl8D3xNH0PUeZwCSc5ppUEMvujeeQv7vDN6b9eu
7b5z11F2vDXdn5PwhhYCbABUkNXQzBVo4tvXHVkFUuljswAroGac5oxwOnq32/TiEP10F9Yvwnk9
dthyjsCDmvyIe+w4iZm7l3t7B7T2QsnRlGD+KqPy2ENGA9Yg4GRP4HaijW/P2xfyT1bJg8sgkQs9
HtTkVoGBu0r4c0qjVMMMxLA0hU37HkxupKAucLAduasGjqnPHvbUYzdSKbtYTFwy4OB1oKvJkbFt
kYa2AIMWCt3EcvqbeZexvzgyXX+DQttnN6rmlionTa3pnI0Q4FiOxl/T2rjUz6h/YpKJEDx4ArFh
vAVvp50dikj3N8a7/4MxYqTJUA1CvSAZM8OBNJaJndnzlQsFalqXBEncpL3wXqr8bO10pWIjYigV
1y3C4x4BAUQrfHiahZEQq+aq4hSIqPdZy/28ykWjZIW/4TyxrrmGYToEalCL6H5cPw5lY5SzhRo6
KQzLl6+NQ5d5pwwbhUll16h0ESq9TeDPxdc/R9G0Ix3ijYawfcScne/vNhs8Y1e6hGOq8rAFRBMo
mj92Ho4a+6rZr+u6QS69vx92mEhTwfLIw8IAZHMS2QdLBrYPPvyK7T+bQoXGrZXc+lRzYklbdx3v
IKHNN0SYLySy7WIpDCYJ/NX9F51YbrnTW7xoY5CsHIPROKtAZKpgoJJ6Hnq/ehC7NWv+l77JmwBo
9YjllfLIzktljkajf9dKEgSOi6gnD5uMnmA4GV2YrRv+objHxYpi6y52edBmhP++jJA9AssP2glg
g9b/0ugwDt3MpiAomlRHzBQjqr+SuUVKgMLRCVO384TZdbiV0bpDka28HAbO9jo7ew/EURmaROhQ
Lk+NOdb/WH/KWR6MSTu6F0aZg3eKTRjxyX5un/3SJob84mRKY4vXI9MBXJbWhiNJqoMWd4MznpUP
IrkmKxkqOs/BU6Z1gJsFu46QzKqsgoofqJLjjqWR9ZDin1tTAf9FLsW/6x7IDsJSTJhZCQtYpynB
CrITXO5NyJYkJjjD3sTnatHLenZmwB7WOLURN5VQ4jWdTtElzxtIv9v1Vm2xgl1pXtkyIOxW2ZZb
yMWrKPvTzekS6N/ffkhjA4b8pWfRsh1rjj/woGvYqNDiylvRb0InCs/JQgMgB2q+AbaqvtRC9SVo
4+cGkV06w9mfjglcMuJpYZMpfBYHPcAp1NfhfJkzewp0dVumt0oz+7y5O3cuTGBbXd2nwXFSUwG1
JC+CVvKBaOYx+rvYl3tZ8J0lk4/eD+tTMPe47eGmiBXkoyx1EwIvCS5K91uwpZymE9gfOfOQurK0
zgkFYrTcauJalmtSG8GxcobCSJnFCQU1QgHzU5ODB3I08vzP81Zr2tlrTSi5KaXSE+tBhXp9ITG1
i5hV+qx110IpkY0dbOIO5SCzY3ZwfyhcSPJUCFmC5SjzM4eJ045D/Qywf99xQqYn0hTN2yCX+6Vb
5XLgjNXLYgip8sKMWyhqbqPH9ZHYyaGNdJYxcDHwEOCXH/RvsWE0gP4VZfm9y7b+XFBPO85Wv13b
cGBbWAyBY9OMCNZT2OTw9+cfgT15flJkXb74ukx0DSkeqIV0w9xqwE7b5Xq7UlJKRffbmoTmULaM
q+9F/5PgghRbiq/xTOu8bGO19HNrPPbn794rL5WppeoVbpBHJTCSwgEuRzUQoYaUs/3808mO6UzN
CwQ02/1w7l1nTWcj6yHlr2Z02/o42KtWG2yyDDIRxQocgY8dWOSw/RHtSCeh8N0e1FdwfiMGniun
dirgczRhUCxcXtwQQElwaJYCxAUnKdNDeujgvd9/nGh8R1inIu4UFXGtFOWMB7G1SR6G7wNZjlCU
DTT0RAt8ZnPKHj23m4VsNY7DY8HGw8IwwquP+NNAk2X9/ZzHkksggHEs4aN35BwR5G3mo2Nn98iF
njgAa2e9WGMxlzX7Jyd4wWAPzXRj2ODbTAHG1UU7Nw1kaoxQp7rCac4vSFfBFM3ij0U4llioMkE2
CqvZw62VWwvdr2eVLEBx5cjYO+CI1vXDzXypyQIiF0u7yciqknPrYPBA01EnPIHH74CS6vxD1BPu
D2Rp8csP/WHLsOjHezQin6+NSlHkiHDFvkq0OR3ydeJe+rq/Zs0H6MZOYWkIb9JXtpwbNApqZH9X
6qJ6sMMnblmr6bN61PzJa5tZFA0w6MMiItsWXmjQ5CQE8V8PqKKEhl+JWh//Ovq5FeB+L9z3HmeH
FgNMYoJAimmTFUGhpleUMTYSvBTVH+ToUv0dS9NLK2VpgfASe8RxIC1octVFfTBwW9UyOSez2YGv
Us6f+ULZm2q6c1jUpe0ZjLyHtttC94bqrASj8ckIa+QWjpbS8lwJEo23wnUWoKvAm5M2ZfgQrmig
F5hPzy+s6YwSceqUBu+JneSiAG0MffL0ncbetTICo95y58so+QGtb109V+zYU9rCJ0oHVykxtr89
sj6XdOfZJIhcIWGFazFLBoEm0aHZ3D9w9jHgvMTeLLZVMxiqEP2QMPygizdug9XgQsoc4nFTVMY8
8FvYKkOv1GDumGeoXl4GyeLw1U3PDczZGAWNlPM4o05rGac+9pqjoAOg4/PIqbEHplST1iAn8TxX
IBo89hUqZU1spPAUBaEBNSooN0ZpwO/8BXObeKW4EwUP0mDJctO5dwqLa3/N0HcDjaB0E4yaeof9
UI65CzANGlv6vPuanSe12TrxXIV3mFp3T9B5UabVo58oH1G/SVxsgbtIcgukblkLQr+r6z+PfpDr
xxA7ReaE4A8yBInZ8+R0T3sbx4sDWYSvV+w7EASe39rLphpDUsk6AjgE7nNMPg+EbawqCDJAlgco
QzwxZ7o2JEEB+DKZBbSigfhHgiWJYSuZJG+Wv+R9+bCQhwR1f5DPYr3EObp+X9p3o8cYW4YaZ2y1
iKN1UnKBRxYTPQkP9f6Z+8MdlGZQf7HBTgwwPb7jieoJmFrPxRL40Pw4XcoR5r+mneZMzglwszBk
qB0B243u3SLbLY1HRe4XhpmEqxXsmgG3kQNQiwmCaipSZRvV3LFU44/RTN0n0+EWa+nwq1Gxb66w
nBHwF+qAH/tSHsnuy563EgMo4VPXvDtUI96C+sX7I3lDqpR2uJIKPlX8pjozP3HQZbVg6zLEnMSq
yk+mW9jdF3KAtU6yPLBdYGHp/upTmI0TpEe9c5MIy2qOeyCOT5DUX4qqj3oEPNFMOyRwJPnUZ/Sc
4HwJhFVyXVKRf9t19m0TaXEE8F4IGu+h0GqUlRj2Rmb6rwkaWhe2e2C0/QB9H9w0jywxXXOXd8/M
fkKp+p+3JLX6lEb+iOUK4C40mHXzSDARjVlb1ZICuPIgPPl1IXRhZxiGB+76B8GnbO/M81yjvOyX
Ty7taK3vBUln8QLQwDa+6rshVBgvbiOgxs2AuKyz9mz9mTKSEijBkRsd9kuKULqyYenj6B/YZJCM
G0ol6tVEe+ufgAIU8FLpxmmorKbXgPeySrHIQOo/XFqbuIhGysdkDI3wZRSUd+0vY2Z1RF/Xyur8
djRguMsOUX18/9xJi+YIKwVBoI5ezIkUdljghu4sq/C+Cf8xBD9gprxXGqEgLJ71a0aKDZ1dt2WY
+XG9jDZkWMZCyyFb6yQ0EdbKGuWR9iPqFmnl3rG6DAHfbI21qjN0/7cWY0sUJRbKnXkkJZRRaNaS
u+4odrmho+QIdfCUNj8E6df8u+r2oCYROti+gEeNhroHNP4qIA7OsXdFbff7udSgqlSe7tx9asI2
wfczQkXJu4y0n3sE3ulh/KwmILqwGW3B5+rzpMXYOJAF+ZOngPbo8QiwejLOfUJ1D4O+LYSdD+zJ
ld4lwCFNHOqI8vfHogSW4uGsAPrkv/v/Qb/tOCrAJduNqsOly2mCPf9knfmRniZtH5jrBrRd3jMZ
qChTHbUwumTz22TJQ7QUJb5OwaCRwLhRd2pzQupuMGFKPxMQhuX0sMgcJjICP+kG/y3rT+tiwset
9WQuXNfLnm7bNGXg+CvQLhZgXTbQHJjy9j8oLU+aNX/0exlAk7Qzpy1m7VmwHv+EFuKU6gyUqCQk
nK8y+km05E0UHy9iLOPg9Voh9clmvScLF+ec8bExoK3XLMrXZ20P3Lg+nl8Oqgx6VTKLJIV2s/hs
ezir5mPOJnkWK+AmBZTfRwzeGEJGXBC++/mS7pkCXBvQ3zuWIqYdl2OFjXit+pxK41HLwhnvboID
2xCOj52Tx0vE/1arO5MyD25wO8pwIUyUCboe8yiJGzKwa5Cb4nBBHDqLLLFjShALSFc3DYjwoTcj
bJDRINYQJBnj9zVjCqKM6Pk6iLHcEg1n2QtZts6ozJN88XWrOFSDaXfb6EPdYkq+iNefnEZQ8lTW
S/vahHQ0QCxkKL9QxY4Qk/jpe6Wizm4LWVXYbjCZo+BFJ0LYwd+FtzNF4I1zn30SyfunacCMW6h9
ORAZazbpJrTH8HrvgWo0P+ygd1TFUmUBuJZ+uzLiz4T0rtmL+HJHsuWeee9FvMnfuK/W0VJZHGP7
o2LOamIlu/uI7zjtTwh0XRQldFncxc21+rr3Fkw3JMwpagRrtT+0E/cxc412LR3NxI8djW3M7AAR
OmX7ZAYximxMMrDx1KjWSrvnj5Z5kpa0TAn7D7Q6JiA/dM4SnaRzQUPU2oxGlnq1G2RZLjhnqLeU
wRA6xDTewcTpaRVJNdZZjGxxvw/ogksaffcsigPov0c5BUCyTuxCwwcHE36eF7iIyl7XwvrSmDXN
UwGOnmw8nT/BghF6JZZVvh88ZVDHBDlpArDkMULvCW5pDvCo1XPt6WZlJDcXEWdGzdYwCfm6zoy8
rG2+Aeb/rRcdm9ykI0VIJm6grS+eJB5IbFELFKsrwqnqV9npls4EudPzATLdNUrInVx3LzOsZ+gl
dzN8NT/whkZqFf2d9yL+sYVhNVIqI/05t2Q/+7Fx0BVXodkILbsXKckzQP8bfIEmJS3aMpwtoT32
id8cg6w073Htsy6MR3S+XlVpzxVftQw8KiqkTcpj+9I+oKbMGzA/OywamzhClBvOxvoej7+HenwI
PgH9Or2ymAN/QWUSvHwHzUTk6NiS4TtNjnzA6uvFSpOny6EqBTCR9b/fpHLB1HE5JBg08edId0Bw
kFCZe0duvkv1F2n4VWx/wyPckzP0cWXB4oA2rC+cjj90tjdKTOWClOceY6FI5FZTch3/A617wF9W
+VOonldemhWPUe+iU9+KqQcRUR9SB0pzDeuXVRxVXC3ZqHUgvidq5D/XOn5a7ebZSGfrDfnaNlnC
ELhdijvgN741f9lllOW3ayK9C4oBh1DWcib18U7WXUKFvHeMwexLo4juhH49c9/0gYB4kkq6Om0/
kSVGyo9hBFX0DsIfxlEuq4AHumsf6q8ZwMOT2JyujIj8kZo1w/wiLuOLITnOmNrzloW+DSKh4BeM
wI+gR0rxNp6Ibf/6IU0ZZptAqY00aRDynkMLUim2Z8sKCjLQPvQ3klkePQTK15eJIBy6EPHHBmvY
rapbD+TgYnqQEomuAiACD/se0lEyGrfLYD74fwZjKuhQ1p97LB7l8hj2e88BHc97ZVHUJmsxD9fg
WxjTFDnXxgKGzBBUW6dPkwwZ/H04u68oNncb9Ujw3ysP60ToW5mik4lcolecBekvIlo8iuxp2p3y
j3SrKupT90SOUtCm235mDqc76V/tmQtxuudE4SMxChaKtOCqLXohUePvGqowYjf71O7HGmjU8PtQ
t4WRxCC443LuqbE5aQQ/1FGdk+xwACazWxVqLjVxh2w4RuF2nYVGc0y4oYb+SOJIf6gYzg568KMl
3iDGAREzygHIxoIzWaCOaQjtrti8Qt6+bYgi8Fp34XQzzbjk+CkwRID9Eanf647CFQArjg/rCv+r
dLA1/M/qbySqRwaW5regTIhHqJXh8I9NRNFLQOIzxRUb/Ao2HKz2N3XWJ8eTVbJwc3s7Chc0Ekb2
eJfJK63M20nj1I0hwU/jfFS7OW7aQen2c3+SpOrw5zJklbR+lzUWA9+6X7Y8RCpX81I9RspS5Q3Z
qCgmdAPThnayMGNUSnqjZ6+QLynEihiGsARS3ky8SWyqLyO9FF5Dt0ycv68ZIc03mj+cuTKe3nBN
UxZIpUDZkz0fRozPzKkwVHSYOBehF2StqVDZ9pB9hUCW+37rcddNYZiRLinZd1BnhZrUg5OI/d1j
v5X/Gix2plgNMQca+CvXzpegNZJgSqE0OeQlurs796Pa0s5kPcw7XOsxBFlgLvPYWiditIXWW9QN
+tM9+iwb4BkiY5tQ+HjpPEsNpQxAuLLvV0g0rDTwnMkGNTDuIoXvYE15I7N5ayDK0xPoLYCsJ4a3
rRpvNuXigc/em1C5ektxw2cSKLZpIIh7gIJtPmQUAjN6IkNUEdTq/u4ZLcykaVLF4XmmWz8qRHTU
bYRERxG4UwSWSQJvyB5j/n1SeVtsG7toz6Myne703jHqmpTMMRgirdyBwHjCLT+grGjj3jSwk9fe
ompdyJ8hxmCVaMuRpYLFRNvC5n/E8DE79d3d5CnhPsm1X0JQakzIEtRWE8yjwY6TgfEaaOSZjwFN
nVG8BD415ySaeQmw30E8qzVvqkrcGl7o2xhQP4xHnGAa7OuO+wruIRD6SIvw8W4nQC4NUf62N6cT
9n6Uh46ADeIqiYobO5oFzxpfSj939ZTBQ2Nl3loUOuommNghfLzNLDcDlUJMgrWrVTvsCj6m33rp
L/Vx6E7o1kqHyghWZc5Odyuy2TdgWVITXNqrLZb3fT7ntqOqSmtmm6HRUrfzSxNtTPG9PFakq26u
N2lCksSzqtAtKCSca5n1DyQDIvPasjVd83gsStkODbH5Fk/qhUzWUoiZFkL2wuNnwHUcZ1jU/h/V
1QZee+PASPFmZrXzlxcmzaBvfpj4oBJUedx/IApHygN14PD/cIwkMEbRhvSAUv+8HwN8w5k/LV0r
CX189Un0yNUW/e25ijdGgAUfIl4zyQbUimR8TXnPEGOS3mqmtyjzDIu9ZeCXrnmpFvo6z3pEPdsZ
LZu2Zklw+iQtUW4ttlvOy4TYmdnTRk/7/UBOKuwtK8gV1fwYvG/0RbuuRIdxq24ElcSYszgKX0w7
/hIYZeu9iZAvpNurGPYzgQqMe7wB318OcyvN5xaWPDWRkQ7KxVlfKEzUBzwv6Np4EzDuLhFbqsSp
sreVfVZR9pNO1ysngkqsf61tn/AW9NRbe49ooQKWkaBKALwM5PgDzbUImgR2ntw+drzzdn+BGJHP
VNZMwfwCaXg2cqoa5LeBpQO5ivhjgXQ6R8MfT6mxQw9J8hz7lGdBdluAtiLLesXQ+l5h4akv8Ocd
Qfqkas4klOO6Y7NCuntJV3PHUXzBTiwGYALBwT20E/pklspv1DEqQfTUV+/qmhMaYH5fToorNioB
tLnWgxWxjwhBgSiAh5JAruUZ9My/Pm++Fp72Yl1lVxXTTV92R1YqqV8dbvr8gUqV8ZZLsqliUviz
VvgcRGK37gf6Kd7x7PDSSf7QYcVwbp5nce/efeMzb4LtqcMkxVH270MD8KPpgQxTNgH0v6lF/ckl
tKOWpCe3nVGtbxyGo1GtACS1NcWLBEadoeUmJbY3G11gbkEPLGe+ntQOVpqy4Rk+gfkjdlB50kln
Qhp4esaVdK/7BkZ6UnKP2J9GnZLuALJp4/fG4NINAxOqRTk0AToW4IKEQE7Ra+onhumGT3cg0zaa
b69py+XzUvNpy5NIKqegCL87ZPljXnFf50PlZhmHe053Tm+RvFG4dZmc3COg+B9eUK50qzfTlF41
+Ey5+ItbyL0K0gudQYiT6Qnu70QFIF1z9YF6ok4i7djWlRcgY/+JvRg1uGzPXY2v9worlmanbiPv
kctSfAZkvRGuFb9KeLJeoxKnC4/UPhUnw4Zj6dAVeWWtRoKsQKC7AjxXSRmvnsvF/nSMKhep/Hp8
lElruzOsoS9jRYOjPSVp8sSBEsIfKZ422QRCFMDX4L6hPO2wBjF2WToWUMzASZW1pSh622PEtnth
XyigNMBX0Pq4dNm1iK1wdG5Wa7y614QDvrsAN2VmokCG37k42h9pCr4y1zVubdvJzk9AYAgU/RKb
5H7+58Fa2XaFh+6H26zs+u//6BDIu7ub85Tn2+XHZsQsXnK+fdVtQBN7B0m3hHP5HPwmW29Y2vqo
0QxbDtAa4mmCI0CcWkStXHjR+brJxGVKXLxyOGgRRLFJu/0DygKkV7o7hfxlxL7pzyB/0mfyho3f
UTWKdFhG6Pqna3eZiO5/bPDHrxfJh2Ve9jFTkgNebd/LuwIMZ1gN8q39bwh2ir0pbRWoCaX9fZDX
Yi1TxyC1k7Qfzm9WxU1U4kRwMMR1X4EqPuIrYbxNJY1eZUA7AkHG8t6brQbvnVpa9ntULsIIz/63
Oorjv/PUKchFgVSCNYEpYw8zvvlFqnyMhRjndpLCZUJnFSiwEy2LxB0rXnEWpctv+/CGHnMXvQpL
oWLJYUyYSw2GaMu00EZHKY9NziQuvlO3TjJL4yDagPgLvJ+oKXoGIqIiuF8bSAmNHuc7p0FSqAQr
HGJ5pu5ZX+F8O1C6FySZctR+MXEgjYKanwBMEUEUG7S7riD/xH8X1WzgrQ7zHzAJa08ivJknV8sx
lmU33jQtiNnNNTjqWP47NNPsFQxPG0Wmrt1NVv/mGSQMt1Dzq5jpswWIlr64mubWZcDgyf9nRFd3
mT6UmQr1+n27XhBkqxhMQ169Smm+le9QyGFSXBt9eWXb9+/DywYqnbtiYpYzbKU+69Xb03u0YVq8
1FhqkhB7EbH305N9WCB1KPBHW4gMCks9XS/mydXrCSlonBUyJU/eBC4ddJnt7LMFP4Ir+suI3Ix4
AB7YgUBfBU57QxpDiP3fS2GCCcFPv+QeB9U6pBqkM2xT52BzNFC5Rxc5JXQQqFgcVhepqwph8xdk
UyjLDS/3KZC5YXVz2hHjROcMYO7niwLbhjf2qLE1nQKzB4swvzPQcR1T6yM9FY5gmFWq22QN37yc
8x372r9+F5Tev3X82utV6yTU/jsi+YukZnexlN0CW8Wb9H8xQ8DL8TGnmog39ahrOXQKW3EjYgLr
G2t3q1eWAY4rHKTbDG+hVzlpNyKq8yQveKdGVfQzviLhOdDNCd7s9o/X8UczvlnXRzytLfnSP6My
zH/ahdgkc+Iowjt/DFQxwt5w56sYvm24HiAbgKa3KrzvI+bUuKaae47zim7HTu5KLj4kH8HI214h
yYNPgZH0/fwSolwg1iBhAqkCB3HnJiKO6R+Qjq+hHXbFY/6++YuT5nBFB6z5TPBXttKz4inR2ltP
NFor3PU+6Xn15OMdYTXL3g+1/bjstTfLgdemvkFgxlhpstwPzx72GoDRGTL3xWMyTE0seIBCu1aA
P3UIhtkw3Owjramw+Vq/5SVYSV1Xu2C9kmp3o4uSHXz5MSyiliMrIWX2FS7McoUGmQIB+/kJbFDd
Y7IGnm7uc7NZRjzhqgz5B0HIFcU0m5iexOPuxtBXolk4SeXd+oJ+zLrBewKG9P087BtZs7qmmuzK
VBI2l/NPeX0e4hzkB01xbidYLgtc8XZWl4UmLvDgp74qs6TrFjsnTTD+vaTvC4x++b9fXNLrHWTJ
cB2lqVW6tucYpFNuZlyvyQadoEAubqUS/3WcgqhpbzHvWWLxemyZNMGM7hVTV0FMlz+Jmt+NpW7J
gM0T1QxmUTNIzB84f5nuA6MBdbX3ILHcF+XP1R7wVl02+2ynxGvcHEYRtAken4nQVAwd7VacR4BL
jNSy65uNgAMyRb1UlwI5iilL0QyIYsgfgQ9M3aKx+gWW8/m3IcppYL+0A54ZSE8QukZkfu4Vu5Em
ReVz1RA1WEbOP7PcMgKf5iTU+AwhByyLYAh/iPjDR16NfvK+ioGKpREvb4ahCJopzuFo0T+RZ3Lp
sHoiYBg3bF9SyXKR3qYDY1SH8sh6i8e/IzYmtuNY6nTMdO/gJmKbmh2e7QmYv0XxVNprjNeah+pV
kW7Hf8Ia+tmdXErOBhhL7RRVpuN3Uvw8EoMvw5430Ehxs7T407ce1NMeBisX1I/iw3BehB1z4Xmo
6/g4Jx7gltSNhHpXTn5rz6S0qE1WIePCn4Ev4JNCETAG2HTC55MMH3EuU8j29u9MDufRtXw+SZIn
2ARW4X2xEODnIa0u08pm2DLaxH8agg92tSL0ucb+MBpoKxpEcr2TBsF0BpqzVOBP20tZD3RhKz8B
IffBwWPtCpXDhmVfQs9V5AjRazrg5fQ/YR/K+alN8T25XMiwEiZkc49eZy/kxtEdWNM8eHTzfcPK
czVc9bHOvWNo22Ws8qtw5r4eNciQU08jJLo2xOYVOu+URxteGIi08mXF/DUtzddUKp0XSzyMB2pc
Zq5u2j6dDmHk0iTOt0K6x5W7lIfgKrmWHyp3uBAL/ie2d0AV0Po8nFeEvGGPtWcxtsvw1/TXKqIj
mhmFEYfYmYfgxaTvMHEbcQCCJX7WsmpOpaEq27ZOd79B+8HRBZ3WVsfusM65aYrQDGeWKM6lxzO2
CFXOytcI4391mdSIrYjiwgzMbWvF6FKiYiqrw+Up2G4gmdGhM1TtsgFUnQXlKuosWNSHVSe4GMT1
/wzbRPDgx5/cs0uHjneM7znpj7dZTk5LQp8MsDjRDekDO+v/Jtcs/x9lQUbYF3AIeXj1owuPxEXB
Z+MFERzsjXVgeIV7Kl5LGgifIPLy/rTVPAzjwGYoOy7rEmpy1ZTWQLk6CXsW0zq6ZFyOwYKRBTqj
9bIb/IlaKxndhGkCBqMGoosW/dgI80YZNfmSYVxuTvyqufqOPAF9nPklchcyrD1I93/rilozTMh2
6ECsOmrJkFBruCsyIG3+k0HuPwMwDhB4UoCDxfniL/nTAWEZURcBDj22+77CibSJFcl28ls+jhpi
eE4aCZSAQCd7KKN5GxrIn3zRt3uEPS5HxGFmwFeubzNKzqcuolmhZPz3Em/OYsFRllo0liAX6P5m
wvD51LGeB93K0C318yo4LpnXvCnQgy8attzulsOzTP8A70eQMoy9OVtPcXX4t1roXph25IB8dw8z
zvknoDao62hSbCqlix0/+Yx0wrnct5wsi929SMx18UyGmgg5MY6CE/3CUED3ojZg1OPEFmKkTr/7
wgvDLuhN7WT9uaHpaj7nq/xB4vCWutTPxhPYqJjbkm2be0FIPYpRl+jVUvSnNFTTLI9LNmDs50nV
rLs/n9OFOPstz0c46BgNSmfYcidTj4FxIyBkUpqiajE9KsMUHYh9MfwNx0iuWVgefgd6dTuQjYwp
SuZubc94H8ejI23eg9aDhj0pIFxVpaQlPrKZTV/5Kyv+rtxPMJ00NjywrQEENMIR0xKW8jnFNYgy
AqzduGAziKiKe0NGlSffTcj2b5DFwJBoX7nCO1Cvtffe6e/UI21bVAH4Rw4VwstHgu7U+jesVGsx
TdjVpVK1xyEjHy9T+UaAA7GGcTaF7+8PENocrAlVZnYB0Ed+gkznAk3Fs51npIkkMHkIrOm289U5
PMnfZJTlI0vvCJutQGylHcXjYaem7WtTmfGeqo1k/6s05Ph6zTX7MivTMjNK6vKmJzfpgDdj4D4p
vnobzn5DDvhzG+lSEWVqBiU41qblWYkDOUNLtjphd7K7OfQKj6W06k5omEah5G7ES6r++XDR0At+
rV/wl7TlhkdL2hQDim16YZyfkpr/zORDtJiY81d+szmQ0c8e7srehLE0m2FPVsh6API4atstLgqm
rSf12EEp2QsJ5Uz3KFosaTI3pdmwrOSyC9PhfNiiLvY515QcGNi7DzC03dyl2TfZ/1cwzPnXKbKQ
/kHTvosbS/ksQ0DuMl/wEw/KQrr+BIY989sxRZ3aKBzhhrvxHlVOMPaPRuDHqsjXeewsX8agmf8z
YnyplFnweuQ3l1RKLFBugMkETB3Inb91s4mcYZ1CnlzPaNGpuCFn34ZZHrj/u9Atdlkcnkc5ezqo
KasZ2rm22joDrFvMfm3AwjMaKLDTMkldQF4AznI/6/MkNTVOVuS2MhMJBXwgTl3wnc8ky9QFx4Q0
5/3t/Im6RtdGPS9ane71mAmZBUawpeLxqWBHahIDCFqe0HSBJ2jTGqOdVayfGlb3MJ9GvQgNLsyz
sKJj1dJ6m/+fwu9XAYbE+l9rjBpI0iJcG8754VGfnAYbq3IY6OIvuWJopftBnriQZeRyLxv7fKgn
yBLzeo07e6Q3HLnW3PsnUVbJPRaomUVhsPwLK0QV+DzY4LMzrIaiL6X87+FXcRMA8wgn+E+/USFB
GxIbVqCqiNBoXx1sZBQED/D1Tw0VNctiTfGxc7B6ZFNodmDNFnQIksaXJ/s5rV/vx5QhGdbdypqA
4qjIHfyicRNqyFVhHXMPnfaowYR507kjZxbq3/nM5O/xNLTHIJaR1rsU8zeFNEAfEziwkQ8l7NMx
1Vjv7HGQrZ1echaFjZ4H9uZqqzJ13dy01qE6A+4nqiqyIbTu9+VmQdNLFLNcCk6GmzZYZlkeYsTH
ZGfdufcsCD7NIw322jvX+Y4aFzcWdE9l/diO+e3NbhOL7C5bcRBWNUM51LdxEhD82gg+T7MeDNB7
j9jpo5dIv25eqR1D8zMsf5WCnMA1S9wQwR6/jRkudkRhIA5amP7I4d05W2Yd4v+ZUg/VlHock2D+
3M+4p6lSa7yne6u/ZOinEoiPe3f6SQd5O8ar8kxYLtsKOZrp1+DiiVksxjyUgnJpx9T6RtNhtrCs
Ph+fPLM3gGobIVP35p9zrfv6sg4l06K8PCjyvYTGGX2lSVVLvGZSmGKlTrfbO4TTpfjuf8RJbc/B
lcqR+Lq+lDGdpWUCOkX9aq4Fwipwyf1RA+RqubtkBUsXR3gAyXuq5j1y0YgLDJdH/Bp6nIPz+JVr
Q0yXsHDkiWT2uIfSdIPLWDXGCODXxKPlZdrCQYuxLehYUUACpKCOAj2jTTpCrgHUkICYn1BKooNn
TLuUZJKXr/uzcLOceLEy/gXqr7IBIAXhhTlfGNrXwJ8WsFFsVatA7/A5rWEdF+68bqwQYrpM32lV
1r8yqbxSCv6luM9J4NnqDla34hWHyp/E8RzNB+Z0rduEqEVI/ZxxTsjD/vhEvUdqWpYXTcSDuysb
QH+2vg0RjfEz23km+Y4LO+BaH8v+9899E+qUX7AHQnPjBbNzhLuZgzhjKF3tZz5pIR51uemOIVPg
eo8tUAvLLqyj1ARYdyrsMXNCs+Kd55WwSBFiNJV6WeRn6zCaf74Av4PqdpeEWRz/9VvTpuJJ7PIW
W8lcodDnooP1En50Hn1vzYy9uECSwhJa/pQhqdmHtK1EaxZgFZHqfsmhNHe6w2xlpnKWoHrXydCI
4goCvT+6GmrSqsO7rncFcgLBKUA2gRjRFLMdtCBoTRmToQEOP2s+HKTjKYlzsuGI9KkySfpx3Rc9
pFSxPLOBsduPUxxHBKXY3C++GR2s+IVMklJBnGd3fKLdfWihUU0NH22SiWzDuUiQ0pjgLy4YBzRk
NMTSXlk32iSj7Tobenv0qzj6HLgjRd5MpbcOHpQeg2jE+fN83WRc/CUjk9lj/0vVJlDIN2+uf9F8
rZPwS+TW+VuRBvgxh+5QevTiuAl8dby2iyhm2/QEUrWvbmjwUcVV4XI6uK9D4PmeHLmwVK5jMvos
zdOAk3BIefggO2X3e4bseQ6gJtpbCd5fT7umdpGSg+F8ML7W9PTdHMXCiiE5LsA48VNJ2iSsTn26
QbFiKW4uutg08JmXhuQJZssLYzGKYE/4brtuxhLSztPOTt5E5YaJp5rYz/SRWYwUStL19vUEfUw6
avgvEZsO57x+nvK0iaglZPwyiyxkvjURAzHVNnT8e6AkH1ANeUdGXTaphYb1v6YyhocySUYtrCZs
LbH6x6spRDLzTJZ4qeU2+XIrVxpBVz002Rj62mVq7iFH6nwWDLMMZwkzMzgw2Bri5OYJRvTJpcEW
Q+zV7pX1Q9uiiRJcpRoA5ukMIbYLLGLchuuNzBNX2Dio74bxJC7RW27Y9r2X7F5wSkqhZ0OT2e7K
L7rdrCj+PAK343naK3UJmNq4vmeKTIIst8F/AQjqGIPTyNurBvcUKlTehg+DMOSz6+1uUSC9kmmG
SAkBlFMDoYNiEQUCtoC072vlG2huU/DfCRYuZP4vRWnJBXz5uvZdSlZ+ovBQLszZRaTatJn2DW1t
QRRHUpS/Uo7UkNogfRfzGATI6f0VxIezyU30uSzfh7rlq8jOWQ+6bisbhTWrpusTNmFhEgGGlCps
ddTxwThQ9z8Xa1js+Y6CX0sZTjvvXzsTJ2aYZxXJ8rshB9gXgY5H9RSHu1S7D7MEbA98W9bRU762
AmwJPv5CUMbHYvwWyQvIPjlyo19gFP9n5cVvfGFgJORchiXYtvHSlg5mlysjNLV6UFx8j01fj2YD
DFgLqMjYa6FZb1N93RYZx5W4w2SIqWBXk1Ehz8Tj+hNN2P8Q9szct62gcQ30TJTMjkacKuMmASG6
7kLUqGOl7Utl00Vos3zrGZkd97cIwyagEuoxvoiOYTS/lbyQV4ulhHS14RWk8c+jHW93HXxaz+tI
X3s4m4cE0Mmkj2GVnaw/Y0MZElqTdyBbzTTHbWEZHxHb+LGgkH6C28znl6fvkBGkIMmIGvVxsIXW
2ZkjBdSf4uVa3cCQhuvkLMEWzUYfXtUigLpHV2kzWyWF1NxmA1tsUPiRsrYTCsnH+9IkkavrUPDR
5n++Bb/xp5jYTdOs/hHUpEz+dDulElB/TrvaAq+r8UeNplfNBjaen9sHLtatgRZqsX+hWfp8ardZ
Jwza/q4Ih7AxYNTMoaUz15XhbMXwiyRDAai9rn+0oXDk38oyvTqhNJB0bvEd9L3nyuyRl/KcB3li
J7FtLXLI4FC3IKSETIoYK/eiGsKZ5yGTOsRe8vrzZ6go0FE+6R5kILZnhEsFPudOKdb6UkrBYZXl
CrxCsmDjFeAp3BOiGFJIzJyUOOlngSeKIrZVv/NvPnWB6lGD7ATHiZu9tXU0nBhMXTRcSxGqC+K4
NMT5mbHrVaYzF+wwUopTpD5ze1UZ8s/lUqwfXNuEfZk0KuX5O9/aczmBrkpe5tvd4AFC+8oYkUSZ
d1pBqeMdkkGrDt+Zi0tGZkD33fXn1Gen8Utz89Q93AYlycb/+eFLz00/8Wi9APFCMsIxzp/Su8ff
hVjN2ag5KLYa1FocwjK/EOIv/l+8Rx2VxEjRXZ15PkR4XBtLW1Vu2TDosH9kdT4dBdgLK4gKXbtB
PATysFFHGzKrDK2ZF9HxeblcNhN3DFS5V7fhNhW41DUXUwlmTT/QRhjFVQEQNVT57vMQjWhIJ7ms
Gotot7Do+pET/wxbpnh3hIgPEXguIrJk7Iu6eQfzxtHxJDSK7EXdc/TfcPd4PGZYfZhZl32uIzUe
yusSUwFMxWn/8IiSU9DklJ4RGWreSbePTirstifZSG60RAo0/l4qp+njd5xiji+OMQWqeDuZCL2h
l7MPoOVPhw6DkkgzJJfsRs5Ny7HIQYpfLntOJbt2MJV7tHgFzdM/PgUtzKtI6j6qBjvyxd3VRMdt
o5z+LWtvI5xI99FiukHYtYab0wobHl3xxgJf3itFjMhqfR5xsMgHgz9QWAJMh/wUpka1WddNMLB1
vMJ4GtuvKYiYwegdi5HWX9if2Wwp+NfqqcQylsnxzAgCfd0qsrzduFZzOgZXC/Q2UZQvkgXMd1f0
CmXM4Vc56R9Rm3qdGytWOPaLeNo74xfxQapdG1TOOZH0mGdSollFtWfqrBs1vQShNmMICU57zc5h
gsxDMgSCRtT0M3IiJ+KEncLq+NjBhtybK2LOYQYjejDK0pWpLxhX8Ah54aL/hlnRqfirr/kBqBWO
lzSLdvcJfVAzagr6vih93svnaYzkSPh/C9c/ct56LU+KRndckUMe9ogbkIF9ttq7Ju5Mw1flTneL
u4cHvaLzbB4zZNb/THQKOwce+/5u/OCyE7bEAgRhkZzMdQRx0xOCgmcZ7AwE0ps2/HHx7hFnNbsL
OYEiYJHb78SiPJKAzdZ+A+o9PIbeK3xqlNT4RhJqTZ9umu4q42kmfGwgx+BfWJ5yXGggKf6qGdYt
j7JLSdFv/H72PTGK5h+MW61QrOLYqt6FHUX+/QqdNh9rFnKGWF8nBuTKeiIk3XfOiLciqdJ/34gV
HXCMsv3eFZr3izG6YLuFOLzFZEUm7sI190RpXeMmgmfWr2NQv756xCU6xzMVnlguotnKoWtit6Uz
7XXq9xqELZyf7IztDDJCD9eFPOv3FdlbVJQwG/1lsTt+KkwQCcJPMu5RMySRWoBiKMmeOylVBTiv
Dub9rhC+sVoyHgFPlNQ3NO414Ln0f2Ehzw3SRmuaS3RFfbM/cxq6UHBNdRCBKrTs2JwVV0VGUfo2
2cx5kSC/vRN0erFEg+MLKIIGhbviW7GXelLvZnOVxxoJBtZ5yS4yQeQdoujybSGxA1f4RgX0dcK4
o53oOZaMAaU4qI1VJKGsy97XcLXZjAsOemwpeW0YBPQSqsbXP7A3Q2LQo4ErkxHocK2SsASjSEIm
RhQLc+SeKrTxuuXto2W30zl4ZK6Crhg9RDbKpaVnp9FiQ6B169tl48oiZIknSOXgj0ops6iQUBDr
6RFNXrBoQTufb+8PhkcVh0ipm7Q9URXNjeZZiB0sfTwN4lLyZoGpwDES6LB0NXuHZqb7BHgbhuD+
vHVsxX223G1cQETCtO8FrmNxPaiu4rJId9ACtSK782m9MYxTFC52g8ApZVj7Um8Z+n3TzZKb33lO
5OdyvI7fqYy5wRVP5YeXcVtgQizj/Dc/KrTg9Y2TlgC7rIzzl4Gt89jzH6M+44g+Z5ebSFzy8Zdc
MBJxMoTgDh49wlUusFC9oEErjR/mH7N3gXKvpcCofIJWYocgan+DBPCtE74StuHgwFcbSlKws2J9
LqyePdvEKQ8+vz2Fa7FW8XAB1YQ6iDRTNboMx5oDOjB4ZxuAtcDJWhxL59PYCSioTyzm0lfNaMzl
O3fNZfPkGJS38XGichpwpJ2GvaqEgZA0Bo7kS0yZsK0o48p4wScuV2VgwA2AQpSrfrl8lsrhBbc1
QFilIfBlv7cnNV7Dgjd81K+vfEMaRMNSV8d1qefjuB7kcbu4SoI3zKCvBVKJ5lhp/k3QhAsku/WV
2l2p7wAarSUWFnMlv3Jv1KCj3GxF9mKRJ5cVtACzICtkbQL0zuAfs+pjg4PjN9I8ac5auYYZ9n5U
a0teOk3Jw+pOdPCvHv1saUl26vACSPJoxU5+ka17Q0dtOrQ89XLish+yCzZg6JodIQRmdRVVVNA9
42iZtdJUnX9+nsBb8VVmYkGlRSyVe1PYAkZK+17UEFJnsIWTJAzEMW9Wo1EdD0Vic05GWI0odOI+
CJvVmipmyTbDK77juwLzjhQwjVbcaImFb9941lEPe8BDHBhWC4PP2u7m6Xhn+K3Xf5l8ia6kvs9B
y/n+Xb6hvAQeZvpNX2olvisVjn1PMH2um2V0jdgWz1j/2ZQDtQCJVBu0gt+MhjS84supoBWs59lY
rHYpBtfTEDNqj85T4sUYjbMiicRPhWr2Jo58nDMoc+Fwb5lFlqge17tM2GJ0XF+8yKQ8gYas0b5F
bbuxALVioSw+fKyVyjoZRMI2ncwNkVZnLJdc2ZrWofDKBY62Zs7EMMCIpNyFop1p6gqFUMZAP5G5
TEw6Ra1nF/vZxy4zZuc4Fmmu/z0iKeSkpUSdVWpU/W5UJqIUdtlCtoawGnCDfRngbb93zrtxKq5S
rCLsX2kWOyIpS5S0papDrNpYs9fUcCjt5G6tdQ06HLU/8qb2lEfrfpWO3OplQ1awjwq6GqMtPwmo
FuYhiTTgYfAKLAzXDvlxxsOxGx0br8FeG6B6dhPXif5bvvIWEtaZyYLhHXdRbmo/mcqqgzgD4LHQ
lh88RhxWrvXTU/q/892l7An9l265YBeKSJeHJzZE1sCOgSwdlGNpCYce7JleEwAje7tOjy0AB+X4
jVs4uRktXlpOMlXHxzSRN3WGP1xVGioi06NmfclMfvHxpPDqm2Y8vmw5TmmS2dYXs/0+Vb9hHIo/
tngbxtXXY6oL4Aa6ph+7Om07hSmObYtOE6RucTjU4/Ng6ITdlKm9w5Ss4o39ICH+sBTOnlxwlQcN
5UMql4xHhj5jhIZS1NktNqy2Eii8BmnhMecFBjKeAb8o7ycHiS6zl06MQ3ObRRockY5gVCFl717R
gXiyMOJBkONPtoEy1iCiOJkMsbN4QNzoORIeBIoGmnby8L2sXtEitHBhcw9/Us41iVT1KuYBCUch
HP1ymBcmGksZmr18R4MgW3r7uMRkQ76XQUwbyp2j+qIPW1UJNwLioQUeVdw1K46neQ66xUSsnAYK
LR6wt0yx/gQADzckj9gFSuxk0LGrVw/Mtr1RBTOrJpLyysn0BYpCcIRmxu3kTFodp0cPXm9Fq5Cx
8QIFKXunCOvUDi5a/2dUNAVTAuQKivU6vYr5czoow7XsF6AL+5wQZB33a6317C838dVTGobwp4w4
GaQlkwyL30d+8322tbseflCxqiyxN6KCcNK3aioMy+Mkuld1MJHxWHhJmuIZXUxVGV7iUSfOziiF
ysIVKyPHDQty19JzesksB3WUH/B7YJq1nCTuE3T4bBdipRsC/upenu7pYHd9WTJiTIaI1memquiV
Ssr9Yn26b1f2YES4xhz/8En9tNecaP2VNaXv1JliJuzh3om6VjHou2BwWWEtnobRoR3+yWQ0JPtb
QfbVUtirs6VPTX1EaPEoCl7UjU2oCuo/G6+czBEuwF6leKRtKt3zYw1GyAN7vqqdzwfQOQHWM6OX
PX9ETlW+19EFobuA57HtFarVouI18fN6JONM0sPE2LNm6RPkJZBazb18OgEW75je03djrGVXrIQR
Hy8bfGf4VZ1FTmTqyq7RlykhkGxcJzXy2GNKndRfNNJhe9+2GSkQCYtf7cQA4NdH4aBZjtrCzkK8
u3fWjWxoi4Rhh93pM807a0SOZg+ld2uo9UXMjiZilQ1bN+r0QJjJu61VCzdPfHuRUCffwzoI7iMh
ESb2tX3laVUyZUYhgTlpryXSn4oFpjfEgE5g0a+3nFuHJhncATbqHl6n+XW5zYB2xzp4tekb20Gl
OTngfZPFngSmQwB8tZwEEM9AEYcK548pDklhf+k2SrMsixP6LtKe9YF7dWjQEp50c9ZUblB5wzb7
a5v54s9Yg9fczIHpK67pDDOAC0FpdaLbE/KxiGBdBHDlk3w8IP1trhViyrJhAL4pqF1MTqQmZs5k
CoU1s2G09RjU7XanBGaoyjCuJ054eUC8PnFyj8Mh4hXZxZ1ik4XcoJqn3k5Rq66w2Sh084naFP3o
BCzVq9g7Z6p3WAM+EAqHjdbXw+DjA8TYjKO/0jQLyjeaCWerq98sdzSnlgeaCP97DZFe7KPc5XkI
VxtsETzPNNBnsl/zE56ziNzTy3hWbxWDRhpsnmXikNRqYUDJCxRSFGwDetzGLG0doDufu9TwIFNv
VGbngtNqSCm+fduxERMglghd/e2vZuIWG2t0yR2yRem8Qt5tE/ATIqaLn9ChfsVI3sbC/9eKRe6G
WuJwUQ4BqKJppcVOHFiFSF9Jl50+DPrnAj+ThqMjyUdmqLWL5QrRpGb/mjb8N/uapQ3UYoiFZ2bl
CrTmNYoLxX2DzYy6aibg/UxupyKNSxJHKubaQ4ZxweRT7dpxpjRL755DezWEVGgKhvBfBCOIW4L0
zzHA0ZOOh8dP3k+jUbiNnRWPnjcCaW3UufvqbKvq67URNXOJDX+bGvP8Wp4ZbtWIDRdHto5kIVPS
kr4RYZpwZpD2FQxwcSWIkOsRL5egn8AdQgYt+id1BefK/7B/9+jsgxw6QFaZawheEWnYVQoALTrX
ZB7gtNFyFHFDFdx5SwsAnGTnuo8OiVEG6ldT5H0uhc0VTeluWC1oEmIeWOartrH+dnONi6pa8A8N
AQz1Zgt5wJexCnKALDGKBFh4ybOr1lFPAmsqC4aljxksoKZbCHp0rZ5ZXYgLMQoWaa5urIZC8FRN
d5iJenIuEWd2T/sro80Io1iEGDUWddZz7zBcYHsg3q62SNJwSm2tv4ymCZ8hei1RlB947YrATRaW
YTwbFYxZcOp8R9GsT4zN+sqDn/1umkdj9tq0sVVkZlDe8Qd1HPCe623yav4jpU8ZtejNhqsTJnKK
fq0snBQ9DDewg4b1yaQg0txTGrcszf1hyIZSqI1J7recWPgUQXVSRtyIA560/slMA1pGKvLFeHLt
2e8CJHekK1ZiJjMivt7vFvgw0ZIiUr7uaORJI6lJdUxqelgrVKvmIikZKmwMh0fBa38n+uIYdzff
beQIyr4P+SS/UeYJ/4D7PrBXnwNQVsG7gFMlhYEd6f4R0gxs+0hdm0pjwHg4VEjBmzG59tcwoc/l
O2lAUqOnReHO8XcSicjnmkfBoKQplnCl2rIaAhyUyPbczzrEcpLUK5BiAvQwhH/TbhY1wa3C7sY0
dSTBNuX0vJt+sRoqS4GJK2C4kBH+D9Oc6zmvLVzDsa25ipa3Kx6PzZXSe40ZiG/GoOGFEah4DNKv
Q121JGKHG3u6xHpR2cBlokEYJ2YfIPOgLDF4OuKoybBu/ZfFH58GFhlaaPhlhYi2KNFlJMypOGGm
ceREFuN/T0lfNbwT99B+XisQoxQzh+EpAmduA+WL29au3qbPwpEvkB6t/okkC6sf1Drot+wAW8qW
fy2u7prLQ/kaNXtLhsLGabOc+BCVltGn9BihHQZO4clfb5AcIzpzjNULxgkzxNaVQGX/EG4u0gcO
8ohNW50CAuLgEs9BZR8DA3BltKH/aLSkgafRiABEvd77joeJuxdeWYnlgk+QvXdhmwzYmkqigrBZ
DkSgcj8/QvVKzGs7Bz1uVhH7aVLCQGpPhTwqkqIwfTc3/2/tBwZSmVETx6MSpyogPDlDwcWKp9wS
/ify/Kx+V/CMiPtCyHaqPhHXALdxr9AmZbyyupL3NQfDH8KlGpJTawrjr3K0IA64SHsrBQPKEEXn
Hxb5sg6uhEJVaoVQblKb2T3fs/FeHk61WuHwh04N+ef80eUMkYZsO1ozUfNrJcoHBJ1HZIf6jx61
na4lnlDgNOetuUQAwM/vbsYE5P41JhYXuaYEoUZlmdNwvLWiJdQbIB1denMHo1L2Hv6gt/DOfAsq
j6qt+6qepQAbqsMFsABHAFX3Ckp3wvHHxWgl/vzJEINDpdaMANuDDj4r25xS4Q+UFWfbJTmYIyKI
7JxEbBGMqGL7XSKunJalULugoGApzZHTnYRAR83hR4madqszqHAnA4myYE5qw9IyMbxLgIYl8iSQ
oPQErYGxKYPnKZsgTxqlydliSAJWy39Cc7nx9DqZV6YdY/slgAV1o2umL4xEztQR2L2I+kOjmdlg
0Ep4abfKZTgY2U55+7PbRGQtc17i+Uyk2BrV6tXRr72KsicltplTsgzL9vsyTos787d7jk+BRihV
Jw5C4xc3PngulFPfmGBSjLxmqgoj0tjutz0JJh7rwQ22IMOTrlAdWnYX/UV+xI5eT4j63v0SvfoW
xsnMu+urvu1gpyYvOFAY65dXKTlj+i4UEj7sZRvy1E39Y2ump4Mll3cjnvCcdgJJ9uFOHtMX+AhG
wxp1amfb7ZZ/FS1dlJdI1M3dy9KpSnSSuYrC2OGjxR4K3kaE43+VZE2RtkvN2chs+3gzQKQICcZs
zvWKnsvdvc75iDf7FAFuJJPBFmeasLyVv+vo113kvMco8SXcFw6CfKIPwLQK4+HR25eHLkMZt+qs
+SaNa1CCItP09xTRuzQ95jjLbwllCeveokXI6m152yO9nTWRt9fnp9TYsOTDgTet9odkQp0edyAn
tsjW6bpTE1Q0Mzia0oDOFRXPsTYKxySjz12agjvjt1GTORzmormv2Z7QModmFpVpafyk/dMyTGbP
nTXgDL/XmwE/MBX6TbS7KrIpLGzcDOQbQQmPY6lXIHTXs/alstquNVUrN5Jfm2jGinmSP49Djjmq
+k8OVFEMzVH0H0/T2lcus3A+p0fFJT80Q7rVxcKy9wS0n5pKQhttSGnbH0HL9T/HdDmM7M6NS5JY
Gi4DYbOKg679f5fmA50fdDu5vSP5C9tPS9cJ4IIHn/iITxECg7UMMIHeDbpxCI1ezYSpuQ24Heyp
pRnDd9GreM3pL5prn8ubd6VVbT8OhU6YyR1Fhq0MLr6wkT+1nIL7AaYlAMKzgt8RMDDxOh45kAa0
KR0AiEuK9+4zZsepc+YNlVDSo0OXzkBsaejBNLaumnRDiwGcVFnClKp3+scyUieg64Ezkyhs25D1
KMBUfCVKzQGzZyZvy56ApYK8y+HQq0liJiUHS8SFCteQBSmKfVNzCm1zWB/SJqmzrr6sIGOL5MY5
d0eHaOAJWprilRJRkBSZv0B/foYW3+e9EduEnw+dGdmOC6Fr0ZUyjxzINhW8JmMO0zB1UpG5p4os
feCnRkvRJ7AedJd7K6a8kFVK5xcMB6HVcGH36AgF7ViHvfvjfD4Vfc+tyTwdBzDPqyhZA65PHlUA
eBnqB2YSSfaaZ8Nwy/zgAKyXJzotQzvDjyw/CT119SGlOAn4Z3/kRqfM2KbYjTi5/ixiMxgH8Z/b
H9DjWwB2EabrCWz2UV3FYUbJeRtksKowl5rA31GXk9mksJwxC9d8GIzWIG6MCeRd7vOqZZ3vmksE
EfNPyKsWaYJzeCHa4xFqQ6qnsTsaad/oBdThSmC7V2BnApaW1wlCssgZJq41NGMYEw2boXyoHUjR
FvjFslUE65u25SSSUo4uZ+yo8Cbrswe0/ktqttHWQ9V/EwJ2jEtNE7SPSC0oek5dyXI3Umejy+sJ
lSKHeFtqpKnkAnPMAEdjd2CmbB3YZQl2X5Jza7XvfDDD0ftc/mJun4mzVTlhH8KlKWlT0Oh89joS
HxbLt/zvlZTXQdbPFO4IzqnhVrTwJCNfyEJl35jjbd5RYM7dxoqG0d/YNDtIMlE8M6ah4bluPnAO
IaW9MC0mK4GY0Ukt6iFrYAgY1sWAAggEcXVGi6Y5DWN7yzuxsVAsBhlZOpkyNhb0TcCRBulTNVso
Jtw/7cvQwUL90Aos1Xob2kNJ092Wk4wsWLuQB2MkhPtudjGY1RvZv0JdCPYr9aSxtCQYtCzvt+77
+Qy+tBXWV8r/ncHkcC2z7vRA33dP9rjHwoNwBedwjNg1WrSnl4QJ+DQxOZgmlWKKiXs90Kn5UIuI
1kMrtp4q5nK3MEO9Zk5XVK67PJ3n6jXFrZGWLKSuQn0ZNe2X7KMOur8ZcL4TDumFV7Y81G7qpqbb
Gx4sbOrIf0flJ9bdIJKzQnEpbzhuJZeNNT5J6j9rW6ryfPoCYmD7egFJ0IJkAjQtgECeBpfmHiEx
2UHfo8dzf38dao5mlBIPynM1A4vN4MNErTx0g1gBKReoSreFoU0EUEUUmUQywnsUzlDbc5S/M2bo
ZWzHfKCmbOJ8xaVN+/gCTY7d5kmzreO9rm6MP9ALZoD3cxLpvm+SUhQJ25NtBfHc8ZGkpDexMW9y
ccBzetGW/5HEQMRgCHtsD/TLgNXa5uQSQ6ALPt7xVtcD5/aoVwIKMU/oiV2KSiTiDMo7cNZohzOA
VRebxoDgwR33C+FGXFgG9zujLGD7/1zoveuioiIc9UtMDAxeL7S5PTp9gN1Ht41fUi+Jqt+V+QJ3
ZJnXS/J51wYl/yVZlnAA8lVAT47QiwgEJOAhS/qdKQpNUPjdgE3+U+XGn35k8xUVzltsWhnLJS5+
jmmoFKDv8PlWR/xrQR0rlXR0Wwe0LAfywo47g3oXngSXf/5vkE2GrUDtFuFFGy404o/NfvkTquSE
GzbJY1ecpl+a4YxLcPxd+mQmWy+Tq+drusb8y95oy3wcHtpXHEj/cXfjH9fL7jEgIoHPGVFsgihz
LsiaMHSdM5d7IF0VhM4qDotmRyt3DipXOByTlrWUn1NilDtSoOK0W3niAvIC1bvUCDkxNU5OaWl1
Ki1B3rZaNDTGJorWUxCFXUOe+CQ/e0zTALc8SAput+s6N1jKKoDE0FKO67amNhmwiblZ8xs7HSmK
JkOL3GysY8nDcEXcrdConie5yULd+GaJUkeYH1VmkS7J7lFktd1buUNOpkXfNMsPJWG1ToBydMHj
7I/XWhOud9j6UKHvZWumOgG4IVSSuvLk+NDqT6XWLYB29nION7thC86Ms3gcMLOORa01Ol52jjHN
01TFyxgLZGI/9o4CoG6AFTjAkYNWQw+DpojelPrYxrNy9OfYWDEWxOSLISCoof3ifacN8qW6gQz/
Ej0zbTfVf4RSj+vxGERKIPDrU7Hc0PeutSMbjnl5zz34/91CZPC9munYOw5/WbPJbrrbL1iXmKE5
CuPyOAZjT6sKM2l3u2IEik4uM4VquYs6A8qja1BNWOICEWM9Kh+AKmKej8LUiJake9TgQbpyfbtn
I4VxO8tEelZI89Gz9ibGrIfZKiWZOmWLnJBdQT4Giw6HM76KOzVO5ibrMCM3L65iU6m/xc7AsYWO
3vjHLhP6pWIn/iIl62u/4MBqweniub5aNpG498Zi1Nw4q26WNj3kLrmo1agoL1iojZWfv+pb91ui
dqFpN2+sJqEgcKytRi1mJuYax+9SpXxP2gy524Sv8bl4KG3sLOOqBYh5gxZE7PF74hK1Fl2SChze
IB8dhOqfWZFljopgUxRIu6+NTXVtwWJR2JR6spFflaBGR5jbeLaUv835XRWZ5Ca9/CQrsM64+xjG
GWr122UM57uNMCplvgqHwwazeu3E9hnL3gjruPhzZ5Oy+ubNV2mgfpAYj3gYMkIaRgq0K4xmklVt
18XiT+MK2mQkHBLIxkoRFV6E1ZHafHalsnx/wAbI438il+gWLnmMtpZ5Brbv0DTgWECE8bLQZTUZ
XmwPPaw3ug7DZNqZopRZlp+zVggaNxM7mS/FUJGMYaT9OqxzM6rdMCAp+zHWNXhZNuOUNZkBYdTz
CkV1VvcR8o9MgSaE2vMiRF9ydp95PbBsDvR5wu8GkT+t6AE59JZb1W737ENIbT6G1zXjQ5s1xlXk
fAX9gtKvylX0JHq18O+ECTMM7xN42mbI9TyumU7rl6x6+n87TqRu57F47IPAV4Tfc7dicllLNfT3
MwQe78xKElH7POkTnVOjXUD+zf9yLKmFpHsC5wo93iGpKH/iSF5jwu5NFs+PNgwDK4FqTMtdRaKn
8tGY2dGbWjHb+DTNGvo7pCUjll/LQ8RYbGb+WLiZSXRpx7z6+5yZ7v5lkZhusYbIljVFpszKETD4
rlikyqQ8ClaBUp1L6cBihtIxC+7qB0J2jqWHNue2ZKvD345o8bpVhRiC2aNCQyRp/aJtrgJI9J3I
le4cYQ4SSdT6OJaRcjlgC4Y2cg1fjy3d5MY6VqLUpQ8VtrnfRLqOqnddQD+FsFBDppMUH/4cDeoO
S+8wKZhg6mOHFREC9PutjzNJMrCowAlFA379pPNCr7IV/wTeK9fxt9MLWLZat9bWbxvg2rRxjnQq
QdI7crHFufiLfN7sTZo4oWOOXJo30VtpdbEhJtjfq20oO2GRuvhz/jvwATfEEVCtb4mvWHd1Ed9N
CnXT5VPTRsXXQQhStm0UG+W0fLwh9rlyCrQDKsG/DOCOKzNsfyYeTUC2GeYMwceA16hrtWR4pqaG
f8gedKrKkyE7DS9u7xlXcHxgyo1kaicRtkA+xuGolpDvuK4D+QC06BvFwTp3UVx9jHPlupS3CU3R
utRwVcn8LhWmGrVIMKqQ0qXdh5hQbDOqrl4DqjL4tz2h1YhcnusImOsBJAju5zhgzyMsL5xPbUhk
fJlp7TilP5PGgdfQilEM1EOoUP+8pItIbuvbH4JjPfMfPyoc//JHwUnHjAX2RPJua09YgcRE8Yfa
jMWM5qhvzcg/hebg/L6tg6I2C9hnp5tR4iReCd0+JfJTkKFhfro+EreuEAUgNEXANp1WHAto+lN8
B1p31fX/k0JeNTqLshxAeQLA+5iOmBcNT2m/jRjNaH+erTTsE9J3uhrmX1a6ckp0VEhhnU/1cZ6b
tnGheCnSi26XOkIyCtqnG9mQkPKG7JhM5tM1+QTmQAA1YUrVQ3l4n0h/nGkouhFuW1RRg+g17vC2
Ts4AzFosC0fKStzBeSdtP8eI1XMNqR3y/TZ+ego/G5Ao//cMRdi4fotQ3ikaGDAeTYiKeKDXbiT0
3RLu2UnYuy26RlGlNLoM0lJgtZw2z10JZE8mA0f7zfc/sevzCetEC8cqxx+F3IFZY6j/cAzWI4CP
bOJy+FYlvNMwg06VqoZibDKe69NKz4ZBV3MLqpYZEcyjx+RNfVxqAD1yQjoA5DDEStRNEPvnFC78
b6eGsnhXL69Zrv0X+J2tGcGDvpWYU1EbOJkPUT0RjLIniCzEz+TtQP7ftdWVROlo0YZqViv8XuTD
RtthkbjobN7+neSbkMFk3KdmoEJc93tXZmIeWkhqtypU26uGdfjIr/uD8It6SKMKe1UDc+GYHO5j
4NP6Rj3TSmLB573z1tk9dESFX8braZHAFaXqCJKwlTgrDusqEICKAImfKWLsC3su5w76s8orksz0
MNp0Rl4Rz3+aL+F0s6LLxmdSLgEWka5HNDB27YqLFXKnTYCsdmKSzI2spWmXhsLSYDkeUHMgC+bW
CyDzMYJM6/mL3snun7FL17HQ/B3mA7WnYGx4jJHm9zpil21dovsg4tA/vC9xdtxs2RV7EixCL4Aj
NxZoh7bmIUcdTb2mF9R0CqN8YmI+smWrnKcch24EEMm25UHyGLRdHw63wcluDUBZtVZLheJQzis0
ofo44p/GwT+OpZLKeXrniC+6oWauhX+CZ5wSZuntxSZT0oBDaOly/4MLh35pf+xJ1ApPQP5U5auT
OWj82y+39YPcDZ3ait/jCPP/R70FAOcjUiCAHK3JgZnLqu0VRSET3RbgBLbnc7wiM7pnPrJkBjPH
NWCKOX1TpA4FU+hawZ0DvQTJHdE/QQUwnGXJI0B5i/qY3vsAtWoaxb0Z+DcjuSgejZvAmNn+tVw6
XE5mG8ifx1z0V4G0554CCzxXnDOuGhSb+sm6ImZCCMXpq2n4mhSnVUPIBRtsVMpjHV6gyF2l54dj
xhb5RaQkYHJdvPlyPp6UP6pcnSraQbXW7w/NpyoQheji1D9gJ6wvLAfUoqcbLxp73nRNFw4GkhU5
yQjRCK+HV1TRZ2mj0ZST7oCtEvAn8GSqYWtjTRIjZOrwgnyFQXGiXs6gtf1iO4jy5Q6Vh2xdeflb
4RO6E0Q/9PQVFjC00zEjg2MLIBlpekxasJIB9/v+YbA8rW1DXhhHlhIHNysr2pcscdM5eOtj8n3V
dEkqdVj4lW4tlxLP9M47zPUWFg2w+AERNHcLu0oMXlqA0o9XVOK9EmnEtrC5PZCvOdgRVle0Lrr4
M0A4sO+3k0zPBYmaM78P66057mM2N0NwVSC6uuTsI5uymAZW0Pmz7CtCQJMHNhflR/FL6UUMoLRN
U3g4CZjpnxITI5llR6XjiAfjsQVJTIxyeTGaijgSql7jS8HLHBuLE/iJM09IWjVMkqf3UOuHNmHF
x1zohk6PCDiOaUEVWmJJANgLImGK3t5GeB5aO+pAEDgHtFYWnavp7Ss6AK6dRvBDxcipb8O6wd9Y
8SlGBu949FEqCeQDkhrV0x+lxC15Mr3PJERiEEPdXf0W7LdXY4a5mTdrCnwXxKYBq2xiexCXomiY
hTa7neslBeNXvxVqLfiTOFKbGxCm91EfSe2L6e5c6/5XX8Kg5MfdNQX7py4fPeiizp7kWvLkzE74
NeaqDWuHEFOr7zh6G8zOhSeounZKGktOe9ZX+6GPzF553pGQ1gCoQpk303kaFVm7DBwZ1J3//qL5
6lf5xzM4jG6dWeIo9rmwu6E/xq42Z+s9Azq8zjehuLWetZETHIhCbcrpl0Vx8kl+JAHw1PD1kafI
6ZrTiBWR5wH6L3CiM38iiG/EsEvID3GBDuhsAbRv5Z0MDH8T5OodZHUwL2FdxG1yxHhGOTXesDOn
mcisdIrxDIIoK1KsxXYiaPF+c9SaVprK6td2ei5M74GlbqHo+btUSnjGsW/MW2q7wDLG1GOl4X/f
4kow/rlo696weUcjirmA0jZPTnZza/fVuWKvhntM+lzyVc03EYEgtHHCPtvRIag6AIk4c4fZwH6c
SPrP23bimOugjZ7G14sEc4OHdq7FFFGeBE8WkrDLi5BqVvA2UAYw/UylFUdGRXJIxR+XGr6wa97j
cvZ2LSsYgIP81i5Bb2CP6pzBo9WGUW84g/BEA3/5rbtX/x2b3He9882kJ8IUgYGXolGqaK0sodFW
hxooTtM5Z8PNLzDFTcxAhAAoJtXuPoJypIwWAcGZd3pQMpBmcPFxYdfIHsNPiRxCe1SA4deX2sQL
pFcfwD7AMola9gwPFtt/vPzT/rc76MIgxjQzF+uyjqCz5gc7iGDU4UqxYaMb6zcixAr/e6LJHqJ8
8rospTZzrsMaLO/ofo65v6/tbtIaPOpLGr/0SiVz0sYlNtNBgN/0e62x9gO4buju+ZZdibJMGonJ
PoKerBZoxfIujkEjvk4M0Nf9F5Mp3QsWxJclFJA3uwxMG95GST49mUULNaKTDYxsUV6AG8druYHY
CJcHBRqFXIUyEL480zTwdqWf8xlh0pmWCymKI1mrN9ufOqdoM0ZMFOKQmOrBjtDRaERRRhoVf6Ci
AjDtg5bmbHJ64opoiebHbym7VFOE6wQthuI69rBwjCTVS+WkULvK01YISeNiwRxtpDmZ8psPq0u5
CIbpx87v37hT1JZMLtGoQ3XeEFzY9th5Bbbj9oVT2PBHRQ9WYlqhi/vu2j236bhJHmh2/KjKbzCs
aOtdFDnSykdbqX2TIiAViwgJoqaYSdEe+zBDbQ3EapfM0mqIXizsWJs0VmIcGoZZMx+gByIi5U3N
Ji1mRyTD4Mmi6QlzSEcJ8eYTzMT71wb48H4OuzaxCZk3zY82jGQSBAWmHI+vxWQRQ+vLLNk18kLG
nBNBMW1O4N1AyrIIMsuZtBYtOe959ZwVJYXm5URYSxZwRpL0WG89ZnV5LKxXkV+PSDXkBRFdizXY
ncaqAoBeAF/zwfsIdymy9RjYUhm/QYbwbjvl7APCbukO3MP4ASlCVm9hmNvIpJC+6DJ1V7X4p45t
pyRd0BLP8sp2/TDTa3VSR0/uAA7EBALV0k7DH5cBYcBEMTGe00eojSwSrbs5cA+4N+vRgqpaVrqg
Y8jxf869hHtUnqOVx8podPAziRV9GQDE37sHvr1Uu4HzWshNVF5Nbigs45NeA86gr0qcpkLm8h+R
JmdTmHmlF57yriwBQgT/TmkdF5tozFLi3PT3aTgtihIZj8XvqiN92GsNEIm8heqAEcqkYgZ67xC8
CtjxMNAAlPFeOYgWUyeGSmxPrYJhKKd+4KBecv70As2oP9bxCw6pWLkjHrhIZQzjJ0Vca2+MhAKl
BxPT/Xt2EXcR0AMVLYnxxDhWFQBsQg3RanzNzMqVs44DMZK8WQQy6awmtqk/1xwmxy2BGU3HTBBi
LeU7HDwxGJna0EqyFGHIU9xDy75OYLJRe4m91YXKxF66olP4KO8oWTGtoUXtqgPCDPXS+mTXhUih
qVXOWHMB8r3HmjXIbDirF4k1jF7MzWnFKYeMMqolcrlhEFrYAPwG0RuFsdIz+dELJpM0Isj2Vn23
tN5LS6WpbDjKruNmpmvdzGWUrLJnPfxrxqOxXeWharcKG6OzfPlynu/2+k1x/6bQuDxD+c8yUoRn
Wip+j4ADieInLawYI4rXhHgtsvK/xpUaliUJrJhVwUvJf6Gw9dRFLCf1Us/VApwZbRSrsV4Dct/C
JE8+RaLER2EkPeAw6uy1ZaDAemOiWArSzO/x+x8859mfbV6uNGuCkQ5jHM8ty+7wBGVEZCSaq4/9
D6uSrtdGCi31dko12JdQIM5qGNS7NKAe5DGZnUC+GM61gD7/aoW9GziTK4haYN21Knjt1ZXljEyM
aoisZF0Z2BKZuhGeMWM2XiDam4H3bjQZlqEu21cjxCt0gsfSQ1ROqD5z/J9gnXImZUPjsNhVWzvP
Rv1pqVAGBLEq2z5GmNpgwLqQm5WtVZbRdstddwYebO6ipU4W8o8SMf8gYw1JQZERHlNRjSjIUrx+
bcQQ5pSxuTdefsR8S6rrrxRhk2+sHedsOw3Cw82vEFKhBARLDA/UFR2YH+aYKy3XwcZUfyflg51k
1kTCv7ncI5A4/qBOFbiLMJHLUEEWG10/CPXImJ12bR3VLRpdKXDd8AOxLVZFT15/LLA8Hj4I+Ugm
SRl9rREM7LkcwNcWfHBd/I5Lw/t2PW/TNkZ5+UW75f9F/XyFrqE8CB72MHEbHPVLp90Hz+ss2yu+
ALfbi140Sb4VTj2yOmLC/8hvmwWm3hJVkI78bpvuk4Vf+GCZ9r391jK2njowD8HLnsmhmhlahwjF
IGmTwrH68zjMYHp3sGX6UsKvjzs81uKG2fJQwxWQpfn2xq/JL5fqjJYvSX6rVa9MWUKvpXVlQjh1
E3iq8OKoTBHtnCff1LGFV1zAyz+/0eZDF32nDYv78VbcHIqxNA0zfo9gnUEeSPLb5kEXRKRZLF9r
unaragJUUKSZoPlUPYgb0QhwA0pJw63fatW5lUB2bMICwqYa/x/mLsyiWCj0CP+VVMMZp1xFp9oY
V51YV4QxG83mULkiLhHhty8Yg7/6GgDqmCfIlEsREA9IDa2UPvOdOY7cxpFwtOClCbnDs1Y/7YhX
1XxeIyBrGhu2M+qL3ejulKoQ7ALj4h834WpDKIri9IHIG5zbuXRNjXEWwxMntodKb74dFw6vD39I
v07T/YbIq1WLyQbA+HnlvX6GoXCIQPG7gBOYKDzOireODx/i7PmKW3kHBb57dGd5Cgxkxt0yqhDy
+1uuOjxaJmnFP+1DW5ckBCT706NK2FQ3lrauHi184pcuJ/SiFv4zu/XAzVMove2Q0ZJpschwcL8S
VyY67aZfXoViJz71JYnPXAOByZD3JEX+qASvUwHR8lTJUStxVVAxr6i73SQpU8CQV0httn6u/6XK
xjdOQTinJeAHR62PGXfMQoOM1iPLuh+W9W9sfWCMKeWQD9G3viH4TRynfrFM6gqmieW2N4PmyRea
lMMi9U1XFclMpUcm+ijtliDAJAUbUVZwTBjobzI5/pN1eyhzI+kQc42uoz2WeImC0T5nt97B9VM9
hkcJHnHgTAYQwhHQaJvBmgd/bncemGub2yh886J+cBaxppH3tvkg5Q6XemzyQXnn5vCBTKs1e/Qm
TkMHYMB5KMpqUrnQ0fe6zlVWLOrgIEXED7sPa9VRHnO107dXNO6ZxgqUfd8/wOX1Q7Tn+KesSaK6
asu2zIN6ab0+lDxrinnN+7sL7RKNvCB06mklgY5u7exsX1oMzFJ03miJ6wh8Zekprm7MwNqrtMf+
DLlEcpGJvyks7p59OWEpsm5wdy9ZTvUC0fzZBDXn9sYFY2SuQ7tgDUxDLzwPCGACX79SYSh9vT18
tlwHbhtF3BO+YJEQ/f2OIMW0M4lZPCpMTn38mC4l5KCQsae4RxbanHTvaGC9Wl0PAx0sVgvm6Tsu
ujG5SrWiCtnm9BWhSHoNI19aNwQn7ly7CUrJAoqjHheuBWC+Bl7hQT2qqqLD51/BWtxOE55I4brz
8qDuh2mY8gqlTx+N9Sify3qL5La5Cz0KoK++x9DtkTluVMBb8RGiNgR0nppVyvOJDBLVUr1FA+34
6ypIag7JpZUFFy2+T+3xNHiQZA5LUP69NjRIstZK611vX2Kd6RvZwifSNR/lqpCaHS8rIhe6ew8U
4cOQgpCGB6BPMzgOrkimj3WvVTxXivprhNW01GMHXH+YCy9cN49dv3eIdLC3i9avm0b4On4yehEG
mTc8YPejvBAKlghUqNz5pHtlBJRefnDRT49rTQWYhjxC9VF0hyFAcV5Hu7HpuEWA2r/OdSQQqQ+J
j/db91ESTa3fbBVVxHEh/llaK0zmDz0KEyoBmt+8pA+tUGRmp8j+wpx4KeU8dbcP/3/vQtfIn8mg
2c5QWMtUgp2UpnkM1xMV3IHbOqr68JV+Dbn2FIKYrVlDS1/stVZ4dEq08cRZ75Vqs7foNVqXwOCF
bBZJt6hCoX4D+2fPCQGygT4VbVrSyJsivdXE9Bd4Uo/bp0QsTsGkoZwPlCwv775cSQR3AVbgsxlm
92yR1PDX3tH1UbcX3Me5UiSxIqznsi5DuEbuyfDX1SWXuslsPxritrum9akiGq4+NDFs6UbIGgfR
uPUb0mVjiJW7eFVl2U81Og9Meoqjn1oAj10yiY7ouwjo9Fhzb8N4gPVoegUdalumhmE+aeVwqQwZ
C+DVxaPzu+lb7Z0DvcK+a101NishtiWcj8MXgCFnkNg481tw+y61v1IusC9WDU19EIIniOd+P7Jf
0/jjfmqScq9N6HJHqMWP3HF0wJ3zFDx5gf8EtNaN/YYHRN3j5Wl9BbmzrtheNfZkYw7S1gB90QYF
OHDrSH0RwzLpwBgHZOjlDy6P99wlEVM96b+oY838QiK2HGKLthMkcxU/SKlafzo+2fDdLbqPGtVP
GJnjXXGOip6ZJQf83XNa3QlehEf+a0YXqHEJOifqEhROF5j/fmUkRalyCD0AATnTBJEx18P4p4ei
haVp3eA95nEQoA5BhK3hgiRjuB42ZPmJSIBj9AvKsS+Vi/fi/MOF5iRrWJp1ns4unz6HxztWwx56
GLvyhmjAg8gcW3fAPGSrME/83YtDRU573waL00R6StkaE0n1S1VFwOrpmyE7re4GRiGacXT57jur
BdRW5ZZQa2ouWsdQWKJjIF2bU0tc2YwKMkyl9v6epa3G2QcXymXEw3NHN1IGJnja9H+16+6WkpWU
pX/SxbsLR9xBvvfABu5dSYkB7N4pBaGzMj8RIs0fHtkWvFfC3tDUn1Z5ESWNH4yIbypUK6kNQKEa
Y+RaGzh6GiO0mIi7m3ad0W8nU4QkmBH5GVTjISBsIzWVKKGmyRzT818E0fYpDtR8OsCVFdI71t8j
2hgffP9A9MHpTAOlJL4lZTjZYMygg2oaDZ1AKaji6EHRVXE3qk605dt6C6B6mFhdNtHadv6c5fIy
7XHB28Hc012lF8ynpEbsFza7uO7jJbTSHTGrVzf4p1qanOafwjGecbG4WkWw1h4/Iiwe+L55XNLO
36n5MY1B+gDzNbbIiE0fB+Pdv5dCIyR0ZIq+77RyRnqYRzIOmmBlvjgcGSzELFoyV29C6L0Ev25f
fQfxS8/C7jNLX0nHMYxGw/U1Kj+uzrTuJjlLo0f6GYV9RT27gWccLoelj/dDjjcVUQzJe9AJBBbo
j1VEVSJkj6c8+wNn9jvmBN/dwz600eQDYoItJl+ObBH4il02wLA5PsUoV9NhoyMo6yDNdp4W/vSY
aGZqIWheITRKL/BOMZH8cYPLMVVpJ6b8f4AaCwuxo09J4sufvaN98U1xOKCJgpJLj4LvwoS0ii5x
/ekAJRil8dF5XY88EDr86lUb9B2NoNa4y4Ck20DtO1C3IIS6U2ug8QTAmXy6/gFnlPU2j5TM1UTy
Stfs1fGwTb+ybtZPFzdvvQGNpwapVQydlQwqoKMQAT5i7pgnOTL+g0G4p2UpOg0+xNgDQP4A4o3w
jMc14gRmf/rR+7hSLSWxkdqWZlUtwdO4Ksq3dbMT61XDshTEpaVRZv3zceAfwLn/uPiGaI4Hr8ZW
e/oLcZGwVj44CZgtNKaTML/pvGP9cjyfQeZ1zH0oWaBcc74bXl7X7F7NxqIejF7d4LIY/Bo3PRZx
ZLvxCYyKvxy6p7yB6pbvawFSidBg2H+j8umpUYkQ61ZDKNYSC+QgMiSqXlEcTDkFeJzveL3kaqcR
aMC4OaX8hctK+67ZQwarVx6zaGgbcSAhf1F4OPYhH2R2rjUOUp1PmFPO+8MU+OA8UyvE7+gTUvJH
9Lfo183A7YbSOZNVzxFJLmlXMBhVAvDaTHKAUg/tj6JDndTgflpwmTpSbe203vovq5yRUna12V8X
+sF/A7Qsm+Ih3zSBbCTG42w5yXn7in8nfsamagjVTvXkg6xsJg1ctntkb7eVjgTr3yKMSrJRp60O
osoZlVsXi2ncBGxlhAL9WStJgECawiWw5IMvPyoUQBJgxTxsC+R630UdWY3fWuR0ZV0eYOVV7xuI
hp+X97P8G3SQ5yccutbTyDAyMn/OzaML5jpHaModziux2mW9GbMgZdR12WKH1EaBBAxsSbbmduvh
N1teVgvkzo9SPlHY4j3gMewl8QgDijhgBTOydNHTGLu3v0ETjkDEqe9m9jHpXT7K3s2ERzb3u9p2
79Ecq0XyU2zqnqn+Tjjv+hxm4UahFRs/PPrNU9PuORVzQukR7f6+PmBRfk3UZrwjCjGn5ClCuKxj
gQNW5lo6WldhKzUcGa4vBylshWt+G0kXpC5flI5bCiA4Yi1U0uuc3h0ktPriaFo3AdrrRN2FyR76
8jqaYUZI7wGPTne04PNxRBcFkQZJKKmfY6CeGfg9oMQS8rq53Pc2zVqkgwt3VwpbpwECU5C6MZdu
wGigv4EczjqWPhzQSnOlOOKjfdn+5kpifyVAOBkyBNKYI3dvFPotVtcsK53vsTdRn95qQsLsRAKV
n26LxhGB7RY9/l/RYKjBQSTldCwa8BO6yNPSgwD969xupQ2GEmiroAcnM9eFKXK63sKYhMgiNVXd
9qIUzJFBLuNzS8iORNManr1Ed9+uYnUPwM9nrrt5Zh9pFzdZ2zyebr04xrgU3kz9yFsfVyoJE4l6
qrmemCV8Kahqu8Nv9kNFaiKejXK7l8QpxzIW5x52iBnh56ZkBVgrAIfoALh6nHK5rfN7t9Bt+6GU
ftCBxFgQ+VRlGs20Y/KFXXg2hHupkxdaqiLf6UXhaUEN29/1cHFIA3JSn6V2aihCpG9FVZhVUvXf
5LnbLNbCE7+B0JZdWCacX1fNB7rWTMmTDcnwJgNYZMykMoKOuQ4nBAldcY5aSGZEDKcQNuNMeRCo
f3+LCq9ilCGS2E9L9iaX1FubZdB++LKJIEP0eZ7ATrjIp5VmI7x51ctSW5sB93dhSllTQ32kfeaq
BkWNGMsD2Ypn+Rvs3WFbjeEBzX9V35GNDyaAq1R6ofXjsiKJN85GTug2zqYX9LQdT8pmWwgb8kcP
BSvulZIThQZBb652b6ohSkP9ob5YPk8H/o6N2S3C/Daw4ggezQk3KfnGnEd1dBEbjuoC8QNKah1U
EdFcCwG+uzh0vFJUbaG3iQaN3yCXU72LY8o4LaQ+/NPEe4vxBmXJSSskCR/oy7Uroy2Dpefo4N/F
1TSOx6VZC5LmFkpzsvt05Dxc7crlLUEQedZGiLN0j1kOR+4hup8RpS8QP/5YVUjozKrYze4an2bk
X2BcCB+H7cQsFGlsXpK8xqSB/wDJg2MnRWtStnLSHEEl9zSS/rrUTFKPEC8Jl6bQzJFkVYpeFPmc
jThRs89sDSH9x2ytyoJESjUYZu48dyHLwfnOE1d/x0NbtnAI++cvdt/1YAtsvR0mSFLSW8YXmb9z
ZNKHw56jQ5HY7kDsbOqOt/ltjnoVGL2/sM42bD+kIPB1WMQkeefbbp+R9ugcj5p/RhM77Omh341e
sA2/0KOaDHJSVNFp59xJkGEQYMTZ55+6xXFOTXf0yMxouMugMjd26ZgHcvkBcJOvD9tl6qsICH1X
4l6m+9EkdMyD5GejYsAQqAWy1RGPSYckFs1WKur/F07E8bI6RmBr0Jly7mfIoULcA7APSkDPNveT
4jau0s3i5Im1XB7fSmX6szefmjvRvbfLiuzxvYB739kEarci1PsEZZAKAIbB8HahjVR5qJ79iDFY
pm+HXF0ZgUIXMi7X4ArnN74gcY7Sj35a4lGETg7uWhwjeNmii2+xTB/9a/WSm1t4xyHQ7OrSYzbP
rHSWGt6wlz9WgdaWZyNoarioAcn1nfduOkEXv2v33XdCLjmwROsT3gymTubP2il0O5wTQHevJMLn
k2W/iUxfDJ8PCdL00QI+bEzsiKdsxIJbvQ4FNnSlvHnmW8PyCK5VecFjmy0xWfkhn132yTp+B02A
Y1SgmjeKa1Z2d4oofloYOLu/QIHSfRxYb1QNzXH9qac001N+2WRDxKAFoxjmW9uH2Dico2ljMlqf
U1yNzGNQrPXaIbLYY9QburGrPVAr2tunc+1aVuhw3JYJSrvLKKfOsLQGjVEY6Y7XBEfnk57dJl6K
9EK5oNBjgUxrCy7aHqOwm/IGPLJnkscU9vZcQTgFKDW+vviEWasVQ63TMHI6tk9epkAxIAE4fNwK
CR1ECeoWpUPFQNTXMoDr/538W5I+kGiMq8weiximO3Y7B7aGiK9cFnkqECAx3n/fpUczz1nP6pAe
Y9TC4S213tlQwecuV8632LixIG6wbXTVnklBBEfrBYjPH6K81zn5T2sfgOVeSLejIAPpSzay1gkc
XoKx08YZxKEnW9ZJV7U2y+mJJMfCR7Opc3/eA5YtrjZphnMtHPsItUj7JkiimdPEI8CuOV3myrzV
vqVg+WnuiuAPOKCgIjYEUMq5kj3STSeVppbAiuDLLiIIGX0/eiubFFNonwxSC0dQGVUggco+jcWj
wudUoJ5sAzxwFXkxOB8UqFehTk7sw0vuC8w319LF2zM2jqBSYmJamB7OmPZt9//ZvsDUftWtnctu
tG1s9Wp34Xc+g6NEHmhnIfRPr9v7ciPO8V1p0H15ayxLGdftGxZMtjGFSByUY+7EhlbrxhXbnArL
IgxRmopzqTXK23bDpx7VV19EF2q2vv1258k2/nR6LQAaG4GnMuQ9zjX3IoBVbHvCkan+ppxQUSUQ
Hd0kWjZLD6SpFeLtQmwN06ZRIqdBnKrqtIHWIiNunWFs1muzOOkcBv+Fu5kPNFcqGw28HIJGMtWG
z11L2Npkjuz43YiA1mxQsJhIOfJv+zBd9cKjtJI3IrP5jhR29K6kV2lGDHC1Rh7aPfs6yC6HJ/86
fCgAXbgXC+RMiMCj+Js5VGJAnhJfoNXeMfg8a8A+hRmrwejKIaMvI9re2Gd8s5x+i5JX05FGJnP5
badbFxVX0hziWXZp1mFju5BG00nnjx3/ImVufBPGf+2tQiLDSCsfUdxFbF8wIYJ7E0rqoTGxJ0uV
L7Octyd/+XZvgUfJu4CoivBvJbVW2e5UGkrGuNkoxWbH6jg0/o9YDP58+y61d9AdR8noHAC8zRMr
VBCCB1EfryQfRXWmw3cFXqCRsC88Gxu73etpoffKV95AdijEPnt/ugACvcdrStYpwfjOiC0p0FhN
O4dyVTKHLO/ogcjrD2PR2B+JfaulYWNgJXgD1JhY9Ba74WnKVbt0pT7wqOVsJtYFLi+9XpuH474E
x5gyeCa1i7EQcO40GPEJGENOZg9NuKIi9VE+wUfWh3XLlftel761QvibPq+OojeDkWl7kwf8pUC4
YG2duopkE5jIit3X5/wvwC3dt3Hif7OPJOFrp3LUb68oUOitHFSisqScHgnvzRlaomnd+m7JTCic
dvvAmfGsqJNhlyJa1glFMLKMWh5kajzJpR3AF4lH+WLO2yt6zdBDDAKz+1+ss18jvJPsvQmE5/of
ldhKwgPlcmcY4RWEcA56N4e0DX464XOnMnu9jB0zAxz15No9DBHAmPsVgql4WdhZYO4hcqHqlzFv
0o2iTbaIVCUSg+pdVsPK1KF2cIiI/32kyOC89GBkigXt/rxB+xDMj08gK4mdTzz2zz4g4vmNqOTm
2d/lkOI5SMrAhu+Wdgh+UopD3SbX6LFy5jccTMD3ONc+mgPWmy/SzQ7xOWC3wid9d2yf9b+Y9oaA
Xk0IFfxQxDO26TY3fQuFH7iWf21JHeGswkNWICbTm0jk3cKsbAMCl0H9dKPbHlgqFswW7ZSKgbIU
IBpqui4anxji+TIu3+ZrtcaFtHIKnj4+pXJil6itu+UL5t12sZAJGujLM2sM5XXmjnojUe03VdFU
eIHEjGxKZsnJr9xtRgC69iuSxUv6RAeyPuC/DWWa12tCmg3dvF4iIwGVVvRiZORbgeUMMj47VrLG
pjadKFBUtT4KRw/s8vqKNxn+iuoPXWAEoyGeqJWorzLayyX622hkpHxeGkp0p5Zqscfsh8tieQB9
zGG4Cu8d/Y1kuoDO7ZOFtPBZTF0/7hqWJdvb+aSV3zZQuVC0RUhSptuW5yvWgf6twrDcZp8bFUHv
itw9eFCjKTrszKWqVy9LAr0/zXWm9QSI9qiV7rlXBGW0gsYUpms5D3W7YvQCKgw5hmjMhjCKQNSo
5s8UXQR/z2HMDmHlE5tBNo6q4AMErkcaB8dgdB5231qdhNzsfvPaH6caj0ntKP8mcfTNCA4PUIU2
46mcRzMvS2y+83pgSY8LXHKO8gjsNAGK7n54ga/+3Iw8AHyTbSs4u1hn01C10igd3poX3OWJ5nJP
kdzKbwznMVAG9tl+Ztrk05S7c7hJJUaTI8pxil9G2NfXkVsQHTuOi1E35vE/uSnGtXNrEbLM4O4G
CNR/zsTEbC4EpqoxOcbgaoLh3yeuTjHualbjb57xHu/oWQL53IT99mN2smnWv/iWdW/jiaGQ8nuM
Qjhg2tAmZiPzkrlWrv/BBMo0Roj0OMfLDW0zkxIFb64uejoHLyPzSx4n6o2YuU1xQvsx74QcJdzN
d5efa3KWtuUiplWvZZN+hj50Jxeww28IjVV4no4uokxPKAxNUJMYOfDItCc3wyETKk26onY45iSa
VABK8+bqnEONXkMGEjDLygr9V58s17R5P6cm/oMGy/JS4oJxYsZW30+BDd/l5l4SRvrpQ0nsgOBP
4ubaprJT874LSYQHCROKfyTsvTRx/JIlL7GkHE85t0uPNJiC4rcWoZvmkYhfhZNgI2RvcjgEHv7D
FXWrTbvvsaVSpQSWFT8qfaQlMadLv/4ekOxkFjQWO2cAzmwZNs+Jdzll5CT2/hc3IKEExc5MDhD7
pkak3S0NXqAJP/zJzb9q8I3ZJilrqhG6yqqpKkVXv1ch2Q4hHbjHrMWZFbKsbyIva2prKTMYkAuo
XPpl/sScVRlKst6z758fXPw7aPPH+IOjVzjXVWI1UKLHPk01g4ajkdec1Kh2N592QYrHrQwq2vgr
X6pFw1dFsPIqYuE4x0f1IZ0VCuDpfN+N9eM0N+dzpJp7mIXNPVmaRJ+kHb+/TLbt87RYfdPtwuQi
IVBWAxaYwXh96P0/zsN4EK6AUYEnCvj6BKzRmccePR7+XvY2hZNym/cWgci0aKxp7957+xSpyEEi
eRqBvJ3uQpB9h7YzfqJz4FmuvoikF0ZKBQEZqIiBCDf9GABPDnMzyrZuJHwXbLXnAVgNWb7TzGST
SYioU+y6s9OjpDzEEZkCiFRfJMSEdUA6jmZuo+LTdB6Bhkf4xKp6P5dFYeqjgnoFANQkG0vr/6x5
uuojye1JNjtnSqj8KMTLxb3v6XNkJ0wZurJvBayaVuDbPJotHlWb+M3/V5fZSqRaCU3VVqVH3UuT
9nSpoiIrVm0Iav7ll8wRP2njO3slKzwAOrhQaXL+Udp8oyr93+zb529pGvXkOPmtihxb8Z2yenKp
1aV3w7H83uurPdMSwXaDNT/h1EayIAtpFj5wuO+TxJw3CFYtf8DgLt8li3z6wGUGi3zvcDD7WSQ4
vGm7U+TB7V7VQ7Ogssl10lJA9MmzBECt+v+kJNFpPQaQg6TvnDTPpGAH8XkWgkJZrtgzzZE2CpZa
KPtafyXOgr4iZakaG96PS86AOBGKMBZZYVQ/FAxT4/sW0+BUSbHnmRfTC8IvYOt5KlW5oILKYdx9
57hOPFAcsWepvBbhxtVlD+TGVNlpGFCp5ZwvX8zrUdeQGMPc+JgQOOU3eszI2PFlEuuGyOmLVG9v
j3hMzsptRjKW5KMIASwtnOYvqnZHAx70ucZnsZrgESRVD89Yq/XVidw0Thyo1R2NrfqtDk0KahRU
G9Owpc5xo8AbhuBJ59dFS4ArbodZ50NcvIlvUKpQjxRcMxiymIKC2Ekl9ag1tXWKqx+bhJ5s38jq
nwuoAbP1FDP6LdQwJpwhehiogSD/RURgdo2vhYiCIG3CueHETP8ACsRgxIIpZ3z4+CclkUr+Ck1F
9Km7ioQGwPJm+pgsUX+2ul4ozNjqsQK9lopvRJqiuVyBo3SD2EpyHygFRoGjS9nLWh75JeJWKD1n
JovIRLnqdnTkrEXwNgwK45v7MXvIe1Wy4sBhAdW16v+pH6KEGU6XLhIFjN/PAc6bhMIXvbMLZIc1
cQIH1HHCSOVaROqqwGxxWwBDqZdwpIozXsL54MwhuKCQLTxVSVwDn0YyF/fZC7RP4am8BNIjgXpQ
rW2DKZkGNlo+o/iaITPFUluL699OEQPVXsofdlLwc1E//AU+mUkAD3E5Ih4rRELUc8J1f2cPO6DE
5L6czmHlT9TpwU8eZZcIIL9HDedE1vrxrCC6NpcjzG//j7SR8sOft5iagCpmglIONhydbm7HnfVM
66tq2WCgIFBq5AvktXQfqXgueFVzm2C1pAa5MKTPSexP5XJvKV1NJTwkwgyT0jI5YpXRHTlT9miL
Ysex759VkYmwmg3Aw+ZyRi78XpVkzj9ZKsIlDco/SZ5wPDbkKdLi3Y/Hh+XT/vAFGpHsd5O4Xw2K
C6ko+qddtkLl/TyMWD+530s5tEKk6skn2g4Hs9TAAlOWxbK0iY67I78/4gbrgLQWzEwO4RBQg2u7
XSqNqDQvJZazpfQlAMKlhbfstlh5KYbsVWXzAWaBO/kHsUBldKs+zl+pgr3rjsc6pA+I14j79TlS
2F/hC7E70cUba81bwcJkf8Zee4iPQ6uPsyz98Qbdz1nx+GgN+0ejlm96GKCEzH9HwG02ThTnNFZd
aUY0M2Rn+v1Rh31oTFfGisi8ejWQnFGb4iRqNykM4rS5lK5ka2WsGWB6B6xcBdWv3Na3u3VlqEgj
67P+JwNMB4pL8n1ks0i8sXId4ft01vKek4vnITIydMqh4qh63EfHzC0bxkh+sN5r1/SXqneUM+uT
EMB9CRBDaR5EfRii+UqF1SZoDpxcJubABGhnvFOWqERUUn4hFQJajHevfpBLkTE8rmZaSJzAJ+pw
J8qvek3eAPneCKtxGHjulC6hxA0HkkoNqR6Qv++GQbMP6Mlp/SUHDaFJH8qsgIPMqkp5mdV/ibzA
ue4uMHrWmzuVw4IGYGeudatK9ndXq0n9otS9xMyRHfd71jVLn0PM69oIiSxm7/8Lo7bp7Z/Cbpxp
ldC/YwJL8QAX+elFBTX8x1x9K0FqtuzCu2UPyv7llBchKozANW+kYKgved8GpBbxXcJ0jx49SICy
Z1C170dAkHR4mZTc7MwR5gWOHYmt93nPHvTa+Vb99wn8aFJXi1vwd9DIqkn7hB/XVHODfFr+qSqi
fRgW+B67jr/4N9Tuge+fHHVS0d//EEjvRcChe2s1hNTqnQv3axowAdJ/QcRRHmIDvyDOoa4G8nGg
IWlG8PCHWEKK9ixYv2bmpElFIceuAbJ5iN28bim51eMYLGd+NqmQ+DQGXCStiYXCAWRX9wSYa9qE
518HPUYVU8X/VtUWwfPORHwUBYGMxy7y2u3j6vN3UOB9irWnC4SRAcBay9Y54GvSfzR8/BEOAPdt
uw3cABjcoD+4WFL5M5M5RbZuQ+Ab5To3nOsKct02e/sESVXwtH3aDUDdJwoeBTTUpuB0R6Sq16hA
uShXLYqy+gSt5aRTvrqH0drVXTaK8i36R6+lUaa5g7WeL7eoY13agTCdeljJAMjN618dS4oupj8O
5jmQIaLSM8b5nSEkMA/H26aHrwunt9ivUcNMKa0AryEb8rWoT4bn2+qknVlUeNIrN/GQcdvAEMCs
u7YkoHW6ghs7OiKDgVg8VZefa9JnBbmKBfG3HKizfNExcRi9XyV5+O+cENnCBMXnPNyJoj1FNJ88
50fk6l3veoceQPbamxqQgb6w9aZ0XK9uqdn0Hoa1fY8ZlsrHgtL2mv4WgUFZTPScd7lfJsc8+r4A
BDfIg6McNlFZ0KxPntUsKgraktG8ZHk/gpayLK1Vjroua0b3YjSl89lU5VN1M3r3/rfJ4ZuGWKk5
I6qjB6Tx3FoREvirCmMFKfsEjw3N0htyr7TQnB3OpsJgbtnmC+4nDGWMGMYEii10jMiTA+YU6pBj
RTxgmaKOXKiey/WzJ0D1Zc/pBrzao0k7JxXyz8JrZLjRV4oPbj2fvZFMoscLEkVT0BpXjcyiYiyi
ixm6DhZBBgQmxjttKTz/GD9s2xDGZgVa6gxv61cKVdsoHhtpN6s+GNc0CGhDPJjB4+DFIUErdA/k
h82VieyeldwpojR+rf1eH7Pk8NwZtwU81JTuf+YjBhcdtiw1qbljZQFqQEbYjEbQ6CODWQx2zkKa
NbIYVC/1ci+Ekcmty6cROu+/mwXNfF8W8PwBTIvD4fDuwdpp0CigtT4rPpe+8Nr6Dtld4UqadFFx
xlkN2aQVZQYhKSaDFPB5MKqUOurxKQ/zLa5hftqz7HUTsJyWUjxIGzww8LQ5GWZ9ji+y2hNbTwpc
kgbRrNH2+UbdcRbBwQKTQLjpSaraYC/dSvqfLWxiTjaYzZiScb/4bKmqiIyg1LorWpefA3yECcJ/
JNPHBlMdFHWN60cPPzQl/vmbhFrPmDHHyMKIwnYRgt0MlV8bLfzUcNW0H7IlTc5VkzcZzudWnUEH
EpG2ViWgP8nIgEs0xwPVKZXP2Q+A4W2rJxfsfsaECfvggccSNVEQBzMSDo6M96hurm7BEKJ6NBSa
FtxjbXPt4AfB1zCLJbyiFS/X/L8uXIgsmbv2KbParmjwmHSVh0SEcvGVz7d95fMXMWBkbbdXn50F
HcJA6o2VSTO0GpXtGFqrx79gUp234M9d63oTwk9B7g1lQz0L1LVn7qns7GPhmz3Iut8c2P6eKaRm
MS3W7hneN63jYwUGzQjKIQO/omXc1I8jDQGgUPzuTMDLisU5pmA1VBYJA/IaO4Zei2QEsZB3nMkW
KcCo6PeKB3aznxg6R4DvAlxYHs3RrxRLb1bgTSlo1yLUs0L2auN/esM4jcbEKbgvaLtFP+8zqkZW
+tWmgD5KEay5B7hL8mkYKwwcZfCOUyokopO2YfJt23lqmOQ0V/gQoF3cS+bn5tErWWKiWhgX0bk6
Pa8a7KWDvCSwpo601J3vtT7SjKRAz68dCv7Hhr4swF5niIrvauOYJBX+S0luq/dZ9W5b57gvrF5p
Ad5PXJjLvzhXaF68R8ktD0n0Zn7RBcwtz0lPLw7uwb0ra0t2mIpaRtGwpCsgjNU2VMXBNOI0Zw2Y
S9CHN1zVGzQjX9wx9XE4rkm2WTkYfkjM4fKT2kzD6xP+WonQQTu8DYW4eavtHP/6ogqe5vUB62oA
gz7LMFfARbjO5J/t3XU60Oh5cBAx6nLUxqDhd2V8GyYM+Phqk8P1VIpUnBjoF+qceWT5qqArRUcs
GN1R/bf9mMULsca/wFZqiVSM7VQl3avT+dADaAW++Gb/LDxaxUTDt99+ftxAa9TXvknRWioAiDkH
bRxYVQUm+UG0HjjWLpuduY7mrhA0E1uIFZB3MKWUG88jdob0X54rvTQe3c8gaSSCxesz0KC/IIZm
f7ZNM4W/z+d2ftHhWPMAJ5/t/u45Bhpq8Siky+RC5g+DZzKayEIRYbKLhpHE7IsPFjbkGC0p/UXM
N1Q3PLmZGphYgvpy9bgWZacaqCefZdfhFUg3XSa15xYTlOhI2JV+f/WVoJIP6xOnheEa8YKc3sWF
bO7lOmmgrmvxTizJJ+LcInXX7WnWlKjHobLTQz4uAGXjJtTgJ3/VA+67h6iGxnoRd7jkz0oQ2Cza
/r6uHsvc5bN8nFai9iZmhX9A5yICo3cluKlGl2JvjTgFc2LfnVsLAiaR1Q/0XHYbJggycVESA+vk
l7NrsrJLFi4oD0l5gYq/Jr2t1ImAzZnr1fXoEZR9vr7k0yXvT4sYSdaUIQmbiw+/GUya1cCVw+YZ
csBTaflE6wqFFR7DMTbx60MYHP4O+hw492Cyhb9NXW59Icpb33qMN17VKZMX4MoDue+PeW6f8RJI
tWtMPDWDpE8q67vmeHp5/0ksPuXoIVENze3iSQo9CGR8MkavD+3WoIgIUMJtOL3xnHJ5o9kadeQN
0e0s8xRIdwslWnrtCNhniYms/IQF2+y7PcbQoTKzNVEncVRe8kX+p8tIqUQmVgZddgwriM24FS4c
oncJykXHR48TmkCCvtxytGl3mMGTAMPgx1twzZKr1A41rbk9JcAbZZH4PvxgBPJrDlyoFHcAeV6e
EjD9LRuFO0xubbjHadjVozw8cWjOUMkrq4ziVUYBDKVKWgc7AZefL9rY1gM9KfTQZl9wCCx+lSp5
9J+f9yHcvbuBhBsKzOgy0aVQR7NN6xIue9QS2nLCFzw2Ksl/J2yqnGKAv2rJ0akD/j9Yyfg2gZd0
TAcIbV9OmI/SE2NGMWitF33iysYpHaynGI1SHKYpm8voxb9FWWfaXcnwuUCIAUyQy2JfFNDyC7bN
AxVQTi2PWRk96EVpI52x2ZksJh9m2tuCY9aYJeOoTiF/XyGLXrMgOJQLpZ18m9EPLNDUrQXL9/BE
7WHD1QbzqeIV07oHPulkn3Lk1C1vVJWX+OHP+gPJw7he7iTcPvtK7PtZ4EhI7KJDZNc0l0a0nYtP
ekvG5ewvt4yOxDKXpFAoihtdmI934QJhM7zuPNwQKKxWm/di3lIV7V+lx+dQdo/3uGbJZnG1OCJJ
BK28aepR/qJSCjfRGX/eMvgkLvVintlK7F0P3tEYN/6g24QaYzBgCHQy5YY66cdn/XwJfXx0La1j
uCd/v3ERqTjE/jk6tw7CW7eESP/j4zpGLDNqM4VLmQiH0c78JWkto68vND7/AW04yES6pZRoxkJh
FmtF4asmouCUZ6pAIK2hVOQH+t6ZJ22rHFl92dS5vnKPvXc0yLFn7MAWKw0YQaoOEtDa0mjkQ9Hi
QNHWRou/CpU56nR1yDyFVAo73YcCFgYXZ89XEsrovIEBixRTzuSKnTcCNU8OyVc1p3XzvuGP1IjG
jNMRkUVzxLZ5E4S4+6RNMAeW/2RtoRsXU9zeojpJURhXlRW+Yla63Ln0yOF+prmGrB0tcoOLL2A0
v1zYzTIixWzIrwDQL3yUZTYYJCb5bmnaCEmP08ttGoexav1v/yoTex2VfNesUyE3PjEr7i2zW7j+
tRatch172Cd+m84wR+SyJLw+jijFHtko+p4pEV0xXyotOSUhJ7hgsaq/ZTWDLqUWd5QRj7NOdbcs
wwdwETJ7g50gLvNPwMQX5hl5cC3zgyAMaqoklc0ASSgF076FhEGIGrEiMb/By0KLUbn14PcJNfqW
obBagqD21dgbw8b6EhDppkelF7gC0ElF5hN2FYLqP1flt4LvlBR+ucdLU+B59qm5c+cij/adh5vs
6kieWY6yL+YSTH8qaLSH8cTxHflRkiut7eGz4F6ZAyW+mO0NyRPDLQNFx76/wP1MsKEAL3uKDjXV
VOa3/O+OGmlfUsAbW0yO4mQUy8uUWRr664hIgM7JunqXWrQe6sPJ0kyhW1AjR5PSpQsJyBNKkcf4
GVvAY+YBPjTE+bkKu5rBHwJFQ6P1asWM1l1va3sq0F32Edra9sZTYBR8Cgtas5dW662FDKLUklMj
djW3j4m2SipTWpaTC2bVcO09cFAFJxi/hmsVor1Z1PjoVXwqLSdfgZWroHvmOuBiqJgdcXu4PawY
h1Qp6cuYtARcFY+YYt1n+x1f1Z6qWzMXAZ1UYmxUdwNUNO69zLLw3BxO00HVfGVkEQRnwkeAFi62
e1SCgsoGyCr/RnSMQ+a/ICXJzdx/QS66aEGxkU4TlHcXTENCqQ4BQpCeXYvSGVApR4fN0W8jtynp
1P1tJbtIAfnv/a/PuRkYi/6SgJalsGBv4Am1YoxY4NaveDvpJcv1JTIf8MGdG/U/xA7131YOY0HX
Ept6wtbWyyhQgU0eIZ2FduAR2+E5TAm1qXLpgoMEEeqyS6lWOpeTkXK9MQILbzaJoppomYQ8qlL6
fH8VNFzNmLdjvjuUa+oI+6Vh+NXZPBLBecB8kPXx/OBgsTFQPwwrKD4D2U6YUN2ERgCNghcFw+6j
D+H8qnXV3plEzA+DwQgXQz4x5Iej25j8h1Jp0DH7rtb6krDmAwSXh1lLMSic0JJGR13EzBqRncS/
650yHELqMdSpwTE2W5T7al2dwfeRrjU9PrYB/fDTFmzZOJ2Z+JkUwTrVBRaJMmilPWOUVwG6wd3+
MUbgIFt0WaWahAj+zngjGVL6HHnf6XaKOG2BOCWW7yFYKw8+jgkBMwk0aYBPibe1p7pJzWM9Oz2/
sRCTDR9PXpIGLJFxBXnLANpiAjrotAKF6wB3dHlqNhulZLUQhTKSi7e2Xe7Es+HaxvWJECuX9sWt
LTHV62GqZYJmBtYOaA7ReR872EagkHvddTsWVSj37smnlbsic77U+EjKJYLDZAFzhIexqP3V4iHI
VRVOYNyaacdbD+du7aLfumw/QXAsmC5OM24In9bjoB1lBzwm5AWzNLJexJffmqTBmvQf3oY46fcC
gADg0YXl9Vznoo1/oZtYWWBMkO7KnIIA1tiGUUFQlV/zV18leBY4t2tDW5VXxZdcTXmjam6zwkUk
uH2sN4ZUP4hd66zedLiPGMp89PB3geVs9SexHuQVuqWZYnt/K8BAdMWNdxFtZBlhJUJeVnFDeKVA
WXxj1rc8VEMtl3LVFiy7p6Q68G4gh+BdsX0MYXa1wnOi/EnVg5x63U8sv9l722iPTJS+IH1GW4nE
b7j9ojv7VXcNOgacuBfEgDai+50qNWqpS8VNPAo8TsJiZFe4NzznEhBohtYO+uD8AcjYYomzMolk
eSrhI3m790Ub6dTMeNpbADGHag+nMMO+CxWPODh4RXc8B8MVGg3RRX6Ci0XT81I8TMXkZJEJNAH7
sIWq3ivtvOkIfiqgONjSsCju1QHH5SLGiA6t/kNa8SbasbbR43W4pX49KrYQD6WYXDbNtqtWMfRj
B2OrWzksHOlRIc4boCkh2jZadDfz612yimrE576z1IXA0P2MtFaOdqq2iWPr2oxb6/+kAzsVthH/
hm5SOYuMGjtGdW/RbXXxyxBPUXMlY59losQVKzGAXRcBmgffGOuarEPz9GPAO2mtERq/lqBiigVZ
o8vVO+DjO6rfE+u/t1GrtVbMJ3C5FdZdpkxRQtzNE7mX5yl8tTgYqwZAlUdPOcms4G1SA2hh8eei
tT8WHyA9tDKN+UgAvvfbQZOcikSGq4uWqklRKDn3QK6F8UFFRwRa6gOfiVzJjpFEuxr8OceX5qBH
UJV94wUPUtdu/bDgHBiIV6swntwm3I201DS21YWe7Ni5G01ewi5IcGmO0Og0y128i/YbkP7jDDtU
f7C7Oh1ec6Ks4jtabGWPeoCRSDy5psvAUvU/ic8YFAQVmrHo3fDguQHrD068sUp8Izk9Lq9/52oy
jWHYjK9B3mc7gxwl+caSKEwjuyw6db4ShJsxI0qzkExvCraKPSvhthf48PMzxUUDbRLgwb1PWulw
2FExgZjOq+3p7+MVApN57cTJj86g2PchNBRZsf2+2K/+oA3LH+Qw32EJkGXUBgHTnJDUM1Bk7FZF
oaffgf5SivOunRTDmk3iHAF73WoEYNl+qVoQYZMWFoRpX1W2Wg4nq+rH84grMc/KTMhNsTPWY/O0
VkZHkVak2rSxKePD50f49IRZWzGQ8C6UaSQjNQrZfIkcHvKok8PeCMC2LgsC4ruW96UA58bUWj4Z
7rTodXtPvnuhOB0d4XLYWPtkJzitvygKswG5XMhv6QEpCJvgj/EsDDjG8uM0/rihB/qvFZegRMzF
Hr9RDYR4KuTapsdjVRdTCOeVSOUtHbieSJHgTwbq2E07YoOUdIPnZlL3+NZkpHlE9A2kJ3bBeFvA
a6WNqm5hUOdCP+S0s1XUgkEQQxqveIAx8An7cIZQPXcmKBWzUDpneC4bQfhg4vVeht9X15zAlcdu
kMyWlzE/pFV22u9Zqocm+UiQK+tZWJVZ3lidT0tL5xU/06vjz5/roCKlHRzPTT+MWCIcHjdEom8l
5AT4IHwkQs8O+GqQ1H3A8t8qQ0nUvtvjPp3++SEaLqdosMG4QKtFnfca7TePRjtOSzpC2cLaECnT
94tL5h4AoTPZZKUlAvjdrTbzYeqtwGFuy6hy9uVqE0gCUno6w1Z2uUluXxEn23Q13OwkbIWC50Fi
0pPZiGPhKEd2CeTC0JDltTi8mNndZvBEEdDUqBzwom/jQOjcFsUZtiS6FXjtLQIf4r0kTLsqDXil
oSh7KtqU5rifMwb9sTiJ/ti8p5b47PcG1BZ+4n+1hg+oJGDTJs2q7+He6hx7HDkvBlB3k59ADtwD
RRHchVI6VUq6ZCdc7XAOv+BTOoE/ffiWeHWHPwoJvyX5x4bmdoCG8s4L1tr9ghB9YvyZ6XwE1pRl
V/M7tiPlTAKqEkh01VD/dzIT6uBR9SDY7ADzQpCHpDPJyIP8E2m2pGkNLcWkywm9pq1g5nSw5Tqd
pErWHJIfosvj9ofj7KPVzU0ZMs6i2hD3E7ZHvEMYA+9+q/udLm2/iz/gMf5NUjapCe+9Ti4jbK/g
PVJg3NPvSC+BwoFjhJxAAOImUpMzia3HTyUCi2rLQeLQR+msS3Hh5SBep9Vb7FNHQMuEydYYr1aJ
ytOElNEaTXfIwJyo3QyRywPtE6C+hjW4plITAhsxAD8ds/jCwbAi1pOuTFBvR6yQf03JuhHatoXe
/sbxMWKiteXcC7ux6IqeQ7Dx2ZHuOu+Yjbf+vi8AIItGkSLPAyFeEvkS0gBRtaWpKMMU5mBBZCj7
qGJoEmIJfc+429MJKm7aTlP/B4MP2f0LJV0cQUeNXcZfniHItz0nH/aDKK2mNxvB4K3a+3j6xGKr
+fGyaRm0p2dF0fnm11j0lVdCFGQNsTwjHbw9yTb4WSQXv/kqt47bNi1kXx9bL2ftQg19H0iIAzwq
6Z4XT48DMKMjG07znfqYUBfwTeHgyg+zw7Hwf4emyG1F1gvGRxuUkMB3ZgJODqMSvSg3CKisF3xR
QYhBDmQeCaxZrEao6ZEH96doTwGNMZIx7d5jtO07Ylu1fXXH8ru4wHKV9cYmreYVx+fIwQ9emYlF
5dz6470yGGwyCyCObsHmlGJjd7MPbn9Ti86iDBdT7tZE/oq7Hy5N6ZsK4MYYBUlmxEs/Y2jGxXxr
DMnNefa01+wX4w8vfpW5oWQ57KDy4uZtNzWtZY4NzKKX6fiNrnFMqVvqcu1/jNOVL9kK0H+A2CCC
2x0t/eOu2QNqnqMyaO5QWzmE5D9X1CufMnJniUBPGHxijkTbhrNNNbfhoT4lnrA5IEl0iMtruRcX
GOj+13inxlPrPmk9sbjzLeM4f8QB1XbNnyeb7gBatjSYp0EHzA58cEhhuFB7Z2woz1945Zr2+COd
1IRhVIb2YzV4LJwyPaEj5cigsIUcqzR9zGnHeyUZ0O8WUwJn6QS6+A3+YYd6D/dqxOQKqzKlVCGL
hlOffETSs9w4X/OSgvte9iNhcmV5vVOXww3v4FbFEweG8nKjdxaPnRHKoKpY2DsCGjc5M5MkKK6X
Qo0LFOe4By3A3YIiNxKRSXnXutmBK1DNNJfWfm7axrwI2v8Nb8dnI2e5uXMkLgeizDCWnYhPf03+
Pr+10L33s5i0LfbmQnPY4YlnT8w0iVP3EYrDqRQsB6EsuoIa1hAfTXKUtwSi/cVxlp5BpufBeJdW
r3gK/2Xuk6Ni2V7o+TpKZFs8Ih4ZOQ7aO/EraPLKJnfS1DhT5LXkCkF6jmSRh5tEen08oKgf/UIB
m7WPEt9vSo+FPU/K/SHPVgdOUT8a3nhySZ34QdyL/8ANt3wP83MyRNUVjophWN9Y2+k+TRueVWZ6
54/c62iHNxPuxuBs3rdPsIoQ7tKmMcaXpCks3YY6dnF1W4kcUTE+GKTuWyg62dbsqbNj+wRpr4l4
kNm5jwKTHYYVzUzsxGXNQqhBVWg6pwIY0ixO9pIQZTCzUYJNNiN17cnTLQVCIZtDjojga46q+mXt
IlQKHFpfpZkRbKp8+JaGuN41FnRy/EfTlW8Tk7Pm4FVh31cgT5RYycO+QhT8Awd9JnVm0YPfbGBZ
HwbQl3S73wlxcvWDlqNfMlMiuRNwgKKZz3dh3KQGlqC7NWXKolkixsGfzzvT1Pd+Tcf2l1uBNHbv
XRwBNeKvQdfmdqNnxUid2K4ve95YcFbnPnbiy7DAG8sngKd0ZOMMfBSsT+bcKMUXv9SuK65Eysiz
ilrU07D5wBatr2E8Ory/EqY0NX4K9EmneN63Q8T1GnC9s5y63l33MVLhh90hw1DlPF49rvjXoVUF
ioAvgALtboHQ0IKsDsylyVaV6MaQNH9TbZhT7IJSlugH3B1TykyGhU4PjBaS2im4VnerxG0WWPzI
06B8KSlZ6nnyHlh/sHoF0QhKYKx3aLLaX5hYZDVoEE8g59/hEcD2/f/QU2K2+Y2E1hSHOkAI2kOB
TGxsA/IVM5cCsdNTRU09/ihR98BzHcf9h9vuN4R/RshNKr3wKixgPFiHeqBFJu37KgZeSNGIYm43
XODU7xuZ8M4ZfBI+pb9pVqR9HRGSwGC9hKDQGv1G7iP1w33qrnxcAOAv21m11y1Ftc56pL6OegBj
vWO3xewF3+Z7mmKrab06xhh1GRMIKefjitgMfcniO5t4WhhTjuLx7nyrzLrTyZZRE+iwHHAhFCf+
1ykABgYqX043MlJeYKbre5VofqRhiHSrGeGqZ2pZ22Dl7MnXn780lIKbpQ0EMh/kvNk76sNnFWHt
1ciGOUz+lTnLL9AkSCwKDGtlNyjAQSHJPVCYopf8082VbheoV0520HpqmoWtYKrf0/2l8ZE32cKp
sXhGB0ZgUhM2JLvD2HIy8yVGvbQS+4YrT/QuoqinSdB6Dz1FiuoTRRAA3+g8F3IRktI8Fi+4c7TB
TdlUDZPnqBBndhzkaodgtq8/16J9csY57I1lQjX8xml1h+vRKh5wusnSI+qpoWzvkcST3va2Zxrv
GZT/LDWSUF3qND8RiYujaAWtuwDPAHU2O3txMt27D9qDXVnxxXNsvG9Cb++Jqyz1S3Vw/5roKH57
O4ICKq+y0Vd6NIburEslPuHh3D/8tjMvobCgwxwhDtgdWSS37hoenbu1LWpzlPIJqeWchggUzGXq
z9jAi9T/s0w/3HU1M7w+HGcVVGvGhrzJ8yZnORjT5uujWviltBnlGkILjkaKB4nkmPtPRxhVYX7k
IrKq4y8BcS5CEcMl8S5gW84xO/EIu7j+EOXPXiDd6bX1f2k0+LsHO6EhQBMNxwa7X1iOwrJe2+1f
eXw4RLF0zdnZ2iMfLZAsr6m2qGbh3mxoyTwO3qgB+bEz10+nNGh7HhShJpcp4Ef6JgxyIKrJuFtl
bt/q/UmQaA39oyVIhp7Fs/1IgOqGvkzEKjZSxfaPWDYB6JqG+oEQxUWPKBEihC9B1e4TBQUa+Asf
zJTTijkn2Ul7aiEfIu2l6Erffop09/4ti7kxvpYr0obrhv8z9XCX9IuUCLbREUn6Rb8KfW27a+tY
8uS9yIueqMTAt/ESjiR7sIoISVe8fitF5dFjMWmHM1F+6LgPAQz9ukbH7SYHPcztoijeuIjdZ2xC
fd/F1DME1/k5EBW2BlFM0EglvjL2JmOPSzXN+RvDIODUyAhPiFW62CskdQxJZEoleljMrXLALUDZ
4xf3xnll8GhfOa+fkRz8H8Z98wBnCsdQbF+FftZ3+lry5hCBrqleu4vrNF3TKTA+hzwwe5v44BWK
HB5relhKUX4RJ/H+4ePhX+0h613ZXalmbXH6dKe1t+Wtch8hsT9tJoyCXbHfpAqeIAi11o4mLEpG
s7dXKTX/yxcRx+e6dzJJxgEwvxyEdBiTiSpMzkN2hE1U77h4RkGOKpc9DVKI/LgObhbcVP3VWaLm
WnrSWAVDZ/mF3IH6bh9LzE40P2dN5gogOsWkHe0qeX3q/q/JsDU9qZNTQVcEOfOSu2yfxWdnpRCa
7i4SlXbQ8jXejiW5LrG/cD9FIOisJIY6qJ1C7wgdYEazWKdOFDIFriM57Bg2v9yEQQVL2AzJLPHq
qOEEYqFy7LqK7eOfkUKuYWRN+nuAwbvruUgx16cfWPmujKSuRh/W+aBaNdV0tU6JNRNNoanjOLDX
pWdpYA39OUBdEQQsJSqb5QfyXS34Td9pSvJ6TQUi/dJ3ZwFM4OpNOpXlgogl3T9nywSJJwcOIN+s
wT15JB4awfbrL3+gdM7mzJ9aWbwCVEulNv1BPe0+1EKToQjZcyF9mNUeoMEY9AajTMfzSNENO08N
FnJTxRODnOp5SnbTUU5X84uz9SJU6rf4Ga3IcdQ/QKsk/V96ZqrpyMpmCJMX5Kdn9eSz0v3UG/2C
FZ3+esWwGjxlByLZcY5TTvmNOAs4f5rcmcft0bYqKnp56X4LKYV7w3iTx0vcbBomEOs/kSaSmywl
vMn9AqyR9Cqjvf06Pv1+uwY9xAkD/JxQ2yz8bMOulIuXGCHog0xAFEUbTE0pv6zutcJJcFxm1GeA
aKqWWWJzeOvJh8K86MFgVD3Abp0pA8PzwrEuAPyH/QgayKlJBpqJ9U0qR8GmR+u5vLtkzT1/EH/l
L9jKLIAAe3MsHOuKA2vyfUv7JoArHaHXO2/alpyJh+2v1epUstAfokzb6WKQf7l1NMSY2wLUhprS
TUjIgUexcbXQGp+uitPgTG9xMcLqeJHordOG96J6Z+Egt+RrDyOq7dCCT6xaE4H2TyNSf+aTPk8K
KLdUWEXe+CBfmqX0RfOMLToMbgwQNvl60Z1NdNvHDNi0oZ28dCQUZaYg6sDrPgp7aP+bMHNPzBYF
tnUBpsyFXF4EyDv2xmPe9NSqbslmK4QvVlKNIrIc/qhoyT7KwNCC+XRyMeQ9ElVDSM9tkT53Ukpy
omWJrnHYzkVFIpLPyZJTKVDDOLzdGQEUKsrExR1rls7RQlZIJWQR13vMyIax9huukAfKAGfgnZXj
QnlAFR7Ya0MzOr0ij6AOOKaGlRTcLsAfkY42XEeEZlvRmAwsufLugq2eS93vixVhh/srCakCBya7
V2UwGzXStPGOYbUs5TPKsGHW67/SbRWqzG5ilu3JoWLRqpYcxd8Ps94JhJgE8vHxA7PcAVcvdBKl
+hyB2reH6A8hWU2PpDjPwT4nDmBWxQfV6O/7hCw5ZYa/4lw+4XEd5qHul5dcRVsxF0uenJSQJJIN
Dm9TQcSq6XtyAeiFvogoXj2W9xpZ57pTapPclcc+W5uiXr2WTXnOe7pupgmXpzFZ+Yqcr+ixdo71
HW2hcaH9duXplvavZOi/vwngbTpv6FPt074ZRsHyGCDlEpx4kLf/leLbJBXUYOQpvylAz5QGxSUH
GEpstxgTHOaORUPtDrtEgyBtYyJFWvSZ+4cbhzOTdKEgmk+KQd/VH8yrTNk2dEBZxurfqjaXl58U
T19MgvndBFXZmkVEJZEITAzvIxNtiZLQudxfkc0wfEsfFeHZ9Zj+s3/ia13ZYLvOJKrg/6GUSyla
161cpak7PGWsahe6YB622pD6Qrj8DtNISL+vPKCWG3Ygqglpo8OkV1HdncmP3VKeEo5btivLn9vR
Kg+676Z6l2rMn3EmVh2uJXI8z7GlH5ZbRkNog/CF0foixvVS7aR4OxumJp/aNVD7NsEFDK70Ex6k
zN5CIyHVCDzp+UxbQS/J5usiT3GdSVgSdYUF1s+6LQvSm1WT0lKDr9wTA3Dm5d01YF+PQscdGlPS
aZdP5xU4yYavhKJv+GIq9tW37KX8wd5JpvEszuCZCatcAg1POxi2pasMBJntVkDPIPnZKYXgn+ao
rWgpKtZ/tYttZJe78Tfa1JCWrEnj0UsTy3YWRcx5gch2KuzygnVmkcOt47yeIbqyCh3c5yT8sqYI
/ufLRhYn2fj7gmWHEgwcFVZAtSffBTWH/niU3pjmxLWFhgciriVXNKumSteN0p1qxLewBeroOy2Y
3etJ/3sZtIsl4FR4xiQA65LzaZ4KI8y60RTDEc1BaxfWl1d0PHwZvpKD1GZTmSsPTYmbDxOjn6ZF
53jX+UODKxt70rxIS10cd8vheMphdzVvDTPhb14nNSoxbOnJPxUYIwpvgncrNkmTjkKczAxChI9o
mglpcx4Ms5hWcsarN9cUw1m9pMqs1dmE0VTpGjMFrvg7TSE/nWJr3erBOMtARIBqDq5vSp+lP9tk
ugB6rWczlyPBJfzKiP9RZokvI7vdkw4vh7FgUq+2tLHoJk2Iq/KuWOrSpElQqpUdmUQwhK7rSehn
Wfmhs2GdoR9GdAaeffiKMRHrI8agMfMDiDP+X/7/l/vHpxvZSn8T8kKQOooZW6FbvrRS/MqzZFCY
wqWfuYOBv41xKpHiqV0A1Xw8ae3Xq9eV+snToSrPilfuh5+4oqsXT9gQ8V9DzjO2B+JfgdJUD/oc
h54no/r4iIkpWSAVvvWzpo0dVqp9fNOB4XJekOUirtMzZkOKw4ORw2cTPVUuskSChjvL2yXY+1sM
uvAm7KanZ2rPYIqkIGHNsoqQQYGSCV7dyKVfm+jwB5w0/yggSPaKKpVT7c3FGW8JUeZPenEBvbKV
E4nwZ7mjMd/M4Yd3oja25MvJfKRJDZbmNrLITs6sWhQy9rWm9PD8lrj3GzXPd5SBRK+9s7jwo7k/
D/oPP6aUVoiIPbd/2Kf91S0T+wSLBbuSVhUWszxsKpxpdnSx794zCp61WzjiJwbh1BnjhdYAv/gl
1aUu0yVqlS/wVjWutkRtIUuvS8/iGVNDjxxoc0IDNXb7b3qPvsvJ/05LgWhPTyya4csno8PLUTLw
P4LCj/IdEE+suiUr1cYaiQgpYLmT0QOGoTk6jdybt3jnAtFDupZazS79MgEs/E922jyB6rq1Twi7
pZItfKR9m+Baybr7I5GFXTXurgftZywP39M/sTzBoam0oP/QF6lLIz4x1LvJ/sYdpKUNFq/8Qvy/
hDrMRlEULbyPB4d0WdHYo6UqZuM+98HKbJdPShJWMperh0i5pVxwH08u9eLr7Sh4Zv5mGbpTsZz0
stptfPr0eE10Mt891VFu9no4fhg8DfUOv+PcY3GXzbYl6k/c6KVh3rYNKbMobZHGIpzado4Umcwu
aJg488zKbXoqNP7WlXb6Q97BPW+tQTYPxuYyZZ6iNKWvOal5vO4eanoe/VScHULrF5Y0qDp0BY9t
zHGd0cByd5SnhyB5uEGpK+v6tEZzoAk+eaK7D2qWNagaptyqVoLZ7LB0i0oKeXFXMvx2p919SK5s
RLqgb5BBIq5W/Se9rkq3ZG8Oc7XkjvjoF4lBf8VuyTeMLVlsHGj+qzJb4vBImjZ3g3923gMzU+6R
gztDAhD23L51mSUY7q+R0b0JwkMzvZncn/icNKPIPEVufK0wk0qP5MbPDFbdsEwiwsuu6l1acT0L
H5157bAI65m+eNoXSQfMkLc+si2jT6bI6NyXCv17BctEVkYvl1VpwSMkhYzNz0eG3M13iTL2HKiG
RtI35hGZHe5xLM4JheND5tL0qfzeQZLz1y8hRgVvJPBMceD0v6EmlsrjXSTLTWVyEVLzqIS4c/q3
QEW5VIGUgsaoVBe8ceKjSKzY9w0TRE9mjlX45ecrAFkXgu7xI/lfTBT4d2U9Hup/57NP+0PYYrnX
FxceWRN76yPRdoM6gslGxEo9U+5FDWRdICdeWxd1S84VGhPK0al0ohWOwk4PW2uXmZlVrb5Teouy
o4K1Sen1EKkG/n303nv3KaDGqbd60BgJq7uIw3kYrpXEcI8KSbMePodCDXv3VMm5prIpT9TXD4BD
aV15VrdQ5p7580SMybUtgR4w4MgEKT7JsT3DAz67SDtleoPNaAfyNz1SIyN/64L9R1J5RuVv6sSl
OT/uxk4gvtvuedbZml+5zT1XnTBcj9oV6Og3Dri4MP6L1w0WztFOf/JgDGf53rp5xAf0pqPyOqze
Ev0JGIdtOa0Gg1Q7rcrutlC4bjGKBUpiXcxpVSwlfgAZlirD6ywJLORWX84bWfRrMUkkWuMx2CLr
nzVx49x2G3E1/BLZI6r7K6mRvOO9Zk3IrBmgZOvFiAMYEmwroEPOxDhdqMMtuD3SGufZIP7SS9mj
l43ufOSdjyfwT3AM1MBzibOXxs21stnEeMhMgJ4yhT9jcGb3hBmFTvk24B+FfK2NEPZ7x09y1CY6
912ZKf+22cASL+L87K+cxf2/hvLv+ThefLs92ZjCvJFRw8kmeGe3H6hZpdCLzlrqOB2n3BD+1UoD
RaFuS0uLK5Ij8X5FRbB3bMWd2kx7xNDUo5BuQj7ptoKvYMo++wr4uKQNcjyOZQ387MwRsc6pwkHK
SYyxvGdaM6+vAHzBhj4vSWgxFynHjCdzi8gF0l34aWo87FZ26EMgCagA4FsHPyVYCnXu7S9N4rBJ
Dds0oT3NnOVKWGCYnM4FVVmMh87qKrJy0Iep1UyJLdWsMYAS8nNky61u9xHUD8yAPKRGK/nsJeuh
UOBXTP17/Ixhp5l8EYUlV03xxN/UFMmNaOqpi23W5UTPKJp69xXYOcSCBQocr8I2R9Ps30M9q5L4
LeCCCYWisTLxrDh+nD2E1VlmqU6CAIWkB0zwHuPXgQ+Sl8OS1jICCFE/Ym9kzVWHgytCGnSh9Zir
OU+I8ntLCY/9E727BpoFgfGhpDkCke9mZhvncCY2kUztsElbKgeYVHmIzD0k3CQ1UUM/4rgkZNRf
bVhzgMKAsiG3zzmdxA5rbsD+UtSkQdIJ5Oqe6A5UZz5EELSnmHyMKs1R53wAWbcB+0kovJcZ8uv/
cDiVRyjxUwrmZ/i9e9R149q2vSEGaXhHnjF5EOB/8LEo7ebkYRxVdIfMSLGg9Py0Memycv/kqzuc
2WvsK8V/7Tj3dehy26ZF2zIoBOABqZOEx2FAOCZo/Dm8WmC4j+9sdGjl3ulAvJJkJ9+gN/Cgm9V7
N65YXqFgxXgPti6Y1S+6CDB6bgL2l2AmwTux+JGbsPrwpyBcpnme3M/ySgEnzhn1coIm8JsJZjCE
uBqn4qz6vRgbj+ZehZL58IQjfFb6uVX96FeCKCNYnrjKf0AMQxKChwJGvvroh4oDOZtYJvU0p/4H
aPUH5qo8czp2j/Xlq3iTIRyTMGiCHhqar7UiRYKVQOSQkqrQ4mPuMpZL1OyzS7R7vIbjA5LE6es/
0vadSc56jB+vugJNrtnjU/GukO/+cVyBdWeS0ME81YnQNu4ksEpzdcMk997CDrCSZ0gmQHt52CzQ
kOumF2BmxmCJWPqrAAfIMkONYq5+n741xMX+4PecTtRbwLUACeY1WSA14ZzGv5xxWnjUAXRY/1eA
nCQaPPtgbZidj4ETzeCX43tJN8a2JGLcfGnno6jNPFwO4n88U/pIM0HFWuKcFdV+4qtGW1lyMsQ0
RlCRkg6KySMJVzQI0nWdbSp42WYDj44rgUwq8aF+32SKIufu5Xfdduwvh/xtC/2y5Cg2ll0yqvLD
z8Q+oL0/9j6B8GfeAcU4M+wf/gJXML0VGbREY+amNDdQ6hkhYxhJSpa2C8rvWG65qGw9KwmyuZWC
1ZIk/RASBM1WFw8AbME0clz2vfUcjX+RH3QIMYxrgDc4qZtt/ptFm9Lc+ZjNsprE1vPJrBlXj78e
GkYxhUYk0mwKVThINla4Gg4MSSykPskecmSpTu4fAyFA5ChYrPSvfDqjnxiL9G6S0dj8mRR3Fd4b
FQ7hqbv0/NptwW0m0da0kgexme+oHbJko2iwIMZHxSqTCTEYY/auUVu0pa896727hOBKr78bfQHL
79DVlsaiZUkRbp4Sc65pllBlplX4l0sbE2P7GEfdJJNF+hfmxFvhuTkrSHF7AlhEHg1SuxZdQhN7
oisK1UqZDaGLJ1nEVHduNvcTX0spy25M0lI71JpnkmoXuO0+YImHESmLzOsdBA81DG8SUH9UrSpO
IiCa0WYhnZ0IL5QesGtT8O/OVMJpLgA0FUhWCKca+P53AcdmrH1pOaxrfL1+ovxfwvxuJTFQK9Ar
dEIT+Nb2L+uTPTEA2u6U7I5VSABFPyUm5iLS7Ye3616Nbzl56hGOnyt6SkypCLh3ByyN4k37c8BT
zJfvChlvl5EoWmglLybKMJNee+gXfE6rMNxlavmIXd5m3G74R7ADbY8razQiQjbK4eki15QALjTI
r+cBYxqsLeN3WomHEK5GkGVcd/6OBVPP8aJCp8UnW2w3NOAU5SNT3oyZU+zKyJlm/0X7LCOHIYaf
OPi1RT/4ZUV0OeybVOdSuAhoOUqkVyY9raXX0DcL00Z5IX3GyRtBJeFO++Zi7WtahE7xXGpR/9Qq
AFnNR0xbwiMD60vHOo8E6Lih7V6tNTcY9FgrJPLTvkmEY9Ubx/lEfTwwhDBkeCd82QVeESKmP1xx
4sWBmiUVK0SYtgoLU2vzBYpylFQoYnPxMOzDraj6dxGYtVKWRiiue86+t63jTVwey3e4/CGQM7jU
hUPXVcntTYZLSA9pLuoR1g6XJf3lwyxikxCqNLk3HSkTvvJcQqaxfqffBLaOlh3IVxEi79KF1qNn
mR0RJ0FzB42d6gsmvVDFODHM6Kvii6aaNpNQT1tLjfcEjvqDM+qi7kUPO+xL5C/45/rX0mpSH3aO
MBg2C77K6QnqSUJVst8Ha4iUO6haWv+GFp1vBriIe9Jt7f7tRtyhfVq8DMT87LwGOC9qwQHYdIfK
IwuXQVwG58fiauCdM/YjyHsVPWvLC671JjGBwF9EArsQamaqK5FUU+p8pO4ZQ9uiB+vsbeZ1y8B+
N/cXJ2T1b6PdQp6sqfa3BysMsX7fPFP5HLrauRCJHK/x4i/qcPBFiZd40qaSBqQVggKRjk3ISasX
VFugdDKTj3g79oa8q9fD7GH7SS8ZvLawywFcRf1Qjn0Cttr2le/jNnVOBNOi8Sp4E5smUv3ThDW1
ZxUz0loSY07cM4ncB1wQ7eeZZ6SXfnJJOHQ0XELIJd4NEBFeYMOif3K88202KNZJaRWWxnJSicox
dR1S+vDsUaZAHqwCm4zOk65uEFdKfVVrVeNaZ/L4lMuwnK0fTMN0qoi3AcRLKAhFu90Fwl0WPBMl
N0fsxnm8JMAIjnVlOXaiGzBcFbwo+2UOYikmHgT+Ody04kOXf5tGcPZ5HQVb0xtb83InQGq/YslF
9RTHNvaMAmfP4luGOiiHeGwk9cJnoWkpLPA6rM3ONWlMAW5LicvfBD/NZSl+79JuEMGlnsoGBRaW
UiT4tdWz/MnqmogGGtglH1I07mtSzL7sl3uCIF9oSBI3NWPxn1QCIju9FDWUZ/0wwB644287Elia
Rdl8smE8CDUIcT852M02Fun3YXy3h4SAHPNm0cuici10yF9jSwJd8r2VMcgXeHtXWrokNdFzz9Yk
nWD0vJcNZDWz+ZmB0ta6UazMjFDtwqCFuJ1IfYHcUz0TVd82dJwsYzRH9fo4adfnJ+Zs7C00kvV1
Nzm/yf7PKeVFuPazyTCHwmj+C6H63IPEoM5zjhGIuhlcYBy0Di2maKDQMyBaOHGgDjjLJXFJfqJ1
xpYZdE2JA9bJBMDtYoBBhTKEA4bTMh/42QmhvREZaJLe8iZ7ZSPmNRWfK/3kmR++B7ih+EOhPEkf
3Bi0kRB4MAWAPZp+fgaMub1HC+w+XKw7bx9TZKJkfjhvJ+GIGTbFBnVudFnI4f4YiLKBHIg8EO1u
to68UFBzc4/7cYSj4LT5N331Ia0d1qMTKo0pQhRy+qLMnWVGnrVFPGHMWXYhkpRFSKw9Ck5TcZj8
uMC/vlSTAHnhsccNZO8UbuwskaCH20a9rKb/b5aCO8ecHCt3ReGPTz9Cel/o1QzMnGIDsRegfPIf
7MVSTNAHWFE6LqTvD8sfzmDxLnbVk6mH8L3oQOtY4cVdlhixoKcpqg6knokoe6LS7zQYUg6YlgzI
jNwZS4mgdO7Q+Va18Ed7g8JlVU2qqYtYCC263hjPVhGUZsmGpdlIVT/3F7RTFzEbV0yDXE6+pRMb
vklMUuRO9YdOI4S2B2Q2+Y7aGnauMJdA4AEv0wKmpQu/xUA/1RJ6eAN5uarYLAVVWVNFyo7+jkq7
hFWxaNcaT0xpA5NpfUUQQVuiefRzhrmCRJRydMm83/gFYYT0B4xGdka4rLLVvcP/DNir3W7JbSRH
Uf7Q+qulWQcqiAgu36x8CRNBgFk+hvPoJ0lvCO0AMHpEmu4pIKNlX0AfYL3a8XSyxyJJmSmrGO47
nWsDOrzVjdvnNhX5YJ/xJ0jmfRW9/yRPDUrOTULAuRoPr2ILBsif8f1+/8KdNFh/2rActMLxEM1+
KU4WnVI4ncpEhp1GCTlrRR5E5ESiOqc3nDfIVkFeBde/SyRaIQLQtBjk/qZRvn1Xm94cSN7nVsNh
QrL+lFa2dAD/eFHnoMD1sxh3TUaoKPVQPcK2HN/ThvqAYM7ctxX03uvp3Hed6xf3To5z6NfjMaOZ
CBbL6mKkxABYaF3xSByN6Y63SHQr+fIdPWf2UX5eJbiojIqw3GVijU5Co5XMyGzUFLY1lUEJROS9
TQ8vkYq1W3+AyfXhJXJ+W8SHU0VYu3KBg2KS2Kd8TZte/mxcVn/KqPZxdPxy0U1KRmf4uJht10up
1H0R7c9De3CIMk6ofUVUG/gWcTIDV9Qf+aLChNECXddoO//tXLMoJVauyLIu4Fv0PbgnakoyFmdP
oKvI1UMfMBWWJS232XSI0LZnEsApMra4laP5YV0r0igDmrRfcUaL/UkEvhCIafjEEfPqef74G7mB
Y4unvZkgXrlSmHb7pqw9fCY2/Of7UKcfax40cvy8XakG7IpfxA6MW9TVWtbK6SD/HYmedkHnm+xe
a+tX5Zn0ODadUnkQcd7F8zfTER2id0lNT8Dmi65ZLieChmXs82jxpnFEdMYvdXt/fbIlkTtNMVwq
7eTkefDHV3UYXCQSQtAuQBBFqhXFHTr2FgC9SrBuefDHccj1IM4xKcw/j8msS/4BBEdL7t5hqxxk
PJCzcOZft82oZ/YzV4oZq7gsILXkkWaY/XFv0VDdsqBa4+U6Ka+U25+ZVgq1OFx0+MXKNVnfswR3
4rPNXEup/U3+1ap8Ju010vcy6vv6w3d1KyXDZq6iEGVG3CmDdSOIfxjaUz7P4yyMS2qHco7Ec+w/
UA5OzAfhIRouFn4LWOHGbZhhiq8NrO4uOvkn+p4YyIHjUvhdyYTPKu2bAl/CDcZau2YHc2jdGCMv
EjS+zq4FcpEamRYARXYupBo35QSA1G525p0VwrZfeN1gzlK+WrOATZpLqQe/F5VI88oOckbgh20t
Ow0Dpfu+xrVSNuD7dIW23xmWvd9EggFESvdgrG5ol77cY6N+f13PMG9nLM+PzMEdhorqI5lsqbnM
51yXQiwTn6/bURRQ0eONYQMVwQQuT3tnhpb1+lVYGea48eBthcINziWHfoHMJj1Xjha1RlibJntj
NaBnhdB5VMlfcuQBdMEckh+ddLbRpihmbJEEWW9tQnrLUrCK5b48mpLLhq3b0XL/B2Zl+JMWokqq
82/t+R7u6oilmu5hoIeRpiDdodhfIx2DAilnwsNsUuE8qyYzYzhrNwnxnP0apHUN0YlpkTU62/nj
OF/GxwyD21lA3+UdQ9udfxbTgIEyA6J5r7fvvpF9QIpbf0OfsJ78v5bma3yYQAZ45uWiA9P/ecgx
Vw/vLf3h5J+dIKcuWw4ZEsm7gf9X2c1v2LehYXpr6NJh+j67CGCWAwgEt0IR4YdQ5OgEO4BrR87n
ir7k4qGEErEV0iRF694Xa2zyVyJj12ahtyPPDCMys+WObA2oq7UfBysM15DQnaJvXgxaZQ1sbWLt
8akGuDFbT9lmloH+df5JjPA8UhqNa+eAp8haBFSR3l+tV7rnK6c6h7IGdIRywnWF82YVjjN6+Mcw
Wc5/DWLm3rUwXoq7jyHWR4RE0Xz0nMFKRRUzoCqD6WGFSmPiuBbHQNwVbHRJANsc11PDALEHvN0C
0Z+/nSJCW6VflSJyvul4A7AXJcUCXOeGo76uZkzgl5i0xOnD2T6BdgX0/M0lBVTSxbo2i2R42TCH
XZLcdB8vwWwYnMkbWUaC7SGpPx2x+qaJBm8ViM/crluOvyUa+O2rlqy26aUwQzAdpgv2rkgq2d97
znq4yMCxLmmhpPb1Xo+Qg9enlSkcZDRyLhtXWSjb+4y1nA4c0JH5VWi17vlq1pbBzTtE5WSm166C
BtJKtJsd5y8qp5v2WWQw3qiorjZ9FnlIA9VO+YVgIokg0DmTN9FPxI3Xle5de9EKytja0VCBog30
ksKz0cq+UHIY5ZF4NOuwiNqe4xhohi8Q1YVnKLdzjZhEtIgXK/muaBDbV1zNZ8cvy3z1iJpFf2i1
XCO8EofluIXY+36SRQIXlc8JK0PKHU0u9CsHEPPvPxND46SRF5Qhrcy0vgxM0/zabuJrUuEGAtQ6
rEe1fm2c33+YhnKZ6uk5Ipx/6DDCiIZkVYkNx6eewOw0LTw7GITXkyt+lWnVsETmxi0plJ7PxzqX
cpc3I1yLDlMhzBRfxt6CNUpgwMZJkq8edlCcaQsMFVGCOycwlOH2hKjdbgkXz5Jat56NvlwG+mmW
GtxUkpcGcJQCHjHBqtt084bLa78LX1dqmYm1T42v4IkAj2thxQZE8vmxRIqSNseRCg5alKhgPxjw
hWIbfD3NeILINEWrNu2RxNDdieQoPWc/cT+w1Y4oGokB3tI0hNKyLUPMSkyyWjU5mHv7vXj81uAS
oDS2L+4Kaa3RV3S/UdLJXh2sITPXmej2xc9+yptzs5w6lh2UTc86Kb6PXskh1HVazy9oKm54vz4z
0bT4fZrzUFGFc7hbplwv1eLboX/EJpBH0V5hBEbowsaNTIvlFsTM7jPpFCDQ8c3qzugH4NBNhS58
fn5NDLC0hak+Jo7DSRMeqxzPviHX4OiqkfE86TdplCmk4xH58qfrQS8J7ANimm9I3xMUb4nnaC33
V9JjKFU72V7fYREaH/qZXpXOb1NVn51cyboLJ2Mw6xpNhXRGQKBcFGknosjnowBE18nhUYOcY8dl
WjdPixzNI45g3dD85bQ40KGPhCqZhyq4PjLaXKbsspttwvvCN80B9W6lipdDpxRZSVNwo7L1n6c0
V9t18t8eK/YWtAyf/pEjVR/iVxR6OAN07ZZsvlZx9qiWsHwGxDckldCdLXOm6PDgCoHkybao4bV6
NOb9HF00UfgdW7u0FSor1/V50ossH1QRRvzE4ZUJRRhLFnRWLQSp+jpnFvQ6EzHqvBhCA9/AvBea
o5K8hItjAHRxDn9irIYvwMmHbO9WFLVy3zWY/Z/vRIz0uIirnCi921hQaF0sXrP1ZwQWPKjbTGpf
gtz6y2nGZy/iiREGvBX3r6rF73cpuPosn6iV+HLvBtzd5OJR2VaA3IOQlinoS0Xb/j8comTqygWc
FafZqph7XN1YUvXG9Vbyt/w4Whp7PL2wYnf551zrQD84ShfFdphxb/eW7zNkPEhENruspggMvMZo
REkoafNkkLCxbPebkLZp1OmqxCX2GyDyDM0kKYClwLc05INoAKRSa/43cYEHjNG4oD+8TX3SZKTh
dDB5xpkxv6xa6KoWHeUhyHeMr4mk3BnQfDQGw0sdKBoqXEEhgCOfWzdBX4Xs1FvfDbgE913ajVxS
QLeZcR8oIJU5PjJlyI35HSVx0sJRm36bPfQ/yf+wYmAgg71PH9Y4ByfL0XKje2UTm/Z2BCvDcl4n
Lop3E8qqN1NHysSAyU/+Wq/TQREcnzMszY4UDR3gtni3esqdNvkC5dMNpYF394glfeeKOEiX+CJu
OxXNtxJVGk29qSj5cRS5Gl9jusQ9v7Ih74F2DTYIAyXiCs5Dbq8algTAYPOBXyQuGeL7ez1vTVtm
8n4wGT+OlMo2QhvdR5lcxtuf6thnUWwUxUi1GFHb6ax7ZSxqGwuLNsXgxoEAXXn389NSAbsRZYjF
dzJoy8/RuQqojTBrlTUe5cbx6NHplvUb6qLp/Orm/Guzb5WxMGNgVAYJ/1dbllxlTKRzJg1ObkKr
/lVDe5A0DWBWkxJCWGsnYsQlMAOuTZmbK+UqUilmyGrHRhpA9I51lRRPXtB2xHKN7aMtdREaZ72G
Mg1HNEQLgoKgNsSJiXz7kEXi4MHMpfYrVsTCwKtPOPRjz3MDfIgQvuSxJjMb0ictcRvsK6DJEvyG
FruC3Ile/5655kihV9jePMVruXW+JHsCRWQVTvF2nRgqdfUW1tddYixQvokSsq4bIWX4M4laiX5N
6zac+D6l5DOdc76+HbpHnMZzueVXnOIwlzrNBEImn78u9fGJUFowzavTTEoL26MD4lq9JO3JgtJf
HqerrpjYkKqVMn2WhYMti3qzKCDA5K1OzRH7LOIk/0oTX6tLBV8pFCXH7M9nz0PDhixtVwua5ugd
Pz93/nCZhU34RXOZQF631O6K3HijtWQ4Tp1s+S6X9vk8KEjGG9J/I2vg5Rvg3YlIgmaR4Ofg65kl
ohfmcnyeoh9k+gChtwcNB+MGzH4C3NAn8UA7nGFeNYbU6rZqCIdD0vPdvFLaa2DX9rtW+ZB7C551
EIzYiX8m5j2bAr2mI2UftltSIUJh2bDg2RiibzIfudha7vhBLGOLjqgSFZo4QwuGGvUivWCYlQ++
cp0UOEF11Myv/9BTQHFbdcREUSFH/tgZ6iUvDWxkcCZupb13dE5cA4UfLqpHel3L6LpodHd7I72l
qwwik3TWkTlWoqXxUKkGEW0kPlrTl9YhfOqx9Ku17Mf+8I09+HaMzLoCFljd4MP6ctUz1Bd3TPQs
kOrPB8O6A97d7a8bdhf6ZX2Zz0e401Nm6ClBLvURIdaBwcj9eLsJ4sSNE39IegO9q0WbjydIuNTc
axkFhwBps4aLiDVySrj7o9l/vzqguUxL2EENEZED9ZfMx8K0tkRb0H1C56EfKQbrNaAupIskuuyW
Gm2H9boDXVd6FuXmKRPm4XsdZZlTSQs9WhKiewJgZ+vYHWbYULfgGaV+AOzpz5VqggPsWXnA7st1
MaUpzatBF1qJemRGSpDMBOUXRGJHZB4ZBB5TVRjRz2Y8Id4RJeyR91vZxbxp1S0oAVm4tG7EiBTA
hAcx7OYr2jDY7IZ2QQEwzzKUbMLC2/hx0WAtnftHxV4CpYNVwbbY/K81zrWr2yCRbeLXIMp3bld4
2QM9FNDyERbVhdlwdStl+ofAMpUw2hkzqAhFSdtjr6w/JTdr1NQwAmiO+xHE612P+YABmiZdxTz5
nL8J/Ls6tzskxmjIg6qi9wMwH3auQ0re3zhYePKEjuwB5gSN5OyRG8sgnU8BwBe+LWFwcIsUt6l3
pc2MS6HQDK0fGjygbpt71PEA30Rps0sKmMYYbbQtSzg0MfrDCOfwE60m9SyjmE1D8sA1i/36UEhR
7anUvjxgAMsQXY/K/XyZKm6t5GuoNLrFDf8Uv309V1RHxCufSYIgxKSa4a/ayXNiTgyezu5vv77M
HHEu1te6JowNmbgW9jrAxTbP2E8JB14IkWUQ60DTge9zF+Bj8swEqdSC7bLaW2p7O4Hmd1Nakcug
cHqKVqXyuVA/eD7UdRkRUayGnWYOs3835F7QSpW8jvtUI31USBLW24mNxY5mEhWFUKdyMa5NLPNe
syHwTmyJ89h5OTA17BVU5EABnZ362wDYPRw1jce43vayyV7TlcsFK/7LW5dbdu4yDsmC03ZfzE8O
MEERb+oMp7sdRMYUw4owdBP0qqMH5lmInYyq/EgriKwM1+a3mz165JHxoz1oQyZG1Yuvii1s4iaZ
lN81z5AqRvGS01gFdmMiEylYrl5akE9DD8scuJ3WS4RtoIUgwi8Ir0iMd4W0vEgkGWm9FwtXsr8X
PSH/7YUhs5ZnHHYSl4N9GHrvPQat7BDVqqMmbCaZFINNrnjRFluvQQLKAxwiSjsXfAfH4ICd43uB
dezRvV0FRy+OmgRDZdrsPJj4VFARWQAN4LIgZElnUSPkQeVl/iU9TiN8Q31LVEfsCCrumCWNKUrD
oH11vFe3ZguVJeaPj/+QjUoqyr8Hh3L0unmpcoXoSUS+Yyo8n2YIZY6YKqp9y1SHsUnvJhP2cPKH
MZllQ3zm9m0QoTobW/Ay0igZ7BC4gdl24eXBgNAQ6ehiDRvt0HhiLQmcI3DogdhYUWayHbawQr5l
bJOw8cDxnknT9pUjxX5CE2Xtfcnr5eKlayoPvDXUY5/I6ddVLDY9vZrUW4ujE0FvKLQjjmZwZXAU
vWUloVN3Mh0Otrv6WOwlqxaf5ILlQp1JQe6Vi/7XEkihNa/ZytQOIHAu9oY85HLlEU4cubYrbxXZ
tb4SX/OfIyBO5U+TKQrdBzGOevSGtbjapAu7hDxV8livFSNXJ415fJ/VhzPLfMn/U+IYddAbXiso
GqpN3+RE0cipBCCVNxKibKoFd2Pqc2an4eogRbYBn0c6D5LCtAlOr7YA1fS2seg2qZA81auS405j
x2snU3xUfr6c2wiR4QuWuZiK1MfQn+X2kH/DBeSDzlQUkIxqG/2p7rIQjHCmcsx3BUCdoEqDW//H
VJ1iJsIF+4I4hYGZhDNt6aaR41sA5mcoyBWvm+hhDjstPwodM3kTMINoar8frUl2nDmsew6PnDbb
X65QSt9bl+3m8hYRhzDww6wYxrgORjjq79kNNyjE6B5UgPH96cobicBNhdK8F7DvmnHEeoTi7t9C
AeOJe8z8p2M5mTLT133EFA1Aq49bM0PpJJYHSNvgM+TBn7FWA/yjp7HCSNeEQtmGTZ1HABtmrV8n
0V+5Mfhd8monKxem03ezMnEmd0sAWbgsIR/DgSglGlBGxm2opOXUmf+7qb1V1bfIj5uEEAaMg8YK
XHmZDNQCHC20neGs+lGG+vdCk8LkV4+nIgPyfCvJJXiHM+otVbZTo2MggJ98nP+bifvxO21waqSK
YhfPTFFuNSlaWQ7ggTIQGIOgWX5HocpFSbJYUC6WvPDIBUKKUCHgmZ/FFvWyRoixOwJg3WWMwCso
NguP3mnjVaUhJbzuqnbsNk8roOdZvjeEhhy92eleXDylQHDUgL49wObhHaWYePyDKXXLDYYjZZih
tPFzi89EYEnGGlkgyxKy9Itn5Dj+xQzU/llK5WJ+LQP1N9Y1B+D1HKmdsjDjCE5FonXohE8iWKxv
ZFTdKTR10dSuoecLgZBy52A+9T249tl2UaqK9vlaOaypVe+lp4aK2Q4lGQg/1ZXFCMl2KXieR91i
+kqA6BYuD/HDRTIb0Mmy9AveL9XcD8PzRRw2/EG8w3YznKfyNM9Jc8d/vbeuaJz3APWgBELWE17X
mfoKLfejVmyweZe1K3nsWFb5HZlwi7ZsxlxEw3LznFB6ONRvdUfmjS+vHf4/VVp6BHQiRzgLzJgU
TpXrRFxyTRUAwDKcp9UqTTDuhwufpVwUo8p0k08uplQCXWhkiXC09iyDJnw74xW5S4/A0c0QiLn0
yyHrnI8SIMt1rEcxsy60VsB7BRPs8BjbLjNmjfgFVEw3aSSJD1hF7DFSsBC6gjpUniUVB080XkU9
yFShkDeBrZq0CtBx6tpjRiOipbJjSv8KRET4NdThI8V8XJE3InQ+zvYsmONCRfNbV39UfErG/QTu
E41DSiOljQMIHdoINpTJ8E1NQGyQL1xLg06aKbKC8w73TbrlDGSa04RYVMUSTKsBFrNcf4qey3kB
tUb3pmrC1vgETtBG4dQc3aJhL3qPlkllOYvmGwdxRyVVuHO4Sd0gTCriPjAiJB4/hjuYy77PmyXf
ErdtiicGbJ7EdHt2sA60eFdQdscVeSxb8jvUz2eoaQ94tuVxUMabKtiu3v+XkOL8/MS8MSA1OD1x
aRQAhYKHmvOkPqPsQu4UEXG9LSCOHl3VnE6LJZToNZCgJUPnHTliZs5okhQmueBF3L6NylJ6uBNX
9JLBootArX9smXRbdsBVqDcvVDe7k8XKrHfTZHrO08dbkkzNI0XUi+dWorKrD13GNn+aHZIkMz/U
uBOgIa2q6BQ5m4nGPMgDAlTFBFB7+37DNDES2TFG/awgPxYC3QuDwBfPQbB0sfOAVmS6GOynlXBM
zdNI76iNFfktsE/Bnb9OjF/SbE3ffXJe+RNKrhvgq1qQ65SWdy/SwFpre5dQQh2fX9BmZGkowQRw
o9JQ63jAIT6pbg71uykcLh8ywlTBur85zeykOPa3NILcqR2fuJA46sFWzC/2dNQo+uC4kJs6lPlG
PI7UguJridySjbckIoC4WGjcLot9BzTXS8CN2ZFhpT1wYKMN9OGT3P8bhCB1o3UOeG46XtGzbdyZ
FbRn0EsPtA1rFKhCRzI69DXb0cehI7anA+v/q79/E4iApcxzW4jcggMwgLbjhIhp0l/S4n0o3uDs
l0sz18OARdFIUnXfD4SnpY0/TAesWfP+wiHUcxsxrAfPXsDWZcJMs8T7RRetOqz2cVyry9oZB2RY
RG5dg9pqkx0bf/fYTYWVn6wJyH9A4SqHQgIgsoNuteh4IoxGhwP3x27D+QSaAXuG1WjzQc6e9aLR
paizfsFnrdSQbSrDiB6I8sLMej/1hVqFG44yWcO+b7qO/jZcMpiEXIjZ0Nj21p/oAyav9EDNb0bH
sTdAmg6T55hYm6MrCEYiwn8iW553SXhHYyfDPr3fho2PN8OtvOun2yRv6683m98cN0Wj2Q1XGmZz
pF1pkB1In4Zxwk+PTMwpVNxYdHUTu6KXU8Du3hcAGsFlL40Rm12GqmRlj/5abfBIES6JsED3EYw5
OlxCOF2plL2bexaAtImQsw9BSrJp/4iOnuHS+ZeNPpiBQ5FnQPsM/o61I7Mb3XtgOBUdTKQY3fKA
FA+QLx3eMQoF/BDVX3CVaecEqEnoMCjIKgZMrLy/k3idMubhm8VeBEy+CzK6f5soDzA+mtieU3dt
/p2NjaZSZyg+p7RaiVb/VgzsJeJOXduSii27Ix7GJYEfXuihrOtrf/jErz7QvkzSy7q5rnmhtZu1
YQkA+SFNtWHkOK4qTmrMxQ/+5fyKLqZWUqq20zty4pTTN4Gqh1DlMd5v/PmfxbtnRqbEmQ32GohE
U6TjNbcxZ2EQ10M1WJKFy8xTAjjBP5J/E2b3pGRNIwFZYXvwWXocZral3B9z/1sEnsy2+PE3nvFO
O6BySa0rzsQF+23EMyyV9C+2DxnM/wCOF3EmldifvXM20Va/RmgVHmbuHErUpzZzUTDv7YLhCFta
qGMx02DkKGRmwpEvgwnvyG0LTTZgIA0kDh1MPRLN1jRyk3GZ97Ijp3HFZ/FfumSomqCqQ638U2Cj
oRH2z9e2v/ADVNjIwdosQddlA101gMNLO/Uhla8k/ECNcplXCUadjxfUr1RKsbIq/neC+Te9b5gY
ae+CjPaSqlJHF/m8W2J/sV8VqoxK9ZH0s1ULOwMjwIarlJibL0tE1JoxW61dxQzdZMdRwRlc/LVW
0U25bV4WWhBvrjyv2wSR5VXgf+WQQMxORCkS/OR9f4YSshqtO9gCSj0zy5LIOXWI5hria3Agm382
YRuGKaPkFHoD8CtWM2NSF+zuxE95eBIp0YYGiHwl2UNMgKfS4+tj8MdtbmGFWg17RYIjrUB+oEqr
eLh4o/HBuGJJTnC32gBX9wZU/Tji6pd/4QNBqv32L1jChzFaSCjxdd7helIPo+Yc9gxfQWmJbzTA
uGHkBgDqjlSLT6a1sw27no4jzdwg43Gg/5yA1M91UXl0awsYNAl/vRgiKXeTUTLED4+Khc42VO/T
Mmyft53K7nA8GgCwRBTasKvCLj8UmtYw8wvPUL32Pw3msYTaTrgjRYnHJMtzTVUEnbK+W1ikZ3Hl
JDYFbqu2V9sIbvIv3WKX520IPi0Lxi7eGmV7YkikzQJFiP9O1/DXq94nTPEzPgktwz4mSAZPOskt
ER147S8GLSiC4LFG2EWUGGL6F7S02+bWPF4j6sUcdUZGKf/TAJHQ2kKbP7x/+X03qSgANdYM7asO
g3jgly10Ir8oGnFKvgWGuROEPPenFONYA/n90bDGh/KIhCtvJHPKtPatQ0MhTvRPogNTY3IO1avu
4p2K/CJCrPO9RpRJyPumgjVYrCuP+hHR08jrWiz2uIhNkPVtUd3yzubPl1YjnIw7W0PQuFr093II
UZ6iRjottM3rQf1ws72C66c6smY+PBl5EovU5uhDp7UUpa97QrcvTEXuX3wlzBlqAay5qufkzSvX
G73SezCxBOCoMzfV2GgJC5aA46E/Ceqssq2IJCmy6vrL0wH8PtMF3++sn8Q+lRqVih/6AfbU3frR
ENNvDJtaJDpja8Bsg02IBiM0VPLOjY3hQUCp1GQWauQGoDxmHaIv362vYIQX70PspJktWdDf5Zce
Sm1pibPzTxqrZfMXsEvuBbBPAM329qB0RFtpzcxCXq7tgmkWHmmuQ2nYthzalwmvfwqLX9l5UHM+
nXeX7Pe2qgO4W1e9Ij530JU/2uHZB9J30gu8qH8UUMHGAyjBZtBbbgtkSvyWY+M6ZEszXhIVgKFW
NKT1cj683k4dJnbzo0fH57NbVblbtmjaFh2H2LTnT9ppK/ozESLsLZ/FCXz9f26oUtWRC7+blijH
gBnN2wnP+1Q87n53HWGuUCprmYBKCnDkrVlUdNCar0q/GwDH7ZgB4vXWBmJKJYAZk1Ab+IkpJhhB
P+LCCciGi3Lv51t6/WVYyHZyybOhRMEGNjARhHnPJIZcK/cRdDtrUHFtmai/BhCRZHUkp5+nmzxE
YOcw2ai/F1jmcyF9kir1T9kX6O+4tPKt6elQlRCeC13agW8nHISqeJDuSH0PS2+MN6cZ09JY0t9L
U9Kr+r4HYrABQnUQWxDgir5rEij/A2wFQ+Nb8QrsipQQHA01AplQOxKR88tZH4kVt9Qqc5SEdF35
UhUgxa+sVEuvG8XXU9RBDlmX5uDeF7DHHe1rFqApWDd5+uNyD6yKsKGxm6X1uDVJQcAmMX3R8AGa
HEzalMh/uYMf+u6DPWb8oBPo+krvuujG4WuIHs5ncr3ELRchFzWPDHd2bhzy+bt7Y+P5zH9LyOFV
fhCpjcay5UrM60QL0cEpzzQayD4kkBfkLmL3KKK7v1ThwHTIZya7C3xYi3Y9hRMvMOxPwVYfFn4x
srcacIQcqa9r9Z0RCSX1uZ7IXu+99uoYWqfTjao+qaEub6K26vweuGUhYw0vNBwja5jrU7AKTLrd
L93WMvWYMCfFs+5PjnSc1GvQKXkEPtX3+1oGYusgcjM/SEtBw3+9IZwAS+hx1vGLovdjePHDoeE1
0gR1LKiAQPMPJ9Buxsz+uzOkIDiAwFTrvZGLCxL3Xi6c2b7vrTk8ZaLShRTkZzEDxzJDmolYHG2m
00uHVjq55po45W1eKwC4c6rRhuqcBwsPLaEsCtl1i7zwFBfia2mPK0aHMQ9X7cyP+6wqGd8VEDRu
XJIoswThXXsWNxhRg7E6KOv1bJBRI3HNLBzfqUFXEY1P7M8KGnG6KzayQ8Pq5+PgyMllODB6shnD
ki/gQIyXmDKGnq3UHreWKmsfX4VytFChc5k5rUBWIHoptartSuVYWJft+TJONojLxji9shtQXh6K
OeHmyd9VkIB7o73L6KTJhdsJqGBVt97VXMT4Oo9IfyyyOg6uRVl/jDTDoY/8DMcguZDfMXcgW5fA
pYygLmTyt1clUw4i+P32+s5mTPBFUalbijUhjqnwbbA09d0Ch1T+SVoj5Lbbjsi9hBGp2Fni8byd
Gz9WiRMNh1kiXNCCmvcuEq58AoAZumwaFPonSI4tnyR5IFbchx287RT731LEehzrY9I8ubZRD4Jg
c57HVWNm5UCWMYMsgD7GadkB2DPQ7KBFSelf2jI1GV0gg1Cl6Cj/3g7HDxDHXtQ1GGqNLzAEV+E4
wBIKjxkrIys5WXAqqNBTOLedK7Qo18YfebwcGxRk6AizRCb8Xb+brV/FrRfNgKsujvPTJZKi+zwL
kl30jj+wab6780gKVG1mVCVQB+DdAQarhx14ZOjMPQsIhQMr+sQK/WS1Kn7YDEoJ99VQDlTrhIyN
hPvzNxzZW3FQQctlLBuGur8j+N/AgD1o72XjqUFA/8bWCvZXgMaF9nufm1TE3MSpMpD1Va/k/RNt
iRV2nJTmPCsjvMjfMV7PEzq73NXJxNH7PuvqkHq0CCIEPL7oagQG4/nR6FFw1E8/x7LrCxrfrtfs
A3PQ5TKNMihk8di0XaGiIrSaJLyrX/fTZCsj8xM58J2sU0abhE2V+vdpvO0tKtrIwjZv3m5qh5nG
rx8JSqxCZQ2aQw+blEVOT+9QzAuhcnLxAIyqJhaU96KFP8u5TDQhMsPyXmRfgkKcojh3pN/TIqer
HVOPGupVW87px0G7GTLuRDuXpdncc6DRr3BMGnmwqwt8augv2ZG84b2TGsBJeXJb4utHGTr4WYIE
2WzD9ZSwjXVHRSu5UCRMVDcYeYGr4x5IQjy32GHKHcgkUYnyW1KE8tuZyCXWtqj5FF80obS8xhuy
JXoDFh4LD2i65iscq2pDW6r5OD9W0N6ixC8QBQuv4Z4NpnuxHOk6hB+BvBzoviHmbD8wrdq8kdjo
zm9xvJ40SR7z+bCDmyHxfBSYujm81Rrhu68SLS7fceI52lIyW4uZ0DPClg7wmmJ8pXyQyBQz6aPO
jU1A4TEe2/3kGyWzZ3LRHxyDqnUrMMCTq+AHwzTJF6qbZnVMySreQyiyETqhN624HP98Hh1+Wc0b
gTC64BXfXMzmxAGbYBX/8ABjoivquqLXMi9nTvzsAFMFbAd9XsoqhaRqt1IRKxvFOZF6IV2PyLsG
XYXhWmMUNmf7DZLyhYU6ntWC9tdqgTYoUcubqmhnU4zW4vO3QAIMZvN5mF0hyMB691a3/imzqYEh
yHFPbKtZZolqsMESJMTWiBRWSN80N7+bJ8dywn3oEkJiL+jH57HosWStJAj3hG1NRIGrSExwWUke
1rOQMKxBQNnpgeztBDtZRN2b+B3D2FtUmchcFk1IYWBjZxYHG0FcvjHoHYkM3F85inxpPyAgAsu3
LnLtQfJpnznlBUMn7GcDcxdh24/nosSZbWmkaPgwUxPJQjZL1uYCg4it8H8TNnf6QaozfPyUBehc
XG3YbkpzeDfD3m6MhSG3uHnqQtvzUzHwtYrhJroHzTtuKJ5MDkunXnWIcYlk4dHQ0Gp2ILA42czD
eKoPUTYL5VsF9rqlzrG4I4j4z9yz8+b6Sb/hfMW5oRqmvQ7wBe1tKKLp2kXD2eFOyicExBDLxDz7
4/TqUAY6/u+rKZWaEI3EzhHxKnL7vepwZwxBLxEy3xb04EdG+nPHx8MGqmZrRdLzuFfZ4Gmhb+Ip
Pkjp3rFI2TdfhKPokyJAyVPFJGi/U9DVP7bmo74WY76j0CzkKnkhiqg37OzWQlKV0bLNmJ4OHQLg
cY+Kj7LxxrJ3uMxwocb1A4CsOy3o8EnMBBV4Ygy+9DacPoWbpJKjohG+jrRNeMY5H041ocEwtdUp
zF4WLsEmLbLf0KoHOn3z/m8lzp3lVDCv5s80ywFrUsiHU2BnohWgHnI7VI+ZZ4aiOZcoSUDwb3jc
XtbEGzz8U7uioH5T4seaEu3fPTw1GzvrW59TXLDtvVLofkO9d8P1s77T99U5chZIQYCykwFxegO+
mvCJC0RmAYiLellU0xcSHTkWCXXID2xtyIUm6YSNQGulbRZNteSp0fL1x6sLU2zv0hCaOWAA/fR5
dLN3ACdbSQuDCRHVOk2CJkB7TlNmqb+MNi7ZZ8YMXBmzobBhOAAlbo6Mbw2tBK5yuHEKtWU/JAmA
5XrJsQwgNbitvwt602XipffW/6BtxzE4+Fj0dZ3iqBR9Wd5oOcNZXrce3keuBSFYpBbXkVF6Gu6P
kTc2ALBzJcwffZpZ0mkZ5LFWwQfeg1R2c9/2wGkxC8GIhgTsGZdyEds8dWWEtzezalzM9+ZrX/YV
SENaXxa/t4PNbjR17ORCunQOJBAcaBMeeuHpLCmRAMpBTx3hgx0D84LLSE1CaqWj9KvC8yXyZHPU
eSMzA4Yt24ICeSKyxM7SRCxbul6DpXzEp1GA/4CoKyygGM+d4ifSM7LX1BqexOSc3+2ikjRK9VLm
2eHxGplyn66ypafKDziP2TNYI2XE3gfePLGdJVmX8d00s1PhqyWgyt2PhAtptvLqe1V087iIw9VD
9nz+eXaJ/eNAkdM3TA4cs3gBrOm8f9CDUkEwBCReMrq6SOVGf2A/fPjy4FEF84dp5r9nK3hHNx7A
vtIlDRrd5GeE2hs+VuEpwwEtBRFtsUPszdqrfxx5P4EXx851RkLb8SbBigJWQWeB/eDUsYp373W1
UpVuTLzEKJnGib+fL/RECgQUi1b3ho3ld7P5H/GGuaT2C5vB7l6Xnzj6Ibfg3yBrlmoRz+S5MHoo
xnCZSHCWqmrM0ytrC8tU9qldeqQMwroRBpUYZ/1p6uvOmnW5FG6SvZ/MMF7n0LE9FKaCUfoGdk0H
UIz2YgstIdWajoZ3+DVt1RC66dUfXobBX295mX0yZbmojt/aeCY4bkwnWqY6IgLmdJuQfBZGt8iL
hCti2OtUVjBJM+2Q5MuyWVvLlYoAef/2CaxIyxpUp7AeNXDExsfj3IDpRJtKXnFZ+9LB1iyRwZ7k
ElwIb1+dP2vF1CU+iOwAOpB/iwwlwcfh5VFo//CyacOmUbYmIMZRcwsMeKlSL9/5zDeuCVFHQeL+
Wr7cCQqOqL20dmQETpJIQSRzolADdJUo357kSxdhBDahXt+O1gRViXLTOmeOiCcu3ExUlkQCjaEl
rwwql8oeGVdOdoavE3eZzcHN3d47qClXIXikB5P3+0FN/kOf/xfmJEinvV4auLf0L7tjZymU+UO/
ZL7LQuurtm+/DIap+5O8xjiwBDmaVz4M7Es5kFPj2qoGwkuhx4e15J3kfa+nO/QXENidQcDVwXV/
Qo8Kh6uiolD4RRRSAuLyg4cTgzA3Z1lA4tq2hbUdP1u5mcF11Q24omkwfw+u1ENdEsC6KI+Hw2TF
b3UgzZGPe2a7Po8VzEyaab1FdGKf2Ep0F3YL0T21Xc0+3G3667I5CqQxd5dNBZ+S2PDfFASmW3T+
MbOG6OEvg+VBwcludOEC9VkHNHrw85mOTV2GguQnZ6ZvXzfY815tpCUixf9Cmu8Ljkjl0g7QkhZz
tuOm2+HoM/DvdesFGkSPQOvQwA5qUMBELu7U5eBpOZklbKYWWxfEhrEXlns6k0FWVXMV8mlLMa3X
AieSKVRMCjdPn13Dfi5iBLUxCa6AZDKC3mTE9LwRFrI/HQkkm5xxn9pETQdjmczGS92Li41kZPAf
uP2I9ivqxDf/Pp+r5ABZoPwjLlrHWmiv8BxXUnULAYWtZT8WGC+JktP1YAMeFzJt0wqgRhyaxhUs
RiwVaCribPPtcXu+Kpc1WZQlv7CDKXJsLWIiuhynXS2TLsKY4RoHSDJbdHwuOTkbkccKne9Cf6yA
6Fha1MqPlzxtg0AG9y7EzSDd3gMtIsCJJARXcWMTA6OnJNYg56kRMJEYTFVk7J0C2waeN4bLn1fL
YjHdTo92Pak3bFIsaOovW1VVpLiouSlKpuD1GBv5aitTP3xoOpqif/rladkCeVit+CUWj6jfrlqR
GPvJINZnOH4JQOiR/KMP+HEpQFFHSmPGRnv2ydY6E9oZBQZUQfPjP3wp1MQQKOZbddbBH9vbqvsw
UNvsFMcUnjkfLdfB3OPg9PHP1gXoB377fdXcoDxcxomDFva7sngYxZTwOQNUhYBXr6jb2Oj+Huro
3pqSopF0ly51UFLCcUhrIMyrWFOQXbWkTZ4rAdZ/dIqKdH1+kQL0X1mnuzfs09B+EVaMCz1VN0Zh
BGGpIjuoJqzsK1ntQCBToGc6uGTWXydEqx3AjXtFqIRAxFwOZjhxsak3CFK2WACifAwDQem75DYD
vLfhWTeAZuJ4aueT009VfMbohKukh2Usmx3yNF5odXLLAXvumrDf/CITGvoZcnhfue7vB+aVLZD5
et+6iLBrD84cc7fgtAXZQbtx7Dmr8ltUyeImC0nQJDD6vKPNrFlg+NkicIeVQqXu3L3QUJ2yxTYX
y65MQZeyx0hxeC8NNS0MgIQ9jKVbFybvyzzJY1yYPusX163HPR5o+l1Gd/eg6M9q6ohkmL08Tr+N
Jh+EjXH1NW2oTwC8v4q8s7P3rA4f81aygpL1DLY4f1gBO89MQUwcS7GmlQYhHZverHHdCvUo3UML
p/u00GZ6BCT5V56a9PjDhxzfjrGGmfmmzUyjeXdTYdSmoAvYwYqJJaCjrDBfYkM7JkvU1DNqv3bS
/EgiNE3hziSgngd+/HVbi8XBT7yUpVYSREnZ00BPhfAvmTHOVXWuOQDJNkjojfpIQ0Qp1AP3faPK
LhyH+l4Nmjrsj7rAUgJocGpyK5MzlSfuXzfWN9KWtgf+usVcg/LaW2Z/Ulz6lHIyXfro0qfqSWvW
RSQmX64yHp+6KyEXeeaWJ+WA68JBOaoAUNSU0rNo5m9T9fYdjLG3OKFTGZAQvYIuufIgMZNt+5EC
QCCE2sM0ySsPROjzYOL3dUzcHMhLFYlawtHp5PafaXCh8LRw38ZF45XcUzAnPhF8OAOUwcKktpbQ
zzD0DEZNQCoatz6linOl0TkUOSlcJrQ/td1UzorwURVKOOqySJlPFzc2ipCmdvCbY9SxctbqToiE
cI7fWZkg08/9fZG0616bPCGYdeSpXd32QDyXQ9K50cfMp3gBAc/zbMiz63f28O7GV3wfedg3v+dj
i01BqlZZpW5fVKhrY9mjDPSeCEHTgAn/W6hLDD3clIOnY31Xh4mVGGC5eY7MOWTp5njFjXBjt/wn
yknf2mqbIPN2qCRMrBUuFB61E1MUSKf9mMzYWJkoM1hMhZeu690GJPg4AbsC2p8ZIb+XxIYLuU12
sP7LypNNUzRtYkYg9Qoe4QVOApTapM/ZocJBSWYYWyKU3EDAQ9HGiPWErXiB7kwzWGG65JhcQ58n
W+sfXy9mbfnfe6O6CQUmYrvd+rLzAmY1MKsz/MQArp96dZ3z+fI51US9/rVJbSUislLIZikOb5fe
WWhnWOqLQtPukLLnrTrA3/GyPdDF+2xMW4QnzvG//m6IcUmEX0sz6+/xm9Koy1slWf0vAkSG/CqT
gTO3rQ6xpRkr64nQICp9C6RH+mN1MJvEu9XA7nzYshVWfilaQiVjNCNc0bwGX7nIaA8aL0V2bIIR
RbmFOeTVYbtWo0MOn941IbqcIHat6vdDItUqXbpHVsz/3kqp7l37UkhjMU5EQwi2XqG/9GGExs4n
ZIerF/gZflk0Jk+pBuiZc6OLhW2MOGLCDLKVFgUHrrL4JFd+uPud07aMQnbyx1UcSBJFlypdAFye
jQe8qyub+CrQubkJloJkQoW9XA6XJPwMtcf3x4WSRSzWytD5XXYDMlFoLmj5hTS3OIfWAj3n2z0T
ar2dKDugaxZ4Gi3fkkaXnsz7msNcSZjNXDfhCGQHe2WeGh8L4Y+7suyi+lCfSgcHxSDwnrMVN7wI
UfkqNVQCbtxMT1cEQvWrhqT0CbOz5psjca4EzRw6m/mLIn9OmBKCHs7YUwQ4OBXtR8Ozifetnkd8
hWiqe3JMgrdtCtryC3XKjivN/jFwA9HOhuiYcnMifP7njj4z10DrpB5apBOIBFagVf7zR7o5PrQ+
6USL0aXQ6rf01uyhnsLoIsPvlauGQ7okvsxcT+gnnrA9qHNbWRqFAN/xlBj4j31WCCLst6LW0Uz+
QRZKXvjL1lWLOzn+mDFulV3lPpDNLSrzp1vAy5prl4srzXIeLmoXrLG6CsjViW/IN67VeuCYHs9p
MontXhKveT74ryosbUiRycvw11KLpaWIGEpG6Xzpe9ttU9uYEzRnj1UQ6c/xyYv7wdtZziF7CDPj
uEIfGolr1lsxssbAHUtLUWbGsjHF61ZT+IR7zk7S19DIR3OkeoMKLWnuj4If9Uo8eUJkWHwQfXW8
5ZiPQTWyfOvGz7QDoou6hWrW1UYetzSg5aauN4GgLaZUUUvlO2zJt2imipRi8nwSO5cHnRzaHKHr
eWImE3rkAvaNI10vEdehgDXWvtKfe+A//hgbpZXYgMubhdXnX1ZQjFgwjfwJIMXPhGSW7h6eLs2x
4utTRifhIzyquR7phCDllqlPEBoILNEBp/FhwG8hdHXTM0q2FosaX0qhV7FH5ZCRJag+tHm/oEf1
AcpGTCXERI98aJxVvqYz25NCTu7AlEGByVTcP7PODudU0KKnlFKZP6ouUXV7OQ2ntMW0aG4DIcnk
RBjbi8JNcBlMbeKg6Z01np1umus+TSIOM326RKcP+XG36va6vSooaWERdSW8sYY1EFzIR3x4m7Xq
aYq2W70ihFwGIlo7/uWGtmtw/jt3/1b9xr4rTshv3/7ZbbdbZKhBWaUpH83tw8d0TkR159WEIHVq
hBc8GYcODPLyxywzcIS8COKiAHIxt0JN1rn1q1V7UlSMGvACq1lOuToXeH8SHFqUtpFm63XFpjhz
V4dvO6LStNno7y5Vy7EYESXfilYk+6XIk6j3Qz+4KzDsr06M/vREyF7Mpp8YYssA9DWkHP06Y32/
AB9KqOGyzT5W+1uIQj9nEzOA+6DsADaqcFaoDaOAwyaA6NZeQ+D4Rc5GepkRCPyIKeh6aA9I7SFl
nyyGS3XvHdv4YbyBcKpLsG9J6bdjxNRfNyYPwSpBhAEgYlcvH8xP9vjZPemg0iFlk4CPSN3jUMk/
JQ6OAMpg+6W0AZJMpHRl/KZwafFWyevK4oNQUtMbzfm8OfLKUeXGnMmeVLe5bs60AvoJ2mVU1bx9
ovqKjjhsjH9Av1dkO+GHhzJdGDlXE+YiVp8+rLoipRS/+gy4JVuH4cccbuMDa70cuDE0WTwrErob
ge+O310IKcyYHk6EO5Ump6EVid4DsCT46PzB7/C+DjEcJhiseVZ9r6SHoS6Al3WGNQQ2sYoZF6jW
0S6GkyLuIqYgK/k0KIBF0YzboRsstAXTHKSrA6bncgwB8+EYABoKoqQ7aIqOjcms3XxE7T2xiZAq
venJno08thaQxvwNnBQnyQrnOQYCANxmUhIhVKMTLOtJ9Cy+sYexGKVdLtCEzTYC+lbiLwakbLs/
0yxPjP2cnKh7gVJBF9kEjUa5P0BaYORRaBn4k8u+FXg5R3uZm1AceDps5nRt5osdqu87hqV8qT9u
i/1dQlaNa1mEhZz2rjQcu6ijbaxzWA3uIUjcaSTvh1H5nNgY61Drlac4sQGoVSnHLODnZx83NRyP
kq2oOa5Xyy0Q+ugdlarT+lqxqk0+r4OrrGprqF0jSKrdQZbVOdv1M8H8zZhB6IE8gEZA6WvrWD/M
qoYTcFg7ELRSA7gUkC+n0bnnQU27crC/0oqFwOyuTYpVcuU00YpXIvfOskCxO1JMI+x9Ezk1PRy5
nJIOTNBQ7eNcIrap6HiQKtKzJekVukPzsvEYzVVAGtZKkm55eRbQg2tlKHH/ZbVqHXDXS1kEord3
LXXfC52Ri38xQg2MhlcIXr1XkqtqtbMzWfEnzo5BUU4MgYABazYBV8E5aR6Mo3aVwvUKFg+zDoPk
Xp1+Fd64JAHNl6X1gRNS5cREn1YwQipb0FVv7BdTYMrKPpnuoQwZrzBLlf1f2NearzM3rb1zVSFK
w7E7gTVff5BFXKbRwETIVp/J/zJTCh07oZgBf5yOSWLpDmv3ySYhF2V52NppUYWv73XYT/gmLQKG
h2fcU8PhF+OLHWBp4bpd+neyazZB2r7GZ7pEUS3MwGDa34j1Z28RWcg1WHal7U4XVe0st1xkCKvP
Ynz+5eJVXy7Duy0oLTAh+3Kp4yysrn7spa6o5h3RfzJt9mIHqXS8vpk7GBa0iWfDe/VJTCurMbiW
VptxOOFNjjHAXk2bwn6S/UcO/89JRPYwKJj3HrfDg3IYeagHCFU18YsdlSkiaKhk+QE1D8FR7RMy
5LWYHk/ZfcCIBLunlNoiuo8IsRQJXcw/QUxVz2EsynRHOm4BQS9bjhXi+Mh8oQrgAzc/6bZTeQVK
i1QkhSIdj7YIAY6OeYLoXf4eTuMttBkaRo7X+/kS1kgLV+qMkuq8UfnPIHffkqEWUNnhRHM4q3uG
+IjE5K5udrqBDUbI8S8o0cC60vku1LXsF1yGtdlhZ849i+gjWXD6Qm6enubw1EGkxGSj1dLSwTFh
9jAkPZP3crVqdBQxtjAwz7iU3eG9o3SwQOTBSAJk9zXnhlNIKTqaBFJFJHmEjBOxL2W9W4zZXcex
wb+CGtcOENscOZqar65ioKaC56Ph2HUgNiPYPaNDwpngBXWNkqSticHKJo0/HyRUMYqu559YnzYr
Wiuoy9eEH+jkF1da0+WftaXVLrBdfihKM1bAnBcnLrcQyDty0MqcnJJHv3t+HvyXOGq4OfyOO0Ol
q9ST4ksKUfDUSDi5aAjZXne8FS9peAyealCd6bnF0z4/i3Pi2gbD/d7/UAzFQozJFxoKNBusqKri
9haPIxFxdK5Zbi1WD0POssrmxa9k9wn1wvwYTxCurjkC/4j2hfM6n61s98HfAz0gso874NBC4vzC
GnCKr8l9Vn11zvF7RCe9vITtRkrFmywFM2jQULQyDpjTloApDii0na54+36jQ4F2jEDZS0hFUKvF
+wMjWFHbUm8c6mUjxg8Di7ZpgV+x32NRFNcyObNaLzAu0MmicioB4V+WgPgIUNgAaN3nU4sAOkUH
3zwx3HEAaAZwBBc6bhhx9VnLIpaGjQb7FP9ePq9+neEp3lvwES9PJw9DOFCS9I0T+aP2sMBaNQPQ
hFf4NpcuP7I+pwar0Veg/RtylyMTDgrIdGhe0n0A171uCucIvALbvyL4/q3qYIL3/GlByfBebizq
frCEw3tq6+t1VBWTl2J/djja/scM9vvZXjdhi1slrsqofdhhMom11jQIzxyyLJq6EmZjyy1gDQFD
YISsWkazfnY8pNUH9s5+CWUoUWlgDFcixAeh/3iZTozuvUffMyHsZ+jrqzl8ArPexDM+ut3JMJDu
MZn8ogomkV5u/4t8160nXucH6pBWxZbbEgvzcYSEZrgWvNvyu4KNLTx8X+FHjZRRNJ27doVCHoZu
HkKEsp6QZ7XFs1St7oPXeVcrQzF2kOzX0u2HZr4ysg6ecq12ZHzsw6BIWj9KBtoE23VaFs0h38lH
+djuPOlyZHGNrYEOM+NP7JWLfvaqtfGZo3hW/yOe8RUvSwN3JEBfvfnYSVH4oBP07ceyOU0SpU2S
ESCecvfh6N15fR5WQTLER1JGaEVDP3WsfDlrQ33kQGn6K6A2xfYvkNvF9+OiN6xi7qmT2hSFvNgQ
YEBvpH7/I3WzCkTvxJcp/LPr4esxpMtGoDtEVrF/QAmpj5MaFNM5YpN7Ud7ehKyPLCBhzRkW8ENB
fZzvpOaXlk4cE9FFn1gMWfIf1oNg3Z0LXRO4ZVuIDR7A/ii3ukFCjRH+vV1xE4VsOflclMgWcj02
4d/WkvZNd7le7GnZbKUtqAv9JF8g5qw895J7fuPVAn6awMAGToDSUUMw+kJpZhIWSAoQqlHSPx8f
wFem8ksUT3HhzkzP4eszyIDIHzZI27p7VIAmT4hvDN6z2XnCzhJbifbw/w2/e+OEYSoi2mhWMi/9
lCMzHUAHVXlFncHz0kvAIFYvOA/Iiw8dFL0ajC1sOhscigznJknF+4uegxjBs+gXcXogIE6SankK
PyBDshSWt9P2EQuZPdTNT4DEu0jqNcQFleyZEidtEuqziepRW/pBgOr4bxho4QLetSriG1j5delG
ASA/EiBsHC8zBF1lVupF5cr0dh0GmWsmT/iaZf4gXbKEV+6Phc3tbs0WrJKksu1BQEI5TuEg6me5
63zEX6de83Zz3vnFMzvsclcZ74zVINUXFFWuRz9kLpxtwtTecffwTpvYEx6uWZtwLHxI3f3WnFBC
0hUKortOZ8dwpNUReE0thKqgs9aVj/AdKfwXLIaWDfqLKmozAawlJGTeqaz53827E7J0NuD6qmu+
x1OmYglnSP+R2ulHaMVyA1BHrLDRNsaCmZ7/M/ktivsBPJNrH+qnPNiPQYG6EG4z1HlC9HWM9CV2
VA0VMb5Ont/cpIDixZ66p99OUdl5PuW/zVpArEqRlXEMRIj53Mxel7R+Eooz5DcwObC/FgMRAlVq
5+LlQ6AnoESOIXKYwzNh3ztL5YN+6pFP85ni7JLjgfQffeg2NCRobtyFnnZ8h8vpHS/o37bxqeoF
ljqE6WuUb4q0OHk3QHP3wMr5j0PP9bQXuA7ms1o4kTqe3dueuj0P96F3YNBgvjgKvfYlpHNdCg/7
bYE6KTXtclq2KXb0FbPM8FdXELa75GjGFwZtG+Fq2LUjG53hmdGT0Om2w/nvqGuO+MvXErbbW64J
zuVCtWCV0Mk4PqQwiQD5PAT0H2w+5CJwF4e7ZVQWykHfMCXG/XCRk0LnplSI+c7G3uYfwjun45OO
DjSvpxxuBZWs2xBUYYJAt0wBk/cwc9TfzyRLij9RaPT6X1eUk+2+3Ply/WkwTCLvaOPwX0tKdC7g
GYLbxPjU879HPirc3LFddUiEXkG/DPH2uFkpwYuNcr18MRjIBmWjj2tINRiQW+MSi2XWzQ8Q4YOQ
VLjvl2ZWoXwc67XHvApne211VBfOs5un4FqOJkEWmt77K3w4SaaKhfQmHMTRu7ogiSmnHE7666SC
/yrUQv2EBwFH4obJ/kL3lgPFGEMMGo9Ang9dwfZYMwBli+xNvT97ryUQ+UpWKDHSkRMrEViKffDr
FXPaEjqiyfYDNPJTbvNrhhAPynDeGUAslZWEAjjCMKqreVm5zdPJWuCIbdgJnPl4MDkruFJ8xv53
6ejJaHdOi4m1+mPNDD4HSpWap7S2bRMo1zxCF8MwCF3hkq959v2BVkWpfpoDRj2YCST+2XbSI7zl
9FpKsaMm0xDKtij5m2n1V9DTVFwAfkHz6yjT7/w75CJVaEu+K5QQtzmnhq6JsUI6IaQBZz9aCyCT
vFjgR/lLWlOpiN6/hQiWqlLWeOeOhkV7mYXB6rB3i7w0jon2+mMcpEAUJTO9MQ0a40+CNC4O252J
oRjgSBMBuNVKVHCOk/p8GrXwCaWE9iOjToajtxuqGeW18EDNEyNwJXaaH3uAVdaq9Uw9JCf8Ba4a
J5XDxqDTBDl1w6QDRrH3LqAikTjiO8zMJIRHgDUjQzRYOV6bRe+iNMEsFjTyin92rJBFxEBiY4i6
UvboUCOIDB0kNhAt6pFSEeUWvfVc9LodSRk6q1sVmt5EaccOTbfHQToO5F7BFO6s/lB6PFlUtmX5
qtqEkgtN/vpXo6W81WChSAoBbbPhJ/QPx5zfmMAAW1LgAAueWuYNK3SdvhQHa2pF60TL3jdl919T
8swiV0gkSW/FApcOxu/Xbwq7wLcEZp87Olvy3HCD3M4LFHKDqGVgw6vBlshXKD7rqYSBoQpX6OzU
hIC1zHiwtx6uSEWqinsMCBBBklWSlNhHja1kORDe/BR5O7cmF8/4fk6SDWj8v5aFYQK2t1e5shK+
tQBRlaqwWe7m0DA/FE2TeKVCOajYF1bYncCACRQsJ0kj0BoIsISENK88wAQLY71uhp98lBCZvQE3
mp4P48H9sJH5sS5c0mIRRkL/48GJynET3bYvbzksKw/pOOhZfFH4slYfnFPGwraI4TO3ndWpK8r6
U5kTB+ispwXntZ2x0kgfuDlVRfFzIsnnRRLKnydDUmJfeLD5gJtD/Go8U5wjAdUWgMSa+txtezYg
RQB8QkCSD6FvLNU5YZ29kvtKqghdnC+L8IJq7dJlikxkgFkvalgc9uqTd0ndeWrk+ajNgCko5Lbd
wJJmi0l2kCB+14I3dXgxiYaonP69xsk6868A5lEmZ+acoRsVdAINlGJa3ZPsdLFKwA6JjqV6xa0x
4XBvB1axbp/MOoNLsYHVwipyPnzN9fY906nO4BmipnZvJ56mArYizPP3Gh+tg2hNojUmmtsdFmlG
+dFLzBZY7EVqGMszPPpD6r2FDek9aBdNVOJZilbBNzS4EeFw+o52gZ8YNivIdrILk0xauNqKr7xt
1yOpkNcA3I61selc/+7z7G4wZRZ7VkWs0h/wCbjJMGvJzb0HhGRREbSbTzA30bk8K0iH1dJiHEUV
xwKwQ3M1EBHZ7643cCiyVa0k9YULj0PUCL/7GWBV032ZLzSJd9U8dNt9WM8Jmhs2Gqwfa7ZVfLLD
vmkse/xNc/TR7Ja7z877mvFXsq0IC41xdL/hRHo++lZyDf6vkIZ/otNsOxSa/OtfiCOZrR+Ka8aY
Iv23/7OrZi+LlSS0t/ZmPZDivLi6xZfH8FykkvQddJQE9xK0isMeJnDGZXoT0I6xuSg1Pie4DN8m
LUVww7YH+7Bbj1FWzRx6JBTJkWo0KJvYO6uZwiARSGGBrZUva9Ryrw11/q8yXlfDOzNuYoUsLTaP
ih1Sg6jZn+CNWMY1xEyHZ2Bqw+tl0saMn10dx8e2R/OMi5xMfE7Iz1lPfSRWZfQY9mTu3u1AUS3Z
j7CPrpwFdg1H8xXD1luuAXzIHRQTw3PW8w66iTlpixZTg5tUIMSpaY31uIjKcWnI+uIEa1F15r7h
mIdDPM00HXqJUly5c5qnYUwUsyrKIfqbZL08NBk7flZ8b7OHleC9wwjvKqbtLQ9YDahgF1x98HfX
GtYLhuu1bjZPhDuFzVbCdavmYWsVlRasPO9X2QL3C68jh/7RBAcCiAiBO0goP48I2ZUIMG59LZAb
s8LLzvBkaMDJhqDXgsgiA416P8US1MuLdWg2kDmyV9hM2gt9bWGpRH31maOxxpLdLaK9FgiC/YIr
njsFRyy7H+qmYM2yE2M/GyoUOJ3Hta6C32cchwSr+ZtGPJu8eero1RI8QDkFmdOhrcN/ZvP+kcfL
GsO4wF0+3AAIEBDDfETMNAFKONq7be72b+SiG9DSeMGB+fhtAVo+pYtKlQ0Yvd2hzBqLHXtFYHlj
CRqsVBkPjnpdN68nMMzd8gstSxJc8PzhxAADevoGr4i+Rpj+xY7ZV+UPgO6D6JbDEgvlvuUg50Ay
M/BNUTiDX/w0VgehCx0SzY6t5fw1XUG9CswQq9KXrDS5n95YgdIGGBRKpru+eqqJsYiKkKaeQ46N
Vc/ws7aDg+jworeQHOHt9D01aWI89x43mTlS7rrSHBCt26KVhB+Q4ABtXEp1jWXmxLh65ysLS+m+
GSwKdy8x6fuZmJdq87XAmSELXPPho3ZVAyaeYSRWLcAIzo1vmNylE/cqWDUgfREKxlt5i5iCk9I8
uGRCzpS/xppDSofklHATk2mOHK0oWuMKL35BScZv4qLbiYXIfEJtwVgnW0oPDk01emnpwiI8qiw6
69yCY1FSrouM6eDFL8/Bo3e6whzfoVq63hkDcQNKEKRMh1fGg/iPzZc1RM/vJvCX0eAkA8XQomOA
REgpa85jCt7JpRqnw0Uyh8M8Ga4sRGfNE8WMu1QFcVD0S83bVdSJIrAJwWbyDlDU3DaqyVEKJDjH
toLHTEjQFxcqzfcJfKbWrPxzC+vdGkbOKxgnJpz/Lu1+VVTzlA69/Zp2rdarqGmZkpdDjII15LLz
iCCbc2ZgEa3r/ycDkloCucJu4bQFnbs1nGmaykdodYu9fhPB4vku04gBqoLphN3HMMSiOIfH/3Jj
P0+44u8bpdjw8r58Ye/yfMqqMrnWLcMNpFfDeU30lPnbgTlcr8BLBscAJxVXjvOifB3dlMzPnfTR
UqylOkzkQoGsnIasSHVcz71TzvS3NlQocWQ8TF7z5nBZj38DigkZExfy6Bjt+VsdR3IQr0dXSe2u
GabnrD8yqSyyQ/T1XppJIMvxGYi4JuyXKE4P327sKT8RnNQsZDF7wH1unVOiMdVFcTi24QRiaxPe
iWsVdK8xaW/+FHuhFPItVRFcV6RGaIaHo4mrTPUh4msXHnNw4yQate6Y2rwg2jr+dSi38jgxTG12
CadlbBohQ/xJ7qNiwBS58hkRZB2iuPc/OkMnYhpPkTgo1VlT+xf0IshOvllNhNDt17xdey7A/Kcb
LBYD1OqoqPHuWDMRiI4jrCOSQ0fgXl9YnB+kS0MiBLiHX+72LMMK30lm2RlRRJGdaaXHqIbyhqcc
Gpsq+6BAxUpoF3z7E0KJsMVhX+lzoF2UoIDlyebt1axRAOYMZ5ICDLJMm8KQOB9AA+FYZCKg+7CC
mWcUshHq8l1lrtuQjDnGOlq95g3lULHZ1c4zgRAefAetNsPfJkqneKeRYwpK+NqxWqwmC51zewTg
gmA0h0Nj0xPerLYtj8P5YJINpKHMbcbPPL7XbPeEa5W6YocRBTFmRRtMM87XQlmYZ9VOPOWYbPIy
ZpXKOs5qEMOrUrzhQZpo7wdqflbAWi+O1kgnux9od/En3nmZO+f8akBZjPxW7Yebrd07UmDqyGxE
nN2/70QAeftpVUss7ZG8m+rg6MO8KjQPxiUrMjZ2yEjSMl8glb+KT6CWiVrGb7YDZ+j3FbROTidC
s36AxmFHJWz7v0EapKa5kfv5qCBdnO/pjCojUSDhTibSRL/HAWv2J3jpnSK4KO3877O9z6Fe8tMB
qtF4MAoquJT+DkgTHWPyDxY+ZXrOhX8vQ4ZFBaMC/uwEnZlpJ2EeKfkN2vcaxEYX+fBFpSi2dheC
Au+EkhyBRa70t2ExZC0jcJt20opnGKE/snHB7imROjQ1ghGRIPLQ7oSfWZg7Ue9kK69f8C2UNBpK
uj+eowhGEbjibvm3GRA8FS9oI2AvA+bry1BAu7uldtx3q23uEjiOGtDmDQT9BbrO+kptkEyPt/eR
k3XDgqXi9f8XJ+11PdrlnMp6+KQn8Nlv4dAs+MF3gbrLCIo/P6iS0PNE9mh15GCvRojbPJlfCZzy
GkVE7Dj4cildHwyhwL9znmNdXETKeEbocHNC6mMZ9gBESNeHpNJjmRGmIBEAtX9fk/3fDpeDBk9C
q03jIgiuMAzThhZV0UplKwduc9NxGzpFINOziQw/dgw6V6KiLA0kT3v85ncSAKGvvGAq4ujQVMq3
cHCydYPf9O5BbFj8eG4oQHQmhaTsIdhEo+XGXL35nF9t0lqAfATkpEs5F4YzwXDpAXvZ/s0i/dy7
F2CvbDVrJGAK5YHR1/2Ll/JKGJVW52yj5kLGqUdCvidLWhMHmdww40qNYSNf2TUZRb7NgRVBVK1r
6rHaEZkODUnMqA28hb8vyv9OnUsXC8gcYxqM01S4SwMSXTJ1DwSztgObIwy6GSMmmuxkTboSuIsF
g67Qc3t1gHW5b3iub6Fs8sHdZAQfzh9kPOwcX1Gcl4IRrs6SSN+IuR9i3R5tbbAyiV75ORyTrTKV
UL26ctvt+sCg323vaeCjy7FFv6zrF6TwWYJYJFTr2mjR+FmgXwYmjAgkw0FD7whR1k3oiSeHvudK
ZY+qKTc7xgTvpUxQ4UL2IGEmyF+IpQxfDoNXYb6JDqckNdwCUwt9Y0vaud2Fr/J/D5beS5IF4Vet
td4zDgmtuqFQsfSNgcPG7uCiZO6WSVAOpTiSe/7dDuTANJUxCUoImkhYTjoZ+tZuDEp9JK6Aw4jX
9XNsq1rc7AMhIXHxSe6biFEIV1rFEFoIHsqVxl+lUbJTqwCz9HOZP4zdxqSlEkiWgLI7yAJfDHQ2
3+vpSvTdJYN/B7ReJkXi/N9Q59VRBbhmtwUPVqy0p4zLDAnveey3wV4jsMnXSvEWtZ1gmY4wKA+H
+r7EFfI5kgqQUvVzI3buhqlMTz/opzX3ivHyVth56MlXH4Eq59CQa3wGqBmgDSz0jPIbRfQUKs+7
A4bP28q8Q8USyOqk6YYWO4nnFtjNB4IUG4ZMLguHr72hLgK8FToHr75p68qS1dzFODmauQfTQEc1
TbMk4C70tED18uQ9FjsEwlKyADD7zAhDbbAEwkY55I9YSoxYFQG+vaiW/ykM6y9akKYClvfMBAey
IE9KxNZPfp86OUvso+jD7TVAptVzqjoxb7E4j9/ys4uLjlZKUFBoSq35GnGRMMcbkJDmlw7qIe4q
+uGxmZJFlt7na5lRuVMc5LgreQfTnDcEMReHJPddCwAU1VF5/8ISCM6iwzHEiAd6FEu9JMXddJ7z
Hu2RBizRbt+rjC9YDcUNGscMv3tiVv38sBOpN59QGrXUZHhrTVlj8UAuj+89rnoepBDKDzVWJ/Rc
KQAZQ1oJDieGBBikirDLrioHpNtIdCo5Rz+DB/Xh1bGsVn08qRTHEJVQK0bkGGfOP9uiWRnbrcsB
uHbP59tqcA4/XoZDHOB4jQqqnuZytAcr3jCqgpbZZJcqdqju+YfrU+7XlC3anYg5ShapXa6wIRNP
QrcQbSNjp2yo954N3K51cq3IjcuVYPY1l83XdKMzwU1QdRGTVD3UcNs2qFFjO5FvyjOWQ2dgIeij
YMWPRIUAGF+rVuIUUQ+7O6M/08ZUdJ9/wsQ1gTQWq/ZXGUPLmTNSXEkS7cgTNP+cUZmUu1j8k+4O
i8qwRACU/L8rF32mbIc6BlbDn4CxirLhnj9gIM3IoAV0kLY/C6r6Ii24jqCj/oj97PhXPX3BeNjF
sWcTNkWMArNsz1d6d3DFyvu2nAtCCXu3xNpnIUWBMtLWxAj15yx4o419fbnY9IeJWZDx5+RtG0y9
J4FNXVdcbNIfiWs1yOWPIEDRVnQoPL/WgYBGHA0VRC08rLVOJx3DeluNB3+GcbvZJYFXboTiDEWN
jeNHTDK8XxBfVusYhUZBpNYKOsXekTVCd9RAoKGdtSjz68jfvt9IlA/tHUdUjkKu132MOIEFClWA
mvH7dDpT1pQVvgTmjHlnCm8kv9J+P+5sE8cbn6tLzCxgENswBfyqZa2leneh42W8cT8q2FoEg0SI
Nnzu9VH91lk6V3jQfZIc5AlraRs8DPfwBuUHLALkCodMAmvR7ebO5uNP6cWTWm3csWuZtOranU5e
t6L1sKKrviWqrGqrYxXcDPz1hjg7e9pXCIr8MjwxP4c/UG1tK4tLWcm7haKYsN8IsXbnrvICMIoL
w5ud95RzsdnYIk22jVx19L4ROMRaPkBUkEkLYFHrb0lMFR5nmFzoRY5yRDcnCnDSOPiUrFR4gmdb
GzI++6gCGQYnSMFTR8rpN5SqRmwGZ5XKtOUX0FC/0YsJiYHlNX0HbM4HqDGRVSiwq0b1bJC055zx
J2RPZylMrnrqEWQinEOcT6dQvChAtCJKHNb/vUriLwFR+gWqiXbXehTq3a2Ce73Mo6v3yqEqntS1
+sR+Wt52K6LVqxH9VR3GEgPmbxx8mi5+XbeG8WMfQU6cXgLaEh85r0LlNZsoLyZyGiJezlZ+dIHA
Y/r4DKHX8tTr+FOy7aG3urWbs7i/r7AKm8UScN3pEo6JCslSfrkqvpxXfFoJrkfM3iqNsfZJSEV2
JgOQq4gEOb0XO9iJyel5nzftlE7yyrx5jd0ga8aTwG3V/FotdHPue8GAN6VSSk9PbInCx+fpv4fR
924+h/CFOHoGNS7mJLvK1BuBYTE8rZgedPUhQwKT+KgMJ9IzqqGoPiMBJdgjSUNiniJq49Cffki+
fmKWp5oixo0m7szg+nGzkF004hM9WTYdG8e7+CqaHxf8K8qRVWZxaKixQ+OKB6MhrRSZ2KK0YcWI
RB+OM24ti84vRrVduJt5H0UAd9gNauK18F2CGru7vnRUa2EiD33vKylYkbdq134q6q7CBBXLN/Wn
J+sEfPj5ZglSGEJx4fI3xOfxWD0A/BBYfzPVMYtejRtdyJPXoaWQO25S9fxc1FK0C5Fs1/g6mDtI
xjfDm4DVfBZTgL73iyfJElULZeVOYvTlxDYrDtG8CL/gVgRtCqsGrtZH763DyWyHXO4wvPqJ87j4
22bbPzzwtiqIoO2/7GCXbunolqU0NVG8sfCGuyiJExJIWzUxYJ+yo0wWBWdF561UHSwrnxXnjVgK
rE2yCCSg5GsxbVVCvVcRYCRkqB2nb2RjqCAgFCTBz78lOZ6v+KdZ0+NN7e6O6Y/fqnmTGerdWEED
Q8CeGeeGyUOIxi5Sk0KMq2nkzBYBCCohBlkxh3i+lBJRTCXVBG7E64fx+1zQhg9RnmR5G22UTLSw
fp2yA8M5hGMIkebdkOsY86RzNYECw453oqhmcf7oP3ebMF6KhgFhWnOdJ+X/DJiXNaFGrxcyxrX1
tY46uuiUGxQ/NvKR7afqjOUsEs6uzDYMmRbdzv1apLtmbDsCAmrgVMWeGUps16XWT254ssASCvDS
46rqJ96oDsoF7xshQtAmXX8WQquQmnQmRShXA66hbOtZs14dHw1srXKzS0td7zSWGGuZ4SvO7EyB
1aNJP5tuVIvlkcXkDhSV+yiwpNTSVbMxMJfdEmoP4AfKrg3fKCFj3VO+s02wcxQ21Dd/RadH60Ml
sRUucz5AO0P148VNnKMNllgQ0zkTj+vXhRq4YdD4P9khXbKirmLYC760AROghhY+ftyl238cxStD
8OtimN+c9XtkMyqgqWs/oeiRcPEEs1Ejo4aZ4Rn/7NrrMevfsmpZiKpyOygCZsQH75SrQUQjyGIa
H793bsna3SVlQ44f6AHlsRTGgCMqhyjtI8oIHsrIarcPaAqQy/a2aBsbhfspXV1Gf59P3jkaSvFE
Ef+c6i8DFCjaefmHJrI2Ij3bqBbf8tOeOXpSg13MHzuyIpvDvjRWnw2Mpkdacuzky3E95JBtF0m8
tNJvDe4d9/8EdApcwAj4vGslDtbrwnSR7O1ujaFS9riv2X68fIoy+o0GsSn5ocPCrx2YLzD9/a48
b7Ina1vGZRuReVDo1JOQeaq8WfL2CZlcgnQN6W1ra3OI0OI9wXBDRUcxu+IoU4Q+yY6g5OKTkVv5
LYTAZjd1cDdturjwM1xIgMrXTHOOCFGEdVkEhA6bsf3Z80lo4TJZeg8J0y9qTiXuPHLj4xdHFXnA
sn+H1js97VB1eEOigy09pg1d4d7Rr0dtnqypy5dHSrBOCC7OqjhmvdlXZ/cuB422zKu4DP+lENzg
tBKSFCcIS/HVguz36YHpga5upnCBy7ug6x9HKPgfWRuKi1kvEcXxEc+8oc1M4+/hNX9Y6Z4VjJBY
OgolI5aaNHqiLRdu3KyIleZI4kBGeNvBF+jRw1MDsZ1F7dlUytl98mmA5b/C6DW3oS2g+lxre/uC
Hm/hXehG4tUuQj6OcZ0/9WwYgFh8V4Y6IUadFXceianCukVTOXa5YZLDQiRgfUoUFeMKtvIpfB36
PhcUD8e++LBPYeaJXYOC+ISpePVABOqh1BLr1jt7ia4wRfppvzUhxA1yNHQyL9tBn/SenYcJu0PY
dNWYUn5nL/wXeFWmzBtvpOoM2BfVoh4QmE2AwsHsDiXpBuq1TDGOAT24MGZDzsfYQI3TkojdgOFC
FeRS3OCThHKB9af+egLDz9DQSkn8P2yqTAxSHOsziYBssssDqG9s37YGSFGpipraS4cej8/iMIYl
Ug3Frg0F1g4rKgYY9Xet8l9hdpL7EctbTKAswgeUdWq6BbEwY2bHpgXZ86Z2cjPL5Ckk82h8oN5h
NfVjzT03eAC0cckyQnB89wuvQN/znISqCOChsCzWzFws2zYYmoVXGy12T5x6UUyc0/vzI5UXQCJQ
dvyjYLZHlyAAk6P9ajsF9sDleSJiiD1r+p/Qo5DZ3sSqWpMCe0jTdohzntwgWTsOvnOy/RfgscdV
EMKn/7/4CURLlcjnVH13qhp9VDFLepamXS/vZju9ELufsiA2wXHEZ758AT6+sEOb7Y05N87Eb1WI
cqUtjs8pQi+Nuf8N8NeNzS18frZOWY5ZWJyMKWq1jMCOk1cpJPqcQX12A6GyIdkCFEbFgYxpuPeB
ChpxaULFXrdqgqpkt5OxfGWtglRhnzLOvL77C605UqfT2PlBXYfsvZlUEDJipMtbSFICzBpHNa61
+HO7oMQveO5UngRXvMUb4vEMGvlNX74S/gn1vj4Gm55eQp6xuprURepHMJkU8/aDesVS1dfK2LfE
Ts/tyo4HKnk82YaGyxQieV+y6HP/3PP+zzPvxMyOyp0Wn6X8B6aTaOIw731YriDJtMNQVoSjRiE6
SzDDtQVuSK67kvrAz6ySVX6/v1aJNZS23rfOruqsE62DkJLXMFUnTjkmpEMib8h310rD3XBvzvzJ
rThx8d4loe8DryNFiVCKBtYru5CuZtFhXdzuQC7kS7mgaH70Nw9ajxASkdd6dmxuO3IjVPXW/j9t
jn62ETexFAMyqRRgQk6E5kpSJCsc4QsjG3zPGR0zU4C/8db9pwTraP3qGSJ+KkmOQ5w0X1cLmcfE
QOq9d4gUgI4HC18bJ+NtTMJb1jFeBuBxRVwvTPbYmOeD05pV5dPiLwlnb1eZm1uVm7W1rTcrQXbd
Idz+Zrb6xjbEMrifvFsPOS3X+f33H3jRZYaAfBM1kZE4Y12cdxZjd0qtjPW5cw3EaV9cUbZ0asG6
PyfPpLWUOB5UR9XJlDUc1rXffKLw8TzfQR16dj06VmUDzCU/PDoZYja22o7Ip+SKYrpZtbfm3aBi
RN589zm36D8QMGLgXsCs+Wgopf9m+6vokeLIEL1i633aM3O6jcNm8QdLgqUOnmQi5r+AvR2PeECU
R8FVpK7T7PL6gPlp0eNCgKODz8OBmXpsebUho34fuvr/Tz0Q7NyeLFiYN2D3BopKdxBzW2+fP2Xd
8uNgkMbzrRfxK+XoErEx3cH/P12F23ctBs0/DYvfMLgXXZ09wXdvzGnuo2GTdutrpJTvzN/KwTG8
bvOf9OUXQcoc0D4oWmi+DlSO5XvNgJILhVf1sy8IvgzzU7nMMgFDs4Ok7lgWakIwIrctTJXHjGtE
25lCSOQ8zc0CDVxl/PkNiUF+ZYtV6ZzQE2QNr9kDOifupKLW/KRDjAi9FsvXaSnGlGtmzpHNnxQU
s/o1/PHsGXKhA5Ng8Oncp4EE+HfCfRzr7Ke3KyE4zo3gx/kQ2cetrddlyxOCYAF33Q0Gc7eQ8NyP
a1TvGRsmZauNPSw/vigRZKp8GpHstI71UK6/ZfF+We+Kn456FI9py8aVwD1Ir3co/fm4TwKsazFz
64wWxPDHU/NsYhdrLRgcsXr5M++xVh+tCxTxgBRCZYtnSL+tQIKHuOQ/35Cq2MPqGh67iggEeuWx
0eE7SEXb8Xy44lhpOjc3LB65FWs3EpFNbmO/Er/ujktlm24ZH92rjvzPGEW2BRdgPs5zIFdxIkqJ
d5EELoAcTRqQAaItdE3kaYMVRi7dkrloDnGB+QcKRQk52sxD19vBRlvpwFkHlbmzOh+4gsRz/KxN
pXaffqWG+CKYlO28Bl/0vIAgkHSxogEnSdTrtgxhXkMZfwaOirEa5NTTMJRNv9pR4xinqzRuerQ6
5DDLueZk1JT06GthOZPj5ODYxmjUbokigkcni7SnJhIO28St/59fJYFCHAwP7rtsmONIeARpelvq
8v7IqRpz5a1yEw9HAMnfRq1aw46qDmlR+O9MqlMIbhjQ83k7teMRtOKP2v6fnXRwPthAQYkCufLZ
l1M53C8EhVMMX+fwmxL0cB/AFYaHVhBLVJFC7p+hBOlklC4o6AEzqA7CsHgd7L0MerRh4NCrvhnw
ViJ9rxD1BIK6Z09+MFhoZwv1/hQNde352IQPGtO+r/814ChUELSvPUuTLHCDTNYcuhy9uYDMuxQE
c0aXuvOJZuO3H4jaAJOOMUCz7eJ5VNYJti875nyqIZpjdwB9xEBg9BnXrg3DjDeXnpXqVOTG4jdf
uGTiGNzh/t6gJYb26fpr/JdIbsdddyLLORgOr+VIO85ilfMQPwFcP8UQIvR5Nbi9MBZD6CKL5Epf
iSc0ch6EXdNVRXd1meBNDjwCp/7Q9yzy7qWD79SXdyHtLNMd5Wz0Kr38MxEtj/evEWyW/v/Iewv3
r9r0pqtcx8qT8KKu1RUkqhZPd7eol/+MrobY3s0cR2ggCN7oyapqn8XERS0YHjJIVQ8Az6zBdePX
eDBYzgcOIatqb+dEW0yCpmKPvt6R1hrSR+rSI4PSsAEw6Vb8FfGm9kcWx3qzNoAUkNXnS49P7lZY
qeindqTeArTVByXkI9x21Qpyo3OZNohMENGw6fQenreaSqsN0nxdv7d24JAMoS/C4554pmLdkjtk
uwtHdueH+UXlOvR6TQCXxZ+KS2MvewIhkhx1R1DmR8reOiA50bOcJwPkTLMr4Rfzw0LHpUrQZ8U/
3+u5A87GCEM14GUjzb0TfnPUMQio5AGBF9Zz8A8NHRUoP14dEQ3oh/JDgbpTqAmugfx7i5WWlDm+
b8hS01ewX+sAdmEAKrNZLOirVKqOmuhD8oeISjlfu1EGhQrP/0+oD0ayipKYV3XD6MPzlEwybqKE
OGEqJM8BnD5K8hAchMW+4F7emp1cQjPwDSoENMRr5qJfUZcgj6FNbqF52uo5ZR2kX3/tcpZS0I66
zj70P/Hcx/zS4rcT6QPpdbreM2JIDiFbRoNvF3pp8F80QKaiuX1fTHWv08+FlG0kg/dzCfGbjWYn
IGpA9OBqM8AIkT4GrMT+KY6A2fnpBLMMuLL1V2bpBIIn+MP13+pUDOjkV8DbKtw1j9+MrIMg01Kh
yXIZKinBl8RCl4TDQvkwBxEWLna1hzJpp9jf/V1eYA2FURbSu/XxZyCS/UvXIxB7rhEN41Chid6x
AMCcaBHXdSwTcYZ8qAd/exPlheXYn5VI61Pep/q7yduUjk0HXIZOdZC1xnQN/xqb90Qlb9RXuQR7
6wmgjRlke6X6l7qfOPitldlfenFiSrhghHyIW17RwozKerkF/VDRVi1SCoBRUC4MbJmNvlHudfXj
qgoIg2mnGe+K2TfSU1DQ5ZT+kjBucUEEqnLcAjKYqJmo31/Q2fb9sIrLpx5UFbcaOjeTFLx0kHRt
ADMyWP50ggTfdvPgmB+dQWJgmp6rWLvd6xE4jd0PqH2IHzS/hV/eCb6nW+6khEW2v/BDEegCK/3L
oJ9bgaAspTt+nHPz29QO0qpTvzjy79GTT0/5iwUXJ8l2hp5wNnjsts3aDHgjPc+WxqenJG6yTn14
Nx+/4hNPj1RTCmq+uD8/wzpB+4BTuIeWdCdMDrviDpr5Tnjb+NoHCBzLpxIBt4DUoGOF/sUQ8heC
FOGM+tmCcjvywxC+uUez+VNRUORO5+Nj10ZXYrcOGymCGwx5Gsve+Ft6FUcbuhT2UvwwQZ7qMyHV
qQAtNgFqcLE5ADTmp7E1r1Xj9B9dwYxo6ZctQSMPj4+MhbUJYoIOhmq0bYx3uw/CtxvE3Uan++US
u7R+uJaHbpDEHe/vhbbXG03ul7pCmuEiZ871vOvudVF645HUWtIrcPaLv6N4HXvmX6pam4q38mlG
IZjd5hEVPDBhOqNpZJ2GZvqayue8L6w/yA0Of0ncayr8EqxSbe6pk3O+/AVhCzFyamEgw0iKO2am
+2k4QQV/UN2Q7Fyo85H6fpNEQANhhfhNwn4k81qxPMITg2LJWFJdh+t+WtmYqpXAsYub8F/9dq/J
TpoKJpEvarevYpOr+1Tr17F50Qno9OZ12gDMAdVs78dc4x0M2UpaM2DWlOYhoan6tcx7ayKP9xLX
cBZjgWS6O3wl8I/nPVVuQhU41vUKA56Zbc1PdreO55J+kd0vv2EeSgSf/H6Xv2uq8Jm63FHEQlml
6skhScOesP17bxa6wWQ6wjVBvmnAsNJOoIF/V0ReUqhgduErZLZ9hR/o7MUzf2QjqUpuT5GkswOJ
smGT8aq74O8gwACMsq3YfMZw2fUWxIizWlrQt6V007oi4AT+P+lLP35C0s7y9h9KPixU2l+Q3SDa
iRV26E3VdmYFlyscJdoXqW7/xqNHry2L5lxYpxQkKpiIO+0L35dvewQY0pfbUOOKPeoauKiV4qlO
tro0mdO5klvHDX5nHXm+LJE7cfxXHXhCa/xauo1IKI6alA1OtmMveiCZadH5e2gWn98zDzFHcjG+
siBqdonZAprkvfJ27ChGkVQhgs4yMdyyRKEqVxlPrJAHOvlaxCn5rkwg08zjOC9M9HJ3w0vHrwix
WzBcI/WeVVP/uDOP0wRnpAUXsU2wbXyFT1yo4lgMWwJX25qjew9/zwtH8K+HYjGTnqycxREKspoj
aIH8UOylz5IpzQq99/2rK1nmxlxCXsOO52V443B+76sOE9NulgjRdK2fZDVdQpIAGJzURV7yjPtj
dFkq4pbzkbElOadHfchrFrs/HLJu+NN8N1+iTHnPpP8/JrJDoZbotGYSbMk1yH/Tq9tkR4AiYM7m
EmCmarHeWj7o/oLYa5JqjyAXVv6MrPCriCl/hwCurLrgd/vt4cBzLR9a1/zrcg+eiPMLn5PAogjK
rkgSPT3G14KeLX5iMeitwCQumSs3VMsxpum0qys83qHYlck7bhD0d1ihZdvNHQilyHKHJLEZUMBs
mir/dmrc6v+9gfMzS4kLHlUc7EbJ7hE9dhXBaFNVRBwHuuM3M14wytIzyxGTRxGd4l4yr49qsUjm
XkJsUlyzrCo4xSlHPID3wLGiIAxpf+dh68kPnJMZgFBljyHujDuJCkpccVvVMeaMX3hCMnDq9Bav
bK5hk9lBzOxZHZn5IV1Exmaeht5Ul1jPpT7M3+MOKqaLNr/Rej5IG/pG5T2XpKbHg1Ff6atAVXEd
2olSdR263Efk+CTMD0xGQTUmdITO3C5PBRbIZi160bVjEqoMcu6pTRsMxfbMM5xL7DWAi930NLCz
cHKiYT0wPjQ2vL1HQ5t+e9yKaLPNZ/7Q/YNhxbJrTjPI7kWypFtUGOpkWbCoAaXyzGBVNaWaTcqx
aaPeulwUE/+v8VkVIV3QB+U5KELKNz4b+LUTYtUFuW6BKeLrHPLaz0gwVZnyNMHZjErwfIQUmYr0
IhTxXQFCM1bC1eZw65Go+FdSeIeeut8JlJ23vh5L4dwvuo2+Nys+v9fcwD5gYqdMi2ILyouFmso2
J2VulUwXOzZ+0VN0weGrTxRpnnMRO4QgtSALegEt8+QY67FJUzs2oCeC7NBjByUhVpH6crXffJ2q
Gwh0wXHdhAB0lQuBZKVLXa50BhcGzK0hgLIxwkd/FoeZPNIJK33uV+/i51Re4gD767jfiRbbz7I5
93ZmiTmothHH/1vJnO3n9AoYpOUtL8vGNqhufiOu5kxvIcT5StDWPEWdrDLal85DI5aICAolRkJq
rwFq5CKezUhanltrlfedpvhQhs5O7IaDJKQRAgcysjw+GZTgzpvB2HY/BZFou1MBUUlUtgvhLOd8
jC9Gw41moszz3Yi36Dho6mKNVoQmvZ2jFloMPo0ubZbc01fJP/J+MUpc1V57KmCjaA7poEnJ/l5i
Jj/mTHNABzHh+pweWtR1Ntx13VcGjpxkHDJ3WYJBAJomz+hchy/wTmieLVUbgoxWPslsHiBD86VK
Or/FDT7hFIhu/58atb9+T+1KgqjJdPhsXUtXkXr72PrnphTtV0gG4cb/928JtJSZxTJeAaggJ20P
3Ipo0FQ/e6/MbpkgiGb1o309jatE2ztrKoauUEFo0ySIUW/2poT9LN8YsfvRUDVXys5xGeIjuISo
pn1u3zKR4chgIJ/7caw85QCm43FrJ52InNjr9jhocbhFLYz7EimafP9HrZt4+nqbsf6qdmLC9i9Z
8fpAwxDAH8c0HUrn6pIbQtJLlhOpoEYaYRKrZ9msZpmxk2RX/t2Gqp1H0/yss4JYAxGej2HGCTiu
zpbG3XHghoi/cEzv1G0YaOKswIVCm988iKA2cSKgxbciEtzmyhKWqHkCgTB8G9ecvUTjc7KithCd
1FaaBCByXrNxVjfiFnKiLgouSDCL1wrOSG4NCrPtYYmu1jhYAkM42YYL73qmly3Q+h7C2ERzCFd4
iwz2VWp+OTPyQYzek5nMO/lJwjboLWBbw2AkYB3kH9jxdFXYH0hd9AAE+kl4I4clV1BUJr1eSNrr
qAZhM4jpIC3pf6ALZF8r8RwUFBB90XUtuscyaxEbX8vWsZsma1EznolcHUMdE6gt6hmZVlasLcAj
QUn5kBKMnO65iRSpT1m1TLhts9juSmy89Z28qHukuoKYmmvbDjji9pravuEB2HzqIEN2gMKjzjFn
UHYSqh8Dc65buCS8kadS45iWERT2Ri6VrNdknfpRpRaq4qujcn6WEMIL6Z54sz1xKHeW7zO4K7lU
wATgyd27uN4Z2233if9Mp98hHAONRRobTIPBLgz/gbw+P1myhqmPdhDtbetObYmLDm3zxfW9853s
zaIWCeIrTvApo/irpUO13mzYrHX6KhXt3vP+L0Nm02gavwBaUOD+uWR7Scg1D06gq4U+5JRxAIQF
2uqDtR5Nw7uCKiDecu9dprJcuREkqrc8QK9+/FxM7uBLDJ7jqWhIyUewJ3WXEFBJfAwIBHEHjS4k
2ZuK1RuUlT8b+iA97upnQ96BCmkp/SYZyeAEBvTfKSBy59ehfFwra3ImmeOktJxXN3NLemX7Ovo0
6RBjRSuJRtX9BTJsUlhxxf/O3ExxoUira+VsEHc/UO0ktLBVzFe044dT3h9mjzAjJ+kGPsZ5vIzV
AMe5L8E1vooCaGOxg2kc6arZL5RcL3DfIkj1cpPI2dCOmlWkL1iqLuc0JTIg13EWjzxqA1CmLK+5
utbfOBgEho1CSFVibuthr9oEjeGsd8n/JDH4U7Qvmw5ypr5KzOKTZ0YYHAJM4vetIUsOotOgNBd0
elP9YKLs452/ls87hPgT+AgHsp0LZNIbn4s537NIyj2ujXG0meEeQRU/MJTGg3znD2+y9D2FsEeX
/UtUNfBxNqw/5JmDOzmwck/WC43lL+JEHj0Jva9cSJYxkJCXVJpFrj2v93Zk9poBzuopX1LYIYMZ
C462tKrAuAiBf3BUvzU1+J39oT/uLABZWjKqIbzzZWl6QwGaaoSmWwCfD+WQZUy2IRDXQ99OR5o6
VpnsOCPbN/wgBPMaYdkHVbs4275g91NjGASV3Uoge8Qi3MYn7mk+wABAgYBoupVes9mGqU4KhR2o
vJuq3ILysvTMvNL8oBUnh7n2o18fmHcGgP2e2GeGtwMwGj9Xanc2KSvoFBL34jXd2Z5Af+gkpVMS
nnZiAw5YwHBhyhYsffiz0v0mme+PlaxkrlR5dInijByyXHXkt35tQoyqTZPRjCerOl0+ejQrXJae
TyIooqpypOeVTSjtehcxOtpoGJFiTcyE6Lx4hC9m1BxgJTtqxWtFwKoiSpGjWg9SN2wrVFCseSOA
Vv2dqLOwNKNwX/7gBVu1x59ceVcFfpqtR5gr98z9VvPcNgUCNVElC1hzMEaS1HK7wRKb2qxm3ZdA
rd7kkLJHOX95lLmm8nSXThsIQUI/UjcqjqdiYCbsy6xRfricoWJGa7Yd8xhuwefAnz0NXeAV5Z7C
ftRGc3UAOnXvJ2rY7TGkP4lh8pF/c91/Px4MNThiFkdqqFeFVz37lC9owexyelQPoUhkB9tjJJyu
CSF+V9UV5tniGS59CYw93V4wWTTHb+AL+pAlnvQGCaYHL+Z2JYDAt/8tBRMOq7efeXVW0yLCaGfE
RFet21BefVgxeH5PFNUjR944pDU7CnsDg4u6tOFUEpbpJ1MQQ5mPY6d/tLoyaP6ddLYo4PXG4BRk
7wKsRgappKo+xzufmMevPttRd9PgZRdL9/ZQETV27fEt11/8fb36kwJQt+6WwX95de1hhsrG9K7v
JzDwuPBMXokMQOW8F1//Nw/ZqV7C86PQOdcM1OWTTW8NRy3Dsa3u3nK5R3IqqxUn46eAoN7BBAOA
8gdjMukevU38/zlHucK0hfuHUT4LtCevMryGRTY0WB8dKcUQ3TZuQmf8f4rZUGs2bFlANzOyBkNX
7OqiF5qWWc7q9KzpXtlWFrTbFAWA78aBmkWUdg48APKKFNys/a7GlOVczojSEZ0ltEvespKzQRAk
v8Qx83Mh+w04l7wQMBVQ6E6JJ9uRCsp0TOyiFv4vgyBzYX3fsNnsfw2s6ch45oXNJHOQY4yml0i1
aAHWPtFSOYLbemBDoOmPUs4pMJ2ZhhaQ1F15zzQB6Zbk+LZhUAhDmBSxmhNvkJaypuKscOuyQKJk
nv2cm4Tf9hIPXxl/RAOzcdV8Ceib6UsYepa5McbYVoUb6kiMQjRhHUI75U7xxS1UpW44HpVNmj4+
8AfV9ZlYA3OuRTJ6BHltKzEZWDKSxM9F4xrZdbosqa6IB4OZ5YY4fV3mvaibWdsQ+0/aKUCGnbnz
O1jGHPLFepukUnl+ME+6E7z4e2U35qvPaw5ebuHEGSWLc+ZmoGRwwsyt8QZtqxylguVC5Y8EI6t7
B096xbYPwhb+FUh+gv6sWti9lWJBlrB5X0C62wH1EeTSVZNcqpwujX6v2URv6JipN7RD5PL8hxiS
kP8shx519qYoB6/nbdWfhZO9G3XgDbfn6t3CoUlIHDLL5WYN2gNLKClHkXCT7oiTd7NO1WlkwJFH
8ifrgmcPQHsELukTFeetuHIyNa0iYx1oQn3TNNoFr2ZMrr3H5QCwG07mUiT48vawElfSc6JjyFOE
D8rHTdi9iOY3n2sxw0hL6AVinaXe5GfbN9c+Ric5hST+RtA0gH92xd68W6wh4ECr8DMwlU74H0v0
SyY7NN5ZEEuFQDZZjdpOg1SSBI6palR+KoOwbdr5U18MgKUXT93EMN2bdGeFsLueHLC8xUiKRyrU
tpDvgj+oRvIkBp5or0HNlrH6Z0QFxiw38nwG/JW4haSgyMeCe81Z69xhLXwzsFSbMMrY/v3A+mjn
BluZP/vh77SuyYl5+4aIL5oiKtav7r+9Br8tVo9Ccqodu2txPtHV3CCH4ZSOcY8n7zuwXSUNd/fV
i+52f8KI2l0r1EvHLLYW7GSuvgnRApWFDSoEreOg10QQREx7U43vTdkW1wp1/j0ypbiL8Sz4iQrq
R76jd3HtMfrkPt1XNjqvtBKA4ssIPn5ATkVhjI4RHhGPZ82YEI6gGPQ025F5i2IDfrz69+Jdr1TB
B/beu/i21fyGbVesCmTxlz7GUuGsh5995ScpUlZMxobE3GaGU1uL1/bs2CRj1ZhSUvXhR7ykQ9e0
00HBFNcMjEX/tiZw/KF/Iq4mylY53eTlmQylv6qoJzlY1j2hIXQdHa/bk0XimTI+r89JlqKGwqHT
dXy0JkZK98SKYPmXKdCH05SHkYF7bbYrmUq2USKbEOlN/jhvSJUvxr1rTvDEgKCEET8pWbEtto7x
Ar39b6FLSWZ2FrBNF1H8cxFhIlDTH5jJVoqgib2aeAZyUH6mjPcuntCc7ZDOg/n3FXS6Na+erYoX
NRHa1LYlZ2hpDeuCnUVZdvNXvWjD6RwDLnQ6UBkI2NLakBf56esG+4tJKlAuxRdtj5YIG82ruYT4
eUsfPnLOXP+VAjP0eDAI5Vn0z0nt7EbRGkM+D5o6U8eKXfHyW74VvoMaYiNDe8UTBncAm3WlsXB1
8EC/mJHSanZ9HuUtzDIwzTUjq+M1D29mUSgVlgoM58M0UhUIbUuklGpcZ+b10DAruY3r1fd1gUP7
PLGnoyx4m/wmWFJ+YxRHudktRtBIKg8iSrUY0My/Y8rA0xxQaFmoPK/TkW+DElAMBvfXMwgDH7XX
Re9UAt+L9SClJIdnafVihdIdRlcrhnaildw1XHZaXqdWQjqD5PmwleXNX79T3Q0kX5fXAl43Mhwr
5br/9n46dJlzLC0hNRHUnmENkOoltIN7ipCVoOUe+D8AqzmQ3fDqxn7sfjSbDjGZaFRR0KAVuRd+
zQaZadzY7x/ts/Qb8KatqeB1AUe+5EkAi8Eq80FUkx0fWSNijVTlq3FMZEuM1Vf0RDRbjBTSZU3k
8GycnDQkpKNF2/H9rRK6FKek9OfuxQQdgAuX2lSzkD6FKlbMa0L4Fs4ZCLWEyWL2HtwFhfaodQeK
oT+WIo8up3OGqXb6p2zdFiV3Q4oEFmlyF/JjDZtejXI5jqlfNXHHdkIroa/jbVs+tH9eB/VqNpxj
l1Y+wGUUrdOvjH4OS0NALOG41co7u0/V5fPwjfgycMFz+jjH9bU1GToPD1PZgUOYI6BFpPJEPzEh
AElGh7jcaluVbsp6AbmYCkVjotlhypeiX47qMDt3B5fV9anX3fRpz27xt/kUPRBwizqSUI4R2RSl
INPEPif9qnR5Y7AU32y5PS/QKWd6S7srOpL5rP3F/O3OqhQTmN+i3Lh8EnuLGhdydMuhDnNSrF/l
tBjzVyvb5qwG1pk+CWHILGe3dsRN8GMMFNNbvwb/q2lOtwjzsliJg3QOr1qWpIZZsb8s2pNePwVR
kRO2pkppO2mUJ7Y+2uZMOYELJfml9/msnt2BtOlue45PnGmobTpH/8PoD2lrJbX0ZRSKkHvsrM0C
fYSax5ST4V/oRxslBoqYuSx23466qcs7s+gtbG5BneQPD5AzLmMt9Objo9pzmVKolcUI+6jMvZyM
QR+UqzxZHC7sFPbZq2lfzE9gf6hErQKdqodm9ye9czmY+16NszQQwim2uItHX5XKUy7jnm8C/zLa
9z+TQ+KJt6q5lU8SbuCwIaJxQe8U4x+X/0uEsTlWxsJGnBFEGG+v8+PErceLYKyL68rf9jYXtZUG
nblRBpSwqikMibQ37x/PUNXDqwqcFR4pDDjUDt7QHh62PSysWB2TW1r1uE/0KjjIETPwsMmJGFsw
hG3sQY1fdlWS3jbqKTd46HXNqBcLSFlx+QHkvDNa2qWWi6YRS0jryqCQhrXqNKavDstdm87/sIR2
1xc7jwRrSs7wqAhw5r6SV60g050JsIdOwNl0xtN4Lrdq3AmXGjXSc2IaAhnfE/U0KQ/dWGdJMcob
YedVP5ouc3VXOEDphElYZWf+RhlBG4PF7Ezr2bAkGKq+zANeSlTJR/ANWw3zIvNimVhh+jzZA/5p
LyqdeoONd/w9pe/69UMokP1AOA/1UOuiBMysfirN6juA3StEQe/bViz3DPl9jiXJqD/cj9ABA0BB
wn5eZNOZv9NMMs9XHgqAmmHVunmbxvWElOI4kL61RL0sbxKHW3vTJVZMThQTyz1Qw5ikYAGCbvW/
0X88gLM5IbIHn1pz4PykbKYNxxCjsyej6RfoIt99GD/zeUzvERenfKm05Vqon/RN2Yaar3tCl64y
04QH0Pjs+/kzcR4IIhPQjPElax/wZsvl0ozbnE03QhiM4qGFTnekp2AR4w/pEsJW1D7KKp5RRf9G
ZnWPesvRMfnXluKco6Fjb8xWGigj+ekXw23gUR2/L2h6vD/ZuB7wpd7oEO7cA1zUC1tBBkr9/GGB
NhgAjlZNQYiGUpNBAKRoTuJpPhS3La6TXIfTtjefoxLKPSRpU7lnYv4/LJ4ous0CHSpaKeJ2/NZA
sFaed6Z0A/cNBdLJM4rmOYMPe3E0E6xboPuP8/OLRxW6U8kq1MjgxAxM6G3SaVMsvUQg77i8x0j3
oPQuV/RljMVIw19tacCmsgTrxBSsb/Kzu/+yiK02jx/cVeeAYp9TcujXbd36BC8qosf6SLkJnPgW
c00a1ulnlYNJ92aW4cDXqKzML7mgknBgesiz9p4Ha9+dAu6Mh/QlEQTe3kE6xbtDsnkDBCqDm7zD
TaHG4xephFHIDX9yvoV+ax+PisiYnIlnz6xYa9pCqnFtiQTv0MAouQ4rJai0x3TsqGTNqz6kBXMs
bKlpOTWoCGL/hpTQy20J2SDXFD5KJ3fMZMCUIZbn6Q6dMxf1ZTQOtseteK8dsWQ+gw4s4pvS6+ak
IByDrq17NnP+Pg9aA+ToqabbDwN4rrw49+dYA6+hsAjnBI0ooFYldwrZ7rf+8gfQ0bSXa32+Tzlo
NRFXm1ul7vedjRM8bHMqGaojmEwESTMNRXJaakZw5PzhfcG8D7JMeb2canCO4A+vKpfSJSYHPHa0
9Cr/VdA29MdJ5Xde0vzTyfeUPywUVnf1k629ybL4XRVbxUG5DpalSgL9yoMEiEIb3hOT3ub0Q/90
rvERcjCbdhq2NxDlQexdneREyg14lcZK+UXvTgbDF4QHeduxIJaSUNZtJU0fLVpkU7HLlxdH6v7E
FiiLiMHIW3w7Uh0rr/V2hSOMOCupWyoQvhGPNLCOseifExuNi5FgPSi5J/fGanJTZp6gD+RdqdSf
PR/To/3HwIN2LKYuwGd3CJG9fc8/1GyAjIZT7EDDyfxBkoirviSHPRsRk3l31ih5YgvCWU6RdFNj
c7ZevuyIRu6Eu22PEp9zkJ2q1+o/SDhKjC7tHlyNx1q+MJ7bh7KQpzhnX/8dLn9h8p9aOjw/lGfb
nw+tsv/DJNTd9I0kpz63BsUFSQvPk7sYVD9quqy5p6Ih1LCDHIH2DqegggmyjhcFC8NKDiLLJnw6
/tk00F6nrLdrT63xV8MxgIa6q2/iCUzdHjaDGuJI2YqlPqbzg+kpbAwQYaP5JjNsp0JpHnr/rbDY
ThkVBUsN0LJniGGZdzsA27TGlDLs92MqPolCitsj/2KnnX7KPmsrnoijOL87tv9REFdnl5WHXieS
u3VDkq7AowZ8fPw6iSaEdTeCn+qiafdb7QRxNPb5bumfMx4aepaXEoUKG+M/CLKdvuwoBuuXD4Wt
hJOri7jQjMEEwHd0nNiIsdRPOFx6wKrGzYckQryv5+NPEdNUwX0BAvrf2ioaeeYrsuly/a0guU6W
w6WJswwk51P+/Tbx5iOmVhkInYiRg6+EMr77hxqGN/tEjopJA86XzEx4hutT4JzCsHGrOgucxPZL
2aGB7hZX/K+tMaInc7ix7vb+TyjdkegyE5AyOWBqcNBXcPRxoaFANxWhlDAXKfjiTp94sokRh441
eZTNN237RA2miu04MuIN18/6lGygGNDpUWYz23OwhxqjI+htprrps+mK8LMuI46qcjt6DVJ1Rsg7
8g11K9j46di/jCFjQJcLo1+tN4qnHrt959HIZFlyl1Hp1WEdJ0QoxdPMjQ8nk9rOlrfwrAehLD8Y
TXuiiGKhlmSPpUsr9ljdP42a+5p9IpOTwiheDLGQUa92hjimZ9wa3gKYPDj6Q3P/JH7eIfZQxBSn
M+DFpucmaBLbIicYS81SXCr57AiNieQN/WDPTICb/UbZID3m5HdjSZzrGyls2hetcZokLGM5n9t4
TfIr0cbZhWuRV+/YSHGfaHaC4WYhYGtUG9poKhLJjKL5nS0ii+g4TMciXLbb7r/60DM8RQmFjoen
+q6B+Q1ZCuoLsGkwmptHb86DC4L2oKB0aF3PA6rVMSfki4Qn/jWdQOq87Boj9jC6syvhI3f6oZkC
l3I4vSn2NziLiY/Bg9C9hxSIvllIKUlqVBT0KYtzTSQF4m63nKtExleaK4mjuURSCpCiIncZTT1s
wp3rHoB2PmXxREcmxGP+BvU7cHuET+ePieQ4mEI2oqCOUuws1PSvjEXWSHpLZ9Y9SG9vn2Ecbiig
zFtSvUEbZ1HdQTsj2Zq66OcH3mhlHH8EJzaCGbedrZZaqdXv7Eyt6pethyJFJcOT90zwYuD2wei7
Ms6G/x9Wj4lYpOV8xFOWXqNXQnAnvrC+I5OO1cBehoP8ZyzPRdOBWnqiFiwRc+HW4ypScrMVbiFf
MOM0DgOJv88OG74NNp2undMZhbMOlyCuUpFy3J2kWXW82+NQJOdct8Z5OTXMPRodloqyPcoOXLeq
OUi4FciEHMgiEN/cF82gWILxCAyuPAWrraehtT0kOFbnlp3UqLiyz33pFNX6ZMdfgsvr8BrZZxQZ
CLWCRgtIm1GKUn5ZhGhBr1HHJeKNGres9XgFb8h6SIIGAtF1XyuM2I90Qp6QuMxc9Vh5uS3MLFie
iiXlQRajRhd/qUVlZ07OVc/GSsq26VuzBgMHaL7ixnn5M1GYIb6/4qfLk3IVF8CNtT120c2oHhhD
7ntNqE+3AKpZ1uNHd2m1fp1u5zAyDLEnSCSTw+qZuxCvr40ncJ82/+1VptLonjS5c0ToeFlA7Ns7
SWraA1RMNB/c68M64dkKo3puzE1o/BsFMg8StQiz5+vOJuZieoHV94I62JjViHJ5nxIiqdBsKmQ+
qr/eKBFatkK9MoKO5LphKJ1s5cakcLY8+M5Y6hB36dPjZElJMhAquIP+dSlrzom0P6JGieu7cQpi
BREoMLParE93kwuFQaA3yUPv+ExglfkqckO6ye8Yz5oj0qH/WQbJEaufv4f2lugY7pw0E33/OU8O
OAyOoUb+tHqelCmmOgu2WvBSlsZ2AcDIFGwhSjlzJCNDvgpo4C5bFBcAIlfdZUE1Ea1NI21WCDOi
gadwH6y6EZGs54gCAchQ2jYk1rLoutU1DXa5iQrmWleXrOooEpb6OnprUjO6gBUh3dTJY6uB8jU8
bUANM6MjHCuel+hP77DyV6hJ3kBWoTD2cCjqiZ7NUjhqcE8lQrHDhfRyLTC9VloSrqTvccIliyEs
heCpSuv3wB0hoFTWg6Xz/xaOw5TFgvQtObB3mCsENo449414CMZhkAV4pjYSL9gUmTIpOW+QiPq6
ThUCMGJAqwOVx9AMHJ/51/1WWbMobSFLYUHcW2gn/yyBGyTJQeVhntdJ7Fmlhf7rpnV8Q62yq4zJ
MVqIkYDM32DGoGKQ976mNGNWtWSijs6StE3xJf6fCjfdBABEV9mtSDRgu7KIJfKJaAJJEVBkNYg1
i8gL0Ld/8SroylJ5NsLoPTHVZQYX93g42KSVbHnPF4wqfs/cdMh3xtOZhINzsUbiKlRd7eMX2LbX
3IVShOtWIiFexE6K9JvhGH+h8VH4IwFgyJxcZNDLmhCnVI8w3/qoFKA7VTws385VR5e9SVr6mDux
FduHiuHgPks6fHMi+0EoxKGqlbRqLuLcxn9zxS6RN85ypD7muz2y/KM7tlHbd1/lpU9Z/Waqm032
YKDGX5LWVYhThWlU0kqy4fLCx3g+iTE3IrN8UoRGX5BIFvFNTkXfvxO+rLlisdfUaEGbA18TXn+k
JpZGcdcJvpL7xj9tfFvix4AlLbtJVsxZrPt7aUubN9B4wM21qWxx5N4+sFxA5cY10qeEXR/raT5i
lraWlmufU98arprPUVtp6XxoExD+YmLuDJ9Engup3qyA4Ndmzr6pO5VOfwi+817idgDQy/PHQ/Ai
QtnrdAZ7uMjQESgmGTVFnKEE4qCDD3H6gka4lRLFn2s8ifypme5gnGVAbzUQaAyOLNn/CmgSjlkw
fpR+pxgm1378NyPkr089tBpkXOjyLiQ/OBpW1lW1l6BwqB7mOPfLTqJZehUpLIicJN9HiBzWcM2/
MUELODvo1K6gkF+766UePfdTjq8PuHuUtdbewsiNjJme4HYmV0FYUCUWMgXjlQ61mCiOUD68Uw42
bWySZKsekytMdPm9sra1w0klMqT2K35Y03RXdTjuZMKkfeiNMiUK/VS2jSzAr4NWrWRSgWu4EsPS
stCt0XGVfKr+5ss9BcbIbIb24nqMNnmQiwuw3zcwHD5MUqCeE1qxscWh9dapiFyOAsuJzT0v2NP1
ViSgaVGPIrCFOC87HIp018OpXMJTR47CqqkWDW74SKA9pIUhtLj1CRH6hJm/ME555WpfmAFpdhra
tkaypopAtvSLkkNowl+ciB/Jh1y5sX8mA43WTpDfxe+7bBrE4BwI6fCe24dB6Ckh1ulZlK65Towe
nPernjkPdYFtrRgIpuI9ywGjElGTqTtq4diI05xpmSdR/Zi+oycDez26gdJDH6jZyKppy+6/qERf
SWMCh0SP2OXmF6HO7HEwY6fDjHhAS0hDIYb2qIRyWCgxGVSxq4tZSKKCK4MIHUXsxFpt9Z0vGBnV
NaD+VfLtg6a9mavAz+7oUA3XDZdllfi63ZpAr+ao3MvCYyQ6HNI+YMFtKT7US5CJf796W18O8f+i
D2a5+nX5LT+uXemhgZ3t8Ab2jtpXcOe4wwBMrkb/+6QhVx1XhvpN1i6bl5AVfUfua8ZqhfOwDMnv
ow+Qe+tDz1rO+uFLQPqisELaJMDtbsv/OtS5aHXgEfdUcJ/bQWW1ZrmHgBJz1+M/TSdn9vTbp7ty
15rK24w2FALce31xRK3HirrBaBOuzikDNks55TNQhZsYxB41Y1MrixJJFrq9Uk7L5XXrLVGGPa3V
hl3j9+Pe6AAv89AOXf+/VqkG5o/7fgnusQ82bBJb3aq1QaaG6DJ++53XhyzQz/dm4KhNw0XOXC5C
I2EJNDYWCQxdD0Kj2ifRMl9CAehlrbq4Hr8XGhLk9/piwogKXU4N5n3GyjaZ743mBnF+bD/YrC8K
GUCjsm3qmhOCEZdZy+ERkFMUpjCCco+JKzvtDcY93euUopV2inUMDQw6bqZbltRKIdI9N14wy3YW
KEknhSNZqyEeAxodxnb3tuUqIg+L0k1ZPAUeXDY7IITIOTUFNeeb9GdsAprYvBBcRQvq+PRVCZaO
XG/BaHomohSTtVoLmVRp0drPXT2kFQ/khNRxNfqLwke7OdYiD9ULOSCKDt4ktzPSi6lw8m6Rmmnu
XSsNpbQ6zfsArYKjwQTMN7rflq9vbO4V0q52XV4lYmWK535DnxCyBxvh/ZY853QcWu3zqrTjcaQ2
ScTtJeluulbCKg5CkBIz3+soVvyZkKfm74U3iJOVZjhDRp4zR6bLpyk0wCrPK2p9jw1OMCE9RjjC
xpNhLIyvGKK2+KMuWPd9lYaH88Ko0pzA963hYQBW9aGEqa/y5w2XQRYt9fxKSx0PY6BOrTbDNtVJ
HP1GQhE8qWvvid00IzBG92T8eY4PPtVgL+jHxjkd5YPRiYQpd6VktRGf2XV8NRXjj0HbUIr3a2us
QGtifyaMYKIhRSFJVb4t8Ow9pRaZ0PkGi5fGpBAxjvTl4QxnLCTebKtollouqmS7Tjz6qjl5e3RS
n1Wyv7rjz2sHH1hOhzrbeGn5w3TqziKbQCFLH8JU/x7dH7aZK1yfPuhZq7J8Nn9O0WyvTf+DXuD9
QU08JWKX++zoa0V3Y7WTgnT8seVydGvXN6usIbGDQZ3Jopv1vv2EYWeuj2ryK2vqPnC14qzshTEo
uP52QAwVbmJqL0C4XIvsbbJW5D5DoW7qkjKHhZCw0p1FWcWL68SJCvUr8OgD83dGVgCaO2JDDFT+
c3jYOrubMqL0A1cv83IM/d0l8z2JJ1lSx7HZ6zOj8AqxSo50Ar5bzGlRKUG6dL8S1rkiPXGVdAna
vMWy9muDFjJ5SeTVKKQlV5JxXjhiFUNdlPv5D8s74I7juMOc4m0iReoO9XJ3CceyBiUlNQd6XceG
YAizufxzyJzPHqAw0YvH0Y5aS6dQwJzN8bB1LgCNlm0ciXf3MM+KLHUHmIXf3Om78/B8qxIEQZ5v
vEa/zQSBdK6zz3IxozhhTVebNueTbbtpTqFVzfxdXXkukFLCkhWpqB22GF20EhnGoAUuOL0l1Ijg
VFAMlLgf7NhDKKCLbEQRCqI52/CkSZGqqrDZnWFM4VhmTPDImS+FtrK+zYoKSjyOfzwuLu+LcmsU
LfBAJt2fHkdGNLr/Ogvnyaiji4w5qjzcCg9p0YwH1eJHXiWDUGHpziRlxLHVeE0nfoHZuQJUjBmG
gVB0yuwveFQ51LoypDT85dKvBMFtZJByXXdnfMmGvoYaGkaoOdkdn9KGzCV0VlU/MIo3uLBGWz35
j6bN3wY2Svrf+skOCIw1nZc63ZfoYOCmEVUKFSi0Wu3flhWe0d+5ayVMB38Pbt74g6Kk4FVvwEvk
6ydi54uiNmrwCz50HqP009m+5A1SsgFDWub77962l2IGWLHbyT51geTwHtt6M70SFBAEEHOhv9EW
Xx4XHXB67Rgi1ii9eEj8GxmtEEbjNBc5SDtSGXK7bZnveH4W/sUTiIgjy+YJj0b8l6b04N6aGBvQ
7kddcgSXBxiOBh5uf9oz5gvr0dbxxPRBHtixjdx7d+dx1qrSd89Y4d9Gns1Olih9ifsDDXGDYQs0
QDAFrTMPavYWJsH8ydlwnERk9MS3awRBqD5dqAV9ZqV6IcSkIgwcdOHaD62YLWwEVKA6F9j9gOFj
DxIllauX0C1A9PgdhiC/L0mb2/9x8sDyBKE9BMxxhIJuVz/RpQo3CTF/xTPB0Bxa+wNvTyyvHgqZ
2oMvLhRP7rrKVU4ceqQBp8REthtN0sD/rVxUXG1ymwVztiTTLZ9kZ9+k5KjlzLInItX845zWp5Zj
uX6D7wQvCcItPMnztcZISwI/gbgswv8TzXO0gT29ZiAnVAHor6LqdWqtZW+xqM8y4cybA8OAOKZ9
DE51u6eFmtnVBR4EqfcBm5bteV75U6oIfi3z4VtnStS+NBa6Ieol//eLDmD6esG8t6Xa8NXZJt8r
eqQ0tkJ1s/lPaLaKoqHJ6I3Ac34mWAxvagjL0K1OVl8awRaKLFWCl0cs0NTVhiqXX1krkHD/8z8K
Yq4VcUX73fKhiaGq6NJqXV0AM3Wuoxgk7IHuUrx5u+EQ0IJmugZt4QxYer9n1QUdCDY9hGzBwhuz
7f7rjjMbCWnO0C58ydhTd5CNKaTYl0IoaMbjqGWLM+rGZMcCEh4uRDFa1G17JbyhY/yIthhZSx8u
wfMBIFBAHGkReMrRFvOlwM0g2OkqvudB5SfhIMQcWO3bZXqmjdpzCn7xt3Tlmj1fDEmE0ToWjHLe
uhBuHErN2x8Psv/6+l+VbrYYLh7nc6fAVXKMqOFAOsbez1yE2wp+NXPo7bCrFkZ+Avft3+Pt7tX9
OfyDhZHhXgMKYYeHPkscW2gES2ALViqke2iHXEtO2vP5J0qd8Pw7ZNLFmvOR5GiTo1gp4IlQBlw8
8wt3zuxqK9+KARtvQRw/ShesJDzHGRH5G6el1zW3DuI41NtcHx51rydur61+aVi6GTl5KA0SQ+oX
V83euIQ8UxWe5QZH9s7/Uri/AeHy3KxC9K5H6kUdP2dnqkpPiF+5tkj/ZG8QF7/Bj2iSxIPizAAx
y/Rd6zXwHuMSON3r7JnKFwOckYeLjFb3beXMNspbd1mq7fhozwtoprBXJKIx6pdMnME6kX3zxQwU
u/0MNKXguhW/ZmB1ZZ2dNHM+XMYwYU/tfsIUM74cjNDDsXwLf+xJochrFNafHNVAIFVawXsQrw0R
ntQ6kHAu0kgHlS2NZnymVPEd/27A9o2NY4PrXizbACsZczHPcwPl5FYME8Qng/yQS6CtbtKmta5Y
E0wYIED+eoTtrj3bDa0My4qf5pzPp4B3ZYqEUauvmwXPWF3zNDjRto/oLCBjZ/k7AU/Ib9UR9f7Z
F3y4pGKvAbBcSelWX4k/2GpSYoewm/Bpcch9IftBQPh1fjeW3NDhWixZZc4dedKYiAqle29PSN4X
W8ME0+GnFDApM3+7j3DNU52T25RYRY2og7dNT4z9S8ICrVjSAI5sTQVDWc13w2rUIL7pv/ljbfGP
w/ECpwCPEOGSCvUQcGfBFhVCLqVpSijcCPm0HnCD5fnQUieKnaqlzC1mXogHLU97BmLLcmVYBPee
sydH+noLNpFIht4rRV/3QIssFKLR0RQF/WBP8nAg713MHnk4KDLpEakti/97rYK1yDAX2LsHHAJt
0KzUtMgAi6NJLw+P0+t12/T0eqZf6UWEqwlSDBqToPrDtovsifcRATfimejdsh55HGfoOLzdAHG5
/yPDufaAVc9PMlpItHxl1sbVPhHoPWQOieB3HDmnqQsBiptq5jhI1g0AE9N/s4tyXfqNi0yq0lR3
5bD3D5pASfcofyyHZ7VzjcTH1WGNu3UpmtYocbxDlBAg9BY9cR5I/NX1GXj/wxVEAZ9GpfnpY7uY
M4FI/buzI/ttYfMTDEaLmRm3f9Nj85qyxbdBtjUeI0adHjofTvhkLNbFEtyAw4vy+UmWtS6eTY9O
8cmi6dbgyIzS6zk3EcE8khAz5AQbM4a9e/T8yg1IYPJ7OnC1nFrqxD4B2sCO8yGszpUQajaQbo/b
NwZ5ZqXwSdRBDl5evaY3jzUeoBpAcqGnVbkjDGY+NdC2wn8SyF++bCWMJXNCe5GjO9seffoTOJyZ
FKuNZBOmez0lzc58Q+PceEgzqc/pajyRi1jTNySa1r87LBeFnO+rnGFyM0FtGtbq0rJVQF5611rZ
DjK4mx73jn38jzrCTHuuAYuHSAsxKCPXjbuP3vv8VUCnt2u7QAzDNytVqryk/wtTnhTPgZhvsPmC
Q/WCHta2uhGHUMccf9wAgR/x24juVtp5INITdvG/jQ4mKBhNKm7VUlAkXGEoPxHyxVyk6XMOq57Y
6jcxWfj8+8ZZ701szwCvtHQlDw14H8YzHVajKh1YkHTE6qnI89B/V7ekyxW+7WI5ExmHl9gr1N4u
xLgP+FO0XftPx7ALw59FdMfwAooYZ5i1erKrxy/No0ubKgSWXaP0m0PFTE4Un7V5OZv2NVWYMqYd
ztbs1eFz4l87nhNEy2JN+Iu8LZ0a6xR9PElpbU0bnKyfdSPLB8oNGRxLT8lNXF2ggnD+og0Rmojl
NaeOwJPwNq9oy9Qzb0HVUBZcf1BWalXsNHUUa4NwyVOcWltr6YazkrUo/ms1o88tAIA4ulOV3hcT
C3Xwg7caRJe+gJTF8InCzAVRGdw+Ei4j36RE26q7/5VjVcZ06BPFXqGPUZuiqdZoc2wIW/s2d7o6
p6EN+hdjrBRAwGfX9z925S+B4242AsXUgky38HpzSOETE6xuJ7PiD4Mu6fwpAlVHvqLXD10oCE8e
UDZD3THPpijmz+KdTZH47k5G4XoHXBmiZZ/TWqDVNpOzTgKCDKtKHUDGwu/ERgZHWPqMlw/DWS7B
s2I7TbNkopBJCbei4n5pbyaY5TyTAmkChT+EeNEAkswzAr5cExIPLSwcI0GygpBz6qP+/ZaHr+7V
dCkTMxrTfwx5E8Dql9Hz4usJggeCXr2AqiizjFKsN57Tc1byE4Y7eyvEkbr2uR2GRHqn5EG2u69+
QRTZP7I09HJoOJcT9JEZYNlEfIDiAOuUZs6CKw7lQlh4++Zl6CtdbdNXF542HfXXLEupg7aOkBbt
VdcTGj+KUC1Q3CbFZqptRUJNc1YqcTFZT2IGXcsuwSY0Kpnj0j1Jw7vCzTTExmhBiv18BMK0zj9u
3b/ePumry/hjX5pHZolIXbM6X5TDImdoZDZ906tHv4ZobfsNaC4UyT2isV3ml3FZkcc9LzF7LX3g
oGktS0+cQhIHkJvb3erob17Snl1Bysk21E9/nrIHPkhIcWMeV7fD9fSCX+wuhbLHLabY9mioE9zD
I+90fzDnp8wP4G7cUjaG4GMUq6pKwmAX2+CscHOXA95UUBPEO/Wa1PMmlSbO01ZcQyIFNOlBuTcP
OHaYIjgmkIEjauIdBJ1dIPew6l9ghpILbVx6//Y6M8TvXxllXmiUkB6SbXScMubAKAkYtsyrs3/2
+8VU//EURKZf5bvzABNVs6sHmKOFSVb7nkptaMgeve5Jtt75YjUOSRr9ie7fU1Joq+MPOqmdnOvC
MfDT0qqNv/9v01IknwL5UKltSq5mSaiCyIpQuK6YRSYN2Cqclx/Enaqiz5Ia1iccJiUukxi/Gh3X
nMAyxZieBaljz/QaYdkEEmbwssncJpMa5N0QBL3DjX2mFqXRNi8GKXCPeefyMCE5Nlohg8GIJVZS
s4YEdWiQq8G+eeXfP3uxNmpDZa9+5ol+EvKmWCXoxxjYbzE0A01dsBWcbvEUaKwEd3jZilgMHqQx
4BWTanZFWZOKUYxnQAFeN7C6+QY9y8aD2YW++DBIAkuR+nIERFjD5sHt5h6eGVo26wu7xhx+LdY6
AjVV6fbBvdJ2LAHJCJBtATbsaygp5ZjWc55xIUn2UeQLmNxqPwP20BRXMcKjYTteAC1B5V4tVVDj
a55gLfGwYWUtyJTdR4h1KlvptuJgtOfrit6dv1PMMwe7KudZ9HQTUgtGRIvEPfa9YKurA6B6/YQc
mCUKfR3IEKrupTTcupYX4Pj76gmJWc1d4InNxNMcGwOvV8dglR53dfeu7ohUn5qM50OEUMqD61/u
u11Be5aBsvaq9Eq0gz2M2v4OWvJHKDmcbkMb9zXyUEohbp6h5e+YcsA7BiRn3A6e6MCi8SQrdIsA
goAQmfPkJ62TxBsKwrWBlQTu1U4HHfyMxVJJLSBM6QeQj4M6pCAa1LqSyOtjw+jD3Rl++JIJUL0p
27YmR0n9O6Wy7uFRDo+gYa9N+x/sIW0waV2x9DBJtKSh35lNKr2t+rkEbmhB8r7uBiEnBxl6iXGp
/g8NMeXWjUq1KMjsSww45M+QiUOyfcGARSFe5gU5n9yyjsPnWHQpU9yWn+lKpvKJ2FIBhd5QTG/r
VyBLQiE4gsJH8/z6vTwv0APvZjORbxuwdzJ5TZVqDMS5Ig3GvgFIg0QPAjqgevJNmdhPwJlio/T+
EELYN5gYCAm/hur1EJeceynFDh8m79jvJ12+dFO2i7e1XUbd+F36MhnXmJkqrcvXuIlmH/eBqyb4
zBp4QA097+PV/hkr/5Ob7Dvzta3sGMEfK/Zt8hov9tJh3oculYpuRUQokg0sIyDLxFpw3XC/8i/7
X/C0L+JiEeESVXpQGMOCXHBpg2aAlh7Gcif6NB9ihe1yQdt7P67/zsxkGg8cq6rZTudgTEKIN9oL
yw3WjaiBKKYCIqFZ9jTqqzvPMOeju9+X2PcuHKOafKary09CftGk/3/S9bmIOa3at0ET9shX6jc9
txVq+2bp1CRvZr5e0hGMW4XLU8Qdld8beVF1ROTkteOm9bRMWW1D3jx5yBwc8e2sm/IBSwEsSvFL
YK8wlkbY7EDdpmMnOcYhEwYJcBiexmTpwjQcebPVJ8doWHIgP9UjOZt2ye0d6l4R3kCK00cMG0rC
kwrtPQDGoPTiU6N4GyAvMKVAtkETo0WHdC1M1wY9TwpdQ/Y8OFCU2ABpdGD2LXcZ4q+dLQgqj0jM
UOjL3XHjmbpI4PKa+za3MycgAOYO43708/rjpSIw1AYJytt/5xwGycAPAPdxKPR0VsSg34lGoFxL
xT96YcGCqofK59DQnX7gPduC6k5/pHsagfnMbFONsxVvU/EpkPFTIIe8BNAzMAOrPJMuKugf88XP
/hBesZarHl7mQKNP2158mHXKwPg7u5yTAbXBHzQqYEsV9KyyehxY7pamEiRcdALsrBCctV4Az55u
DNyZene8wWhhFOWFEdch4lPS2S8sqF/LHMcelN97+oepAewCHl2mr+9MGMyAuVBZYSd8TAaal/jf
QTWIL0qkxHm3l8jfhpvV7a9nWLc3JkF8egSfrGtTNMG64OXK6n3YPkNPlG1tbiyR9GH53ejDHwOx
EvzjRfPv8tvEPJmkBpgCkSXUdxDOwe++SPxDdgwMAKiRyJwMn/IOYUoPVcduYUylMHiKSsUg/lX1
Cxx7VF5I4CRfkD49jp9X5ZtE8H5oEHmPibjdD0ZI5X9+n35pfr9Lofi16nPSkhdxVeC2GLVlrVaT
jqlr65KkQr7RhMMpkqGVvhqZan1C2wflAplqdNIeMOEtmI3Fr5CuZT3MLSyH8c2ZeizcHq6jRlTE
e5Ih5lUhYSjtN0IDxe4kHX3196lZ5ixy1BV0+7kozpSsLrarHm9Uq8dYfoadjf8DxkIdJcGhRGXE
23RR/GObpYSKRTiY3sLdh6kxPtY4ggMshLf74vtwht3eHN2ItBpVDP70AhAy7OL5FSBuNmmtKN6C
EGL8TOEWq5kx7+zA1fxww5L2zCT46IyicmWa9U7g7le6jt8R47RUhSymKmg5gt+SdFy93zL27plU
QL5rvXQ1wl738Z1wS+ufUs3bNkHpz8/yLu9BV0HbO9Dp2BY730lgZJibL+hMLJtnTxcIEQvlVw8M
/gHluFkBu2FDhGM4wIfhI0Grklcchnx6wRVFjF20Q+AkWFqpxvz1Iyv6DglU9lOSNmOub+Dol4Rp
cOozfCOHSSR6ITX1qeS/bjJMNpycWngYRZWwBND/OVXHqCXyVi3iUU+/rjOyksGkI7mzE8biD5R2
qtIAMwMUVIxHuETjDrI6e23YC5eIj7j2ldneoBH2dqQQa1/VsdtHrrcypY4tTAZljjuV+ZCq35XA
1p4SnGSfxsy7zYM6aVb8a9XOV2ZQL1SaqrVY+2pA1Sfi0hxyqERLo68/z5vYoimJotlC9o/qEzTL
HGWk5mNr7cL5NC9LSSXfTKtV5WY7cCc6+FUUZWMKZ5s8SzxGMxqzFFG1nzCZN9JAGH2vexLwwNoq
d8TwxCjZzYq6ygaGW/dGfDYzw5eYuNCVN129dPEn23ZybTeTfys0wPNqvogpvjoIswb77qDtYs1W
rZV1TRfUQEklONBjXUXEb+mP1wHU4TLFRBZTGdf0247hQ5RpcLxmbW3FfyUFvoJcDZrhl5+kQ1Zp
YW1OXsgPTWfvG+QNUHkUbRV1yvRNQR4TfLKvMAJ2k93lPRU2DdGEMybxLh/ZhmU7Zw/q75FHwAuh
Xif77w+uZYhbSGHE0ej0P18FT+Bsu+VLA813zxYQJRfBzgNe0rkbkvkXv91/7dFdOl7c37/6Motc
/UB92AN4bdNaudm8JDfrm3cwaT03MPuJ5CmEB7VmKZFjV0lmN6BRhzD7GcgaZ+uq1J2P7kytvE5Z
/afg7BBKFstCoR2W9txniZJLTAlc/HvvJ8z4UY0WSORr4A0+KdDVNsiRQQZ6tSXsE7oSKHjrLBrV
h/hHRtNdzzrq5KHTpA0atErpH6VsMjawe8ZuKbGyWSff8VEzke8MNhk41lSWgFhdCve64gZmtujK
lbV+J5W3//S6AAa1LR4pAcS14RSJnoU3jlLtfAAYmkM40/q7FKE2V4v3afGX7PpcBsTCFeyZo2V9
PgUMgCFE3vWIqX38JzsrNWGxWLpopWU/16YcHTJKhxmTtyguZpXk2gRBLD80CXnnbFhmHIGuvyk3
y6tWgO7dVfXt5nIaKeDPn82qCLWButTHcrR0ynhHiDA1luW2HoIfGqhuxFGv5a/ZffD/XEF5VTiD
XLb3Mb1P3ov7IDMKQZaQq0cyMLgAp783SFjLxpyQXboFcYx9fZnrvSEsa0Mcrgt3+tUUN+1Sv7o7
yAxDW9YH88eLSEl2jqDaJgsnHoWpaAhI9KjkeAxifIc2EE1jIqacV/2bLQq2q1+SMc1uWQwjm6lR
WnBJtDtsdtyPlKw+R4S1ut+PuKtKYK7Y21MzcgqKv+D4kdMog4DFlMMWcgmLdlrxqxoxs12UNz/t
pQaALwfXOeRswOLEtP576oM+tMdscJPkolG43j1aDEr/pqAWkzrD7Iwf8djAk4JOslgVj98zCEiE
d4UrsQj9TVwxXY1XlEYuAT0PDFuWe9uNFSvSdlJi4txarDOuUp2oc1FOfv6MRXzdx9gOVMmrP4ys
yZInmf6frLXi3eIaomGALVesUbTXInqtxLhk6PIBAUbuafB4iMMMz3na37Y2Vc58e8x1Ydyn2332
h9cy7UTqoBfBEMEPtx73Sq9nP1r3n9XNinQZ65fdquE00xO6JGlgoSqfj5jJSbUS+9g4DLuasW1H
/Nkb77Ybo0qX5tGfV/Y5AQbAyDeleEE9iHfa2HQXzFMyBXy5Ti+UhQtwN6MFtpG20n2SRhUKrofZ
nT+vCH1NBETMsBcDEaMHNN8MohLpuIdgKU6piyLn5KgujptUc1946NKYgkKJllIxd7lcd3ywj7Rh
WpeHamvtcmjenGGCY8pjyJvd5xKJixIpnt/lWLpbScY0tQ6kMwu29xDUMv3q4ov03G/8Dyut4SYu
/DHaTRNm5QfCuWvKyw9ISuO4S7wkaxpjppXdwCikX9EJWeF8hbfKaSKZP4LiAW0aiLWqidUgXCBw
v5kVYeAQRtJgGy/dAWzNJI1cEHW8suveg8dJaV+CBiSyZo2PNsRALwKxwLIatKnpq5nI9xTN7FZL
eylFcN1u5hsHmxI+xuU2ih7gEe9ygqxoY5ZYYMBDBD8Lugmvu+pG7ACqRJBqE7fjwOmZOhfmeb7T
Mgyb/t49gxTrNBMzGjxwU84TD/heNsSHPuAdJ+oLG9QZHSFiW+XJjp+dhppa6ZAa/AbhrHzkjak8
QPFb/MiQEtakZSVfIEj3qFvMrAFNMhSCPJrF1XN4OHCmYf3wvP5BVfnPnTfzkaIqzyJAYCyW0TdY
uu7uSL8hS2yWLGuOxf+oHQJpReeSzM1JJWFeeNYJqZdj4+zToVAOo7JjJX+YkSHzhGCr6Nv5wopR
h8PgUd4TbvqyXaxFLqc3zKnjTe3AW0fefev/zV7SRzULWRCwr0mJ07IqmhJHl1DFtF+MqaqTwIqc
HNhNDqfbjNkwVIVoHjxrdqdTlx5aVTY6cKRsUSqXrCPqjD1FvBwcI4NkTxIfJfIvEmHMIHFFqvpu
TflDmYqMW6X5vUdju+hUZ+sGzZooAXuyrFmR5nJRnLpXAEEHxNEKrkmmFM34IpQ0F7aa+fKlr23j
gSQK8ki5oCIBig6CRqCwtyeHGd8/ITKlk0iRRY5u2ozyjFDGCcl6nbaM7zB+E2DGFc4pj5yavftx
WqBGGye39xof7T2qaQuruEQ/EsqByoV206Gjr5vg0gPcMpjo79TkQfN9dm6Ef8Rr13RSW4ESTX+O
4fgC8xNnuGJSd1cwXD71DP01zyuAfuGH72+7Q6oqwDuFCMKokvvpWYycnGWv+AeK0wEXG7Es5b87
aXpkrm23n6LQ/nuz9qsl1dzyGj3mYps/roHRPs9JUBsILzKT099uGBWXSUtayHplM2w0ClCFpiih
lZSBCbJ5MHS7s08Bzzy/6oU0X3hY8wnIfScLgECBhJiuBxNl3VjoUSQit14ipofoW3j7RQSITt+x
7+uF/FX6hCvCG0JCrAup0oKaM0awBV9hTPcQVdq7T+WOk70E54ehuzCSsnCyx4SC5lwVZ/uu86w4
HoMLDmpLctyu+CEyMnYPfQaKog0/ybOyCJilghwxPrDWraE22PuB3dbEIrfpnFhihl9109D17pZp
qRCOdqrQyYol3M15gYUExnLl5+nBS72054bL8t1TG3alW8/MI0iYc9nRS0+zmMSiriM/t66UOdrf
sw0RUlU9pV+tGRrYwmrbxc2OowHZxZsSMw9brNaMkGqY6U+MY4DEXzj94CQEcJ1iqeLOKu+Wc4nf
mabNxJdJaeKKmW4vSAPAAE1Wmd0DlrTN+262wsa883CmsC3p7ggyUZoTNOT7FWwAhCMbhrBIQCva
kHPiGTQUB2N16GGIouXnfsSYdy4iwNCYiViS0U0sVcczPYZBcsym58BJMEpNrqFn5U6hePHNVcZ2
sOXBa4jNn0/oyk94bhA01SEZaf/VRj5ODldBk/lMC/+Kci4EfhyS1SzUAdPLGdFNwWHnyq7zizL/
UGB9kBlKOVM9DkJDWK5FoPuZJ/yGXvToHqUjeu4hYBblYXq8+Ubx2OhgFR4gMTUwNxi0ESyX2b1c
T80zXrokl+8NP/DU07QpH/dRgdUjB1jrgmVz5MS8/x4oam9cEPGyoMv7Iqwn8A48rWkMghzXLCxY
lcvk3p/V01fhO4MV76rNjQmVI/h+QRMlnJz1m3XySpHvOIjGL6VB6+vpmwTzr22UP5D3vACCa7UQ
p2loxmyxYIBtJeW3LarMPd0QgZxDlvFPQEgTpUCq2hUM2pXq8c/VA28obkBdRtV0qmDpFjsZUiHA
tWKFkOPf5RGywh/NKEqZ1W1BNZaNO5KgqgxNo+LLCliCt7Z3NFDPzUHh7vwLXqdsQRrrm+wGy1aR
xcUbjipR9Qjx33YxiSV70hPTflJIettHDj8NnZB+J8PPobF4GGy9V2hzEzvmDH06D1E2Ph9JafyS
cpyo11a8SMofQ+9+AkrTO4RjlE3XF3C6Wt7OC+tOsjYe417ZbXrGPNv5nIgExboqUCbKrRqKb9cx
U3FEnAQ0sg6jsIJY/OuyNuqL3iNDCuolZFZKvkiP9zqrRsigEshxaPtl1eLkR85WQ0FbRg/O22iv
NF/Hk7pnsx5dzKcLGaJ+CAvmJQ+yan6eAOS8xSkWgQqkGhHjsduQjow6dFr6I7ml2KyX+VE2DVAF
qq7dSlpKmxlOJkUgRyGndvM2LoTJk/xT8rS5SxVezLK0sMOCOQMB8+Rhm1TP1ECDmMFHmK6vIg7s
LxGPt7osofEEr33Np1/3U+jkA2/T2z+redlk5vR3gE20PnxyzG/ntGKyrrdngWnFACMVFZtSPTZJ
R2TclUHAn/Xk3cPzy+5uQMiTtp1qt5v6pJ0lAxLu7ZGmFMhLEKVhSxccdNU/ACwLynpLts+8MdsW
m6zZjGxtdRfaLN/6qnyVK2s8qtf4cLbiVQVG5zuN5qpce+C3zQ+WtItsPXahlX7NiUU138Cil1of
D6muHfkYYLB5zvQMGKiw6Jlv0FJ1qU/cOrf9Zit3PyAH801UySSbpz+3ITZmBKQhku9BXeC4zMx3
0FD6l1jaMkmLM7uP1fpJY7WrHbF2IhNPoBp1wUxN9g5B64bqTqWvM2jrEBlExo3CkB8V3oDCjhsH
Ih/f/4ieg4SS+2cbJ0BiNG8CTfZyBa1f2gOTGThqMxxw6sl9VshUwTWEkDkKgdUjwANeZ0ZOE7hL
20eBzWHi5hvTOdiBXnsCMpRkuBJrVQpHPQ+8J49I0Ci1BZoEcPF9qvRdr/N6VAhAvEk+B7KjunKT
TNwc8Ky3QumNEHXS+KyFjL3hKEsFDbAVScd4rOtJoUaKipX/INe9YOcYU3pFqO+P19JsMKW0BKb5
XEeOuWgqVAFHfvJGMcGtNV7mle0b6G5xnEWgnYM/5Tjdy5iYHEvnZjTuYcoDfyhXnLrC5k93Zs25
gECCW7orWuRCuE6H9tGdKydWMowQYay5aOgiA28uGkx3utE9ryrlumZT3L96uhuy3lGmJVPHYcJ9
kHDnj6SHqg6yBNs9vPl7RPOgcMnHcp+SIt1z1tUbr1Zhg71loT+1MzaXZ5V7Rfmjk6uKpTUDSqlY
DGT2sANB94ueZ/tAXCJOI4aPLb8Yozcmo2+x109380X+IpyebRT6G+7GhFWi56ENPjIoLj+cFoG9
Bj1in4hNK1bEW5VExXzYzlILbttwptWvHZz8Z+IK2UmDU6P2lvfIV9BZtRWfGHsUsRggnZ/nf89f
SbZFUdNbRldUytqKCjFmQqYXpDBDrohqy8A7J1BA6tQGdp/zocrwIgTaZrnqhGBCFsls5ymmbWXa
Qp8n7ZEe2kauPZ96jxODn1qpfMqq7/M9OdCwtGsOwTgdHvJmDNEOwlMla0/ZTwO4unJXIgFLsShK
LIlVxGYS42BMQdaaaEz6a5y7ni0PmNSAw7LiY8v6rnmSYGCueBP7ViTgp/WeVIkoLABZnIH1ruUa
tOlp/n+qDSsZdGULkT5tRCw+bN4Dzx2030GNWPnfv5iits5aKZbA4MU5HuJ3IrOV0WziWT5Ju8+n
YrlgyFyNpq6D+fH3hRIp+FZaxAsGx1QwlBBl2dDpHGyMipdTFWjbKHqFZgN7WFVkHOsw9JS1bObg
ASTl7tokm3whMVVylvF/g28FvyEClzq93/eEEUuA8YVwR+4gSUoo20SqHfgLl8PILrzfsjSD/Uet
Q9VtbilW34BnKAMaM3h00B3f6yy5Pr6FCknxUMwhQqIa+ENB6nQ7MAEbXp2M/RneIEJCpYEQmyRr
98MFwRrbttXSb+225Ui2Gn2uUTDvdyxGUtTogbDGsk8fw0k317DXKlJWn/b42tj01+JZqAFur5X4
03rV6EpzKAegyzQjgM5qOcRqA6sO395qFvR8YFOQgCgtXHU9nINaq6hfsQ1irgLAoBCQlBxyXRfW
SbFOm0vAhM488WIr1cKJmd2xzFCBvvfwXE5JsFO+LSb6JPj2c+etoCZIHQo8RzQYBDiyDfn78NhZ
WcKj8mgClWaNXfO29sitwZelB7LD+MVZ87yTS3zm0Ei3YWur5CeXw3UWPYDuFngw/xOLVDbK38Na
+p4pM8R9gLIiZzpSDM/1sqJotSDoAAJLmD2o8R1fXE1UPsbo/4b5vhrIsyondWguIbpvLu78Z2T7
jcU/S9/GyFVJ9Pe+/Ti37Z/9vzuM/9UDZf4Tx0faZBJTMB7A+cwLGXVGoShvQQLGD3yae2jjLp2V
Rwe27FyBHZIpwpQ54zm0PKEivYUga0zsCjh+Vdsd/vlixKMva+uM/Azq7g2YgvZJS+8VqMUX1ICQ
Fde6+7ztIaeVtJRmhzSXTjQXcIhuhbbDkj+/3nYroZu0257ujbD8NboihUHZgMixUbp8D1iqeH9+
gUgrDEM9MvZGV7HwbmNb6RzYpPGT0tin8VnM+8XsQRZP+EdRVae9e2HDnI3BwKb75Es/IMFPRHmy
vxrfFzAikGJr5vlnaq9zz+I7PNFQ22X41JLTcm/URAe98erj7BLEK9asukFNykCvxAWxgECRwMkV
SnB1VG5hfx04XzPI88viiFXqD3I2lB1dlpquj9t1z3pkf4QolCVECus40lkhw79v9RCx0KWi8W1m
XqAlK6LC5xa8N9m5ETsIhhTQWiWbYdvujGLsgoIDZr+Gps0mdYyni1rUWzQA+j7XN6UpFNpJU8wX
VEvkV0oNvRSS0eSLvwgHselbswknXw2AYidh9cx1XvAIug71+/Y9s5HPMIXHKgGm0jnuHUa1yEHC
Ipzpmi9R5pfTsd3ySENCX2Jj42BghcTfZvywseBLdBK1FzP1MW2tRc5NZdfwwBTswnU6FghU0s1a
raDPI7Du/fJ+izNYqwi+dGLEyvTS2RT95rUDvlZSh8Pm7h68dZ4yxfLnYjRsQRCDPILKYSQftLhD
E5eSOhrUHuxldwMIFfJTrot0m7ZuSKfV6LvCfji6XnsGEOzu0QA/btVy/Rtb2oKCt6qrfIOwlDV1
OX83+fHcdVaZOaHqX2ZI15pdd32ifeQgZS6D4Qx6/R9HXHDapRxrNM18fHBfM/8bngi6yk04rTVA
QC1/yzTOiGTyMOjGXBJuZeMmOb8Gjvl4JDmLBO0o8irjUruxeL0P8QMDnGUnRieXdWu21BSd665r
LQYNlqYus6rx4gpmswtwDDZSdibB4Q5LbOq9H1sbYKdbVsL8pDI98DZpLVpBieg+nwoKsq2yi0iA
z5QqCiAuzPjik2yWzMD7Y65Oev329ow28DNN+sDFEiR/iMvQ8KmDwnAJwGyD53jnUmXOdQHG6q3I
Rp2f3Nd7dHOBjpS3ZmFugYryvjuVis7+MEGoWm9lBLuh2z3fKTx56H+d5lXDOSYJDbvZe1RFI+Tg
rxBofR/z8GQQewbw6TPMNIx3pPCUpr0/HAQSfLNfTSmjjsr3Of1UxyD/njYgu4CFBbmmMZM7AnND
RvbgNCKuAI2hNvQfZ+2NkA5drol9wyGoHXKUMW8DzaHxpPDj6XrL883Oi4BFyBd5dZ0wpPUwBgPZ
QKFzda48y5Cb1/YXLY0L4EMJERXxWZW0EkJWdYe0G9n4wAc73uNiuaNgNV+fUwiiyE3mPuX4D6eQ
bzw9NEVNYh5o07rtBajO69+qgdEJJqBaNyRgoRyuUHhiuFlg9M+GSUi0YOAfR+pVIPsLgDsrKTqN
XI/OI2GUu2B35duRNRQ7SqseavtqY1LLny3j+3serthi/vat8jFzKlgrQicI4+dUXlkN2F5K6PFh
zz4cD0KYbhF22Y0YFWhnH2UtKr3U0+ojbZFrSW+Swl5dt5C/BEq5nMruEzT6Pk3z+a3Tkaj+XPx6
keufTE0Dd9mekmSzsEgJ42YFV20UmL709IC594TCc51/fk02IjsbqknWslGsT9uAL2WbiKUOIRJd
OIyVl8sSWoFl5D3GPP4TJSuox6aFHOYWBrrjdwH/fCevmxn778oMFUrGsEily3vecfMn9Yzef6IJ
Wg0D6F2OdXCnnb/qPaG1SiEdv5vpT0XqAVfPqN8n4L47R+saf15vGOq/9iBDG4air4KcZryPsG5m
DPrhczPxoSDqKGDahLGUJa9UM1kefQ0oKCzoRlbj5mLv2KfPJPyEbCgX6B+2T/HvntJL1m+pQAXb
Ctpx+xDqbGoFCxG094PUPZiuR64GXFI/6CmpcPbOdbsQJ+cD7jKlAJFmAgqffxF5yicTGbZtB3lU
BxNBbAs30IOlTYsICmnOn3zHNQc8R1VEV5rw1aBBUWvek9nSZmWrcpLfSf66PJTIw2KQwOxKViR7
1J/kEODIf5zTsmbzu5d6LjBljyTdbvW5Mh1u1zrqHXmIWW+q2wlalUJREYxzWnW42GchUsObKo4S
vpMpWB3fOD16dZn2yBmk4nsfmZ2cQ9BganV+SHa3l/TQEtz7OtWbnDMchvzfxA91W8KiGhlbzvLM
cYaBkFCIRYurp413PDaFGq+Nn+oAfWjobzKsHwtrwdLBZZgf3M+8g3TkqB8sL5pfEaYdcU76adkt
UOUVGK0/uI4dwYjzZfsB1IMc0mn6iZt0f6LFldkGjCSmaEVoS+3o6AjIgZdjDfpfHQ7nYe+uH69O
Y/YkQCV85Sz3cfH6OLP4/IRn7MwwrZoZ8V/NUX0LN0+BnrRxGqeJSTf9ic9nkc0/SY84vwEpsgBV
IkCxWT1JZt+U2XrUPCy4A9yPfe2MU5vvARd1JlPkZfPsmaQspdX05nLLbQn8qRMY7KPPAh33ohCs
bq7W2pnxP9IZoZNDe5MV3Pl0IApj/vbw4x1jtLhj1X1EkrSWSCTu+Mr8vPEDn85C77GolunBDBD+
8Q23I5tKH3M89swPZIgeYjQjGmXGL4i6QOrbD1Wi+Lno+GhxKgOEIoi74wSPI6tt+8kd2u4pNWtY
K0/4KOF5fcwAqrUN8ODsxUoDujP9bg+NJJ6q1dnCFbVJiK0dKObd3qNHeYkJA8Lg7l6b5qv4sg/N
y4RqScPWsdnRuKHoUV6L3Yl5EZCCdpczQuCH4MBuGizTSn0iE+BoZhY1s8rhKYxYbkZYapmAJ1/C
Itae5eUrMEpriRdNFtC+1zKYK1rgG9HyVkMzcpA9BEUPqtnZqPpi7FHyXaLpdV4tYX4K+vfJ0vtg
6pCCFMXCyCocqodjBqHodnlZsv1p9MNIpLKmsPu/Y0fP/+XnfIcEi/oF9UbMLaCQkllfE2CRT2AZ
UtPTFMdNczGcJGFvH2juLEv0+zQYjKoL+jIDDlc3fm5h02fLlEghN+p+qVT537LSJ8qviWfIdeRV
CzA9NeKZx254WAYB7qexsUwcPBhhkz4WzVa+OlJTiT3TY8UBXHxqi5qv2Bj3nlrWxiTnSmH8/p8R
+VK0pmcRnEFThjBCLt4mMCyRE9JiXf/u4Dmf6PsEBAPKFXq3AIdGwh/0AN1D6ZqgJw7h0S9Wb/Gn
z5PbF8dIadrQjDbi6v1glk3JWbx6NMjzm/7Pb9yKfAcoWIt/Tn7sRfqJDwetfiadVn9SQqKC1t9v
NedM47QD1Cg9IPEFJMHwR0pMNHL5c+WrEFZ7CTwGxwInbAoOWTFJSTpIlgQEIsubreoVrl9WjDAB
aGfTlwq7nugjkfDUxorpjuqKLibxGyloNhvQEOVHBA3mJX3SXucUWOUmYaMVQMjHdFjPP53gHoCx
UdLe2EpznqBGuHKu59vjcxqzDYOJsXOV404R2KasKbmjtEd56zGGHINeqnsqLEZ4UX68nt5ecxyD
3quVpVcExXSxmzKYDo849+QMIzAGHMAE4KBaFrpVMiEvxTMsXIgO+Cvrh8Y8Un/ilmjDn2gZCMT2
ArlDtZHu6tCXJsuju/ZCcMkWdVGX5j027YpYHCXyC95mebWSUP4nDsmDHBzUWoAyYgxMpga2xjWP
zmxy1o4A+jkMAaym9gBiXUWtbP089kYbeJWSqt0LXih4aRaEYNRu38fzelCOfRsNBGDcOhftP2X+
wj8En7koL/D2dT+JLYppFRyVWgGG+WhogY7KXUycMPDYrWSLyf3d1/1zP5k7lrvvmTbyaPoE6cYi
CKCQThDoXMmBJyAJhIWfDC5e3tj5pMmYKaJsRxRT+duuTsyX9+q555fW5i70c82fYGU4kOnY9Vho
4jWKDQrzdlMJG1Ung1kdCAokRkC16QSVLsDteXwWEVJpF3cqJDhnFud17/HZX+wM8z6TaoeFj5xt
Zl1cwOXkh4hvOQAb1KMexNX7LLjCqYORxTB0Ml9CcgLbw3d7N0LyJ4+SizC5CiblAm2SEuVZZuxF
AUmQlQVaYM2Ljph1HJqhMAdVKbvFkaPMmogYWBqZcWbk/AJBdXR7nUktKoeXozmgc1QR9xNPF9as
7CWTsNT6e+gnmm7ss3lCCZQRxkgHXD91/IqZJ2zU4MQvE6DdPkuc0W/ZVXejxSEEZlZn8BsPBgzE
dTy8+MpFBOj3uUcFj6i18Y9IR2+O5nR2D4M9hJDEkg0nQID/kIXezzNN+8Xr9l0UBf4IP+11lHB6
J+ERlW9L1FF6edk3vYdMK9hue3nt1PLx+5OoDNi19h2Bg44j82xw4ZV1J7B7Xqus0fzo1qtbcjXF
en0KoBUBF3ParytNFAs7LRxUFVYaezx4CjPakEpOu2kf+BhWuns20Io81jrnuGPglyFxNZDLRaVs
MlFImm3EVgXTVy3GUmgB6FIEl0gTRGQEJLSV1P+Xm1r4zyfS58FHFlSk3GoASl1FVu/GMRuifHoB
oGkGKTBiMKzcNA6xwq745s2rDVnebm2gBW2x7PP7dFwTSDkbQ4FIkuBx5o8pJHNRsFXZapNTTYMh
DC7E0Mcws+tIFGdLo3vP2Y52OlRkw0gfUb4Wcsrl5K+EAagvfDkUK2T904HXLlS7uola4nFTkqpZ
Le5yTUJOhlZy2dyZKguSP3EzWHRizLM2xc/I/kmmoOA2Qs7bya8B2oxwH0N4T2cKY/+wtmmngfeh
hTPf/3LkhXJ+Lzo6C67vRCWcjYcrQhE+udLbkxBEKmu3Cm9qIexT/6JwtAb70kOV4X2o4AQGdIeB
FbFXwFZBv3c/XJ1h/IzQQOUMyfn2qNBlJ62DlFkLs//TUzeEaPdZQZwdXRjNr9B5amdVFhuFfAiu
Cnq5r74iUBAJCFFcFG6UXWLSOyg621/P20mubYCPD9YXI/d3jdjrbS0m9UNec/JR6kibdgwKCJ3m
uAjPGy/QmN8wpRqYAyKjgIKRxwzHL6QWq/mE43K/UQF5UWkBx1hxT19wcYaSbbjiBu9Db4DRzXDw
JbXmvKkQPdonA1yojiyXAuvNyZNbSUKpYWZNyjXM3uifJ4Itl5KAoF97F+5tlqzTiblC8Zl8YvF9
8VgVcOwCGMjtjWW4/emir5A9WT352bSITJLAivIkI0gIYRI53FL2UncWNfFD8Aw/rL4mdjh3BZct
CDUAYZdwEAyWwvlKJ2yO869OrcwYQn4Q6aHBqpJrgpT4iGUYWENzKX+1P9+SdRVZg/FuwU3tPrtv
51HkqPFIT/JIdx7ult4EHMRfDkMG4siYQkhJVij+ed2uEYlkbv7duoe2ZtvbhBc9VADsFwORlBpQ
Y51xZ+xq+9nclVbVZH64ZdvGuW6ClCUa5UWP+RTf1Oe3V5YVV5agC4lcXamDQaG7m50s7oXnCbJv
O5hcnXEd8uyt26RHfsji8U9Vgdja5mB9NjqJhEkQtD9ZLuOniecMKXcym4dRleGbLGw588DLI3eZ
2CpZXujZQdgkN5imft0FidChEhIl0UC5JIlg4m5fl27mKJifGH+3DMwVWmDIaLRdfRwL5JgrTKmp
bc4hxXr22X6nAMzu7cBc/5yJgcggUaWZbb7KDjJTo6xKa9tULbbXHeB/rOXHq+WtSI6KlWjQda07
3/B1FfFSkf2hBBCO/0l4MrpIoqLoyJ0xvPtWD/GSbVzKEb1yoWwlkeFRD2Zs6EIGnNhd1da1jSRM
NeKOdRCZFl9M4ykLIakbslvhV0HMqRk4rebO0m8xyALF5zA2tjg32pu1RdogFfDPkhJX8Rm59Gbd
BpfDNLqodRh+7SmZcMaG0lQawghvsFndJk6ieezROPUffwo4m5tILoc1C8O7D0+C8kEki2fZVxYD
Aeihly0xi0klAR0LvlWad+Sj4yAVapuV9M+xvm0597RqBgiaLlsxHQP3TzSPhblGlACJ3q6E+Z34
MPlpdmBFUoUuB8xO1FFg1O551/FpVs/y24t4kHG0LhcKjZckeWfRuR7Nl7YNjJpXf+Irv+CFoNlO
4ubw4SmRiNgn/0xTZ+WoTutyiV6ByS5GjLnWuZAvYiW/c7tiSr3wl0Wh2Ou/35fRzj/2MCz8x1p6
1//q+JIpDCXlAVi0Owz20ErMk/Ky8mhzo1GJl59kj1k7I1mfN0XH+37XNOPNngsD5XyPgCAWRs6B
7SsZ0bPqtJ+PoUyrdgGHEveyHQ5Mzqm/GnwSQZOfNyBO6g2eG3bwrLBi2ECUbfIlX6121GUrEbH3
5MBeiGuhzYuvIa2pksy78V6gWcMLxMHnvyFkKKdQfJdIOgjcMP5PL0/FfiMpap5rjGEURAYKrdIQ
dRgstNgO83N2vDZLd8ox39dBiWaws1Vl+gXfJCKqqdxc8QXBptK4EsVezPYlXpLWj+e4j5Z4KbJ9
F0wbD8RVnYZx5Js3Te96uQKjQTr+L0hES3sM5spaAkryBCnHeaYpUsctMd1iBft7SxxChmPVJd88
kyh2Tw4cdDnFpoqHgS5sEsE1cBGQ6ea19sCIRYReMx/SvayjGLh3dNHROc8dgQfCHAP87QkQ4E3M
L92ZKvmUMb7/xEZiMA5JGXqI57Pi1zD6Y+cXFr0s+4t0uvsXyNSO8lQVghP8pGJHObhOhv98w9gb
guScLsyz8vOAtFjmqLhBNE/gsPamuXZ+Vv3gNoIVKvsa9j7t2cRCd9V7mHWi8w7KWoIzdZMutH7c
AVcHtq6HQtA4re8MUE3Kv/BPmwpaBFc7iNJsgU2Xl9hqsOB1rKJlJHV9F6H6f9nEfkio+161J6Op
mcik16H937VFDmslJqV8VIHQHl+gv6cVEbTYHS54QewDnqXXAnc6b72Kxyg+TvCT1V15kw45PTza
U9erbYf5p0BkwXuzsXarsrMiwhaVsKoSSNISZJ9T9GZgje/Rubj3RL6pACHmvGNu2c44C7W6hzKf
JRtlFTaFys2itBDJRdv9rZYtlTTiBfFPthRdttOhOyUVGDmC1oGRg+Ynd6ULof3E4vYRTTgTH/SI
tf0Up/JiEHL0+AYFSfe50dyvmr/CY+E5y4JlHPUAxZERI/nXppH8Ko+31vBV7k6pV3E7vVLeo4AZ
lHCLtNzlp+WKm5gwEtpvx9SAbYvxNg2g05D//oCUgHe6gytC0cmUi2KwjIaSFr3TLO6s4w0BAESn
uk/wmCWS68nxRS+vOjkEvp4e+Y7jlYTGU1QbTJOdItU1fqmTk2DLDEsQYcv4MWAopKP5SYNrJHaZ
QumQqeGsWjxcrZylOM5oVKmneYPcFRR5SX/lHvBWcOoDdTg87588taXXAr1cGXchxNBUH+8tCA4J
XhPRHuBkmG8ZMCnT+nHpGj4UDHgSsCD4FYRV70skPEVZylbi9bi+M4CJwedxSONsyx3tnNe2wxz7
Msq/vJXoY+44/r/2Gm8ys0VBUnXXnx35bE9Zo334cdQruqkUvjeZawrYnu70H45aMXJq0MB3dbe6
sxa9I6sbLJ7miXQyAikCPHreSZtbEVRahhJ8RZWf4K3Q2ceubq38jcuwm0TeMvROGw2+pX/ueCFr
DpCNbFttlbQSGrQdLo97GXA+ySodapZy3CWzW6FlMtXfT1Nrak1M6OdIMuzobyTMIYEDG10e4Ijy
egVVKaXB/PmjZQexUjUcJk+leRl5pLdfGYbIfOViYn0uC6oLJVZLox9w+4ZdOhPA+zjwJnd17++5
gyjZ0TY3RQmxdj1QsNmEof4ofCEfsPipVSOvrL97KJLFBrwfFOTNUZz6X+C7q3c84B2PpTz7weT1
xMbwC517xFyl3JDFJw7QQINLyxNzABKEOyJqQIX6UpkWnOu91wEwUVhPMxJPRJVRxcanIk10einv
Aal5JznaVVbtoEJNtAck7oQWMmEemqoLY7woz18y+9SiKFad7kMkS4CH5c0uu7jK0V8rhXLH8c1G
/XYxxPjUiBCaZyQDkR4j/4caE3UYaBnCo0Al4eYyZXWNre3axqOixFQbUtpnNq5bWTHp1dMUSY41
hnKDNCHb4DygdlIJ8c1kYOhOcTrw35ef0+z8gA7rAs2xSzqJPTeHpx7JqK1u8FD4qHSXBEL6VP01
n+grTxt3DQuNpBkkCX15oz+hf+SIM4KivGHRTGpU3MNWcghCUyXZMNaNR2roSqBTXJfE/GAjKcIu
AmqZHCmsCNaA4/ijQi03hJphQXqe6tvnFt3WU3sRmHst1UYY3xge42XvuPJkT5Cztf3vKvjuQxfr
ydUlock5l+50bu6UmyxM+fEsAH8mJKQy0dLP1mXKc6UrxVLmMmj1ImCnXBFK7CfGrBrVoldTv47Z
p5ZUO63zkS1mfZZ8oIMkZpV+oN6iCvhLDRliyiE7Spms8CfoY3YADipuSdtVxbQnb8sEZkej8582
JmhW3qxu9xDPPTVaPL/DqNPsvnwB36kAPRUWOsMHdnlKrNz8jQNoxydsSP7ZyyXn3okLn4loeajD
xOXnEvUxA1cxsDEJdK67AFtbkQxEzhJvAKTVu4eYZAKfi09Oys59+PhGdBxUkgt8qBXAwpUwVPHi
n45sbHw975QFUiu5BcBfPNUyS7k5Z+aQNmYMgV0BArZ/A4JimAhgjt47UWHPgri4ER7dFhti5vfI
+I5UvDULrtQkN8co4TlUWTruLupQ5Yfr3ZTm1EN7o80uRD8iBFL7pPzh1NM6N/nXuegJSVj7YDkM
CmdVkn43OIQX7xJcSkNpVyHEKF39JYoYLbo24FZxxNtW5EoE4oFwu/GU35uGxSavUXfRObXL8hJ5
IJ4hP6mOSi107H1AdIFkOEmmGucVLbUy2njkdpY3Zzt5107DxpTMeSKfMSAzaUFock7oV6HF/BoO
esJHIw4dR9BUSpX29AmOIExS6biaDnslI/Iwpe+ICIUHvnaMAum7wlQpJffHz2Gpe3Jnhpp8J4A+
DAY2poag3uvXZx3duhRkgOZ0F+jflWTttqfbZnMsKuoP8++rMSa3UisEDpx0WOw8x09vfaYRl0L7
vzpyx/PVtSx+OBFlqRlQTB9WNA2WDUzLsV+AU4c58UKAcs7lIpnOyoOHJfg2M5T0fKuog90LrxKD
iHj7ws22WrT6NLsaTaZVQY2XyC9VzKgwn6W0sb2OisOuqxNsr75jEhL48ystJgpdK2WFJQhGayzJ
bnbfgItMl5360Ul/9lAGZJ1CHqstcY48abrYfbsEbNWbMPYhIip/RTEzIJJfJTvRTInnNaVasrdJ
TL1K6FuhfDz1RTpv0LIdGh/oqwg+v7I+fEa+viI4r6ChV/NcipGZsYHAtfdSw62FYJSGWFw62Vql
2O6qy2LjS/YsjvwExeJ69+wMXdV8mGKCI2Z7cBsVwM7kJq1nCGeAfzLGKricR4JBuEzt0Z6bvFo2
RJQtaejGUAGpXcVXSbP+hq7RMuNL5DV5blzUhXfGRDyU/+BuPsCkCGIBMtazpXV9ELgmY5qaKtPc
ZLTKaFZONmlAtcc2ZYy0iLYQ9FDfCfLaSDrichk9oY40KQqgVE3NlqbPuG9ppGqCFApM6iTh2O5/
yz4pPaElWwKREzT+S7Oeflr7yVHgB23blP8FYG/GKKgIDUNsG8hh3XK6Uz6SQUaaCJNSVsHtMd9B
V3LL8x5Z8r6ng8WbCbNYID91SafuxiCWCX/vllo33AyAQ2TIjmcCWGMCysjenx6so6Vfo1M9FO29
GGchD8ylDXdrkZy9EOwDVf26l7nTwLtUUiOebMgo6ij8js7+sk+qc1S4xLmTZxR6UiFJWZkfmYA+
L7OfBdA/uCUcxvF4Wp4EbWA/lrhAQl75h1CJ93cBIIkQeE4teNCsQHfGF5TN+sTIPIkxYc3u+nll
eJ4c6nBuy1Gg18rKqKeR1tNUNKSwGwg+tFnV9Uyo1CYQ9nenrCiDHgStCh5ywK/s+QuLBXGUPHKI
/pdVF8gU2SYH8BvMqWAsLOWi50zyk4Z7rPzGX4FZcXgdkdhQRDxZg+ImDdfNUmUiBgg+Cpg1/OdK
NXFPOUkPFY/gpnyLTVi8Hgfo5c25HxUVVD4TrT8UQajEy+g93AE9X4IDDkgkn3QtWux83CXN3AJW
VEAoSbso9Bk5EX3cwUSnTpvYE6G4hwMb+VaXVIU0GgGLvEb7LVcinMbNF8pV1P0gXzMnBiKgzJqO
oVvGC20dh2EGencW83lNX8xI7fOoiYJLkmwzlVgr8A3zB6gIQOQp6rEBScBm9W2Z4MrOtoFRbW+R
Fe8t9N8s98mVquCAHiKpE75QPWw+r51k2PoXNt8AWWK7xVVAFASy+v5KSTmqpMGrX7w7pWNF50rQ
MPNJuCDuGXTi46R4Phn0MbfxTJih3tT/bdmb4kZq6y4ixP23L56H9LSOYMJIyPPEkwMiw4qc0Yq8
F9KydmIvXGonFipfQFdYJ3Py/QZ6NsnMEAVe9Frjp4rUAkHLSsLvXwP4MBXIMbYZVxwdgs10Yo0g
w+EArNP+oMUY8lfNQGkSipmtthKptu2GWzlFEAjSVYKevwgQxbzNfs2bJ4zoGd/Ueq5iYQxuKNx2
aE7n42d/Rc/6JNpSULjYYls8QdsJHXPpeK9OEaL7pmiBInPOM3VDlFycw30QwU0JTviTOvBsny33
FNreTd6WoUqXtZAkPa+PPjMHzxmFyb3d3PkzOQgP6BtQKg9WDBQ9993Zmke7+FU68cVB+nmDiNvO
vngDK4M4bIDSJ+yR41ukK32LF6NGn6d/Y6vhU0tvkZoGDBdsihXPsGrGKp0J2k8gVbu2n+3LK9ib
yy6xGUlWvf8X9ZGhgk88Sem/EiA+8eExIWHeZjqBEWfit5RQisuIlGApeEO/nBDNTw/4El4I3pz4
O+RwMl6DM3kFCHyZFqu77M6JBaUOo4C2IOr7BaUMqSBsos4Gh+TH6lAiw8pU6KWkE2zT0chCVK9u
7xNydNlqQQubo50gzFj6amf5hL5hj0tHbjTlmKtOjVqF9z7ateKcVsF9sYVMfjzliiD7EDutfmOG
ZVJMIlmdtbzEvcQe/uQI8v7UtfkAegwUPF/bdS9dw+3SobCJDQoYr47ap5UJHPmeAmS/uyrJbEJk
Q3HEkMfSb3aSZyOFLPawBdsx7ulmmZ9XPZHJbmHxz8tcwDmHak/Z5v/DJeZyV4jumrrx2Zs27YAx
MaNMi00DK9+XjrSFKro/kVqMzZTIb3pk21AAvcM6VwQjk9OG78WH7qqh84wY9zZZpJ7phO+2KKBx
4RX1McoVmXzDuu7CM+lg8JQWLOZvkMNDAnClNeub+Ifq2b/FeNrvI+wzA/axAlTOei/0cIGrUHo5
OhHG4ue0cozgXrmAVMexJ+k2bcVZejbHMq3uyPHthNos+KZBKH8zT9PD0AZ2keWSCCFPfe2q1sdi
IhSfDLRFA2FvX/biFDsN9BG0gg9VKnvLJS+Wr88tQgMTyyfva+TZfAWiKhsg+oSCCmK0oeaCQYqP
5/q5ZO1y6YL1Qx/Y7VyTWbZkvWHvQYF8rCN/P+RPnp1lhd59IZXsLaVWkeRhbewXSck1zL05y+pc
eqGNZG5ypNYvxClTMTKLVLdwtDrPtMHUIS1qDjsh38Q1lyvEK3O7DC8LquvAiaCkFzm3V+bF/vuj
1cCmjRGU5/n3CYrDcmMZudXTNb6cIz39SxTJtgSqkHsOsWnluUlyjWnzaR7SNMqt1Q7Ell6SADZ3
W9uDg5tNxkwtGBQRONsRO53HKNsAxUPuS5vbDsdj8hoCtKCN6usKsG5BQLyR5hTrCsa/hWqbcrEC
tvtiwvaL+qbFCAsECndDFrY2/SRDsH6gyDgivPhLatKDgvK1nBaHQtq3GTHtHHvnmdGidBKYs1EN
/3U0vPuDWBKuFq6affnHrTxIq+MLf4vHzE/qN86oc530WuTc2cOAp8uNopvL83dVnhd/Y5FN8PCS
jQpmTGy2V9zRJI0X+8mbwgSRo2S9AwHsQijO2UIFbd6uWcmGVaUD90/160sPKplKNpT4v3vI96Ua
YOjICrSxOE8qOiOqV6JDP9Bkfcg/ulRRsF9Fsu5lq9NbTwlCH4GDKgO4KYG3bD+ySrOf7U35EsGd
nnOaWBtNgVNK5ArSWQNsiFGV7DnIZ+yvZwg16RBHbR6huNqjvRbZ1chLfba9fvIl7h+CHR2FwSSc
IR5ZhuU7X0skOgCjzp+6VWjbSP3ltf3QKx+pxQInuAmFQrwiBk6zxdNr6zCbsLY3Ub8HfongxH+1
8S/AgkOIlRlTwVBxCoMhCleG5xKpxt8hTfZjjKjakTjh4gQg3A/M6ApFAqPreVxUknFP7qOkYfbd
G6mIXad1YjWh/DotI0vq2Z02QEWI3Pcncal5zxjnrJG7pw44HqkmWPEZRMO+mSz4mj0nrixksWPw
bAx+MTKhtBQ2Cx5qDXyXaXIvWX1f+ki7HJa3SKWpenWHigbN0lPCTHx1pyDmwx9Yx9W8mpiZ0QYW
A4rHlvuX52NGsV+wGu+0to3pYihbkgYRVU5sdsIQqSCoRoKD+xzBicxOk5yvRDR+e/jFh430W8cU
d7VJ63t2LdwibDGXUCm1A8wag89EnYW4E3NvMNXlIp/tnwWy+LcM3Xi6U1rfWDiC2z+fzHGdOC33
yTyNMdlJ7GN3d9MVOJQGOwsj8h8fNZM/7zAzVGwoOUsFdcTSK085xv/uiKbu4V8s+t9Cqnmdn7Ew
6KaK+D/D1o+qo6pHPAJU5JPxCMd3vfYU9HJ7mk41625KTK8Vh+2nnMrbMN/5Dz7T6Ds5Th34Ztw8
LwREiTCgMn3Qu723bZLmurQkhPwnXvnAriu886MJch40UF1FJocF+S/5jSnKRDE9QOlmATqHqLVM
F9B5j39UTJUjMbVv44qa5xHBSV/IvswCWyRPrE+x6MWysNTX4Ob/FVlVs+bYsLRReNBdDvRNj/wq
rA2hiqNxVrJ/TtNswQJYgMi/YPeFFcIjGn7PsJrfM2Z06eRKFLGmy26cBZV9+gVOTj/LB7P++fzr
rH1Z3ijg1H6pWhyg2C4W8khtkKfu9pHP6a0jbf5OrlrHqoIhbXr1WuRo5QPUh9lG1wX/VzLvjqLr
4us55Zk/MSxchLLTTI5GkkpwCc0J5ucBeqbznCoSiJ60d+h1BV59Kw9RYdd65JzhTqIrHqgIVy42
aBNHtGyP6tFiwxClM6EB56iAK4zp7pjliJC7Hkimno20HR5RzIASxsQvXcDkw/o008a6EogIxPga
A4Aleawbk/yWRFbcIB7K6OC+drLKUPDzRcPmzsZGU3UUdQEb+6/ei5rswYAA07uKKbLXPX4ZhZZz
Pp4epw1nwYpVStUdeE/qrwO5ZDWzxl0G21I3+iHerp3uZClTWC1dvoCgXAOs+eLARz+xfniwUArt
8y7ucVOtnIDuz3qhPbkouhlAltJeMdrGNR9vR4HBKBeir0DcIP3btUugv9/AkVYTjMVEprentWbj
3qSF/zJ8N/oqA3DrNMj66B9o8AI8/aBys1/wBu3NB6jws47cAe4vsa0wfdi/po2EUfGAPId/sr9D
6GyDctUu8FB/VEkdWNYXTxO5kH+bL5vGBaJu0seUVYwk7EUya6ZOBDlX/GxxXVc3K1aCY6z0Aahw
9O4sYrjvx2ESQxjYIk5ITtF+VYrsttiNvEgjPTdRtGl0YLYUp8miEtQV/RRVdsnWVeGCYy0QUMZW
QXVj5OyvA10cgF3ZzyOvVXP6aKOpIPLFpXxpMSkBAOXj5zT45F4FvNcfsGmotBn6RQ5hQ1mRnOm4
JOQkMCJtN2/WwjF07AdHJBkHpK9owb6IgRBRWiIHZcrxFECAV2Wz4zK40t4CIbQ4DmhY1sdPKkc1
36H60+i2GOl9PUEZtxJS5t091eFVmyHAFpgn9hiY9BpPy8gqOCpzY1WAT8GFsN20NZHSJyoXx9wE
vlVJhG01AvbYGEEovWzK78YIFKaI4yLrLi7Qsi9jBtzLgJYWrkPyAOIixKRMIidgrqmlwdvseS4w
2IgjrdBa+rtA9JipTotvTYTHys3fUlb/zk0T29Lx+Y3u2IO3FNK1j5Tw+1WbJcnls+I6ICi/2niO
8ae24PDjxCegIuYqx1SKlBowsqpLeCLMPSjjU5CdAdNIfXQQz7y9jykUlX5gg529078viQBx2OWi
FihWR6slY4ubiG8lIWL0PPhjtWCoWnPRMe5IUUvuN8+ARMcbB5onnfRUloG+OP0JdY5PAZg8Xl3K
t0j80k75NbmgkfnCxDIRaRvEF6j20xKycGG02iMQHi13OmsCT5Obl/9rdzwPMAlMRsmeBoEQu24t
9yrWbleiYFfq7UBWe2GjowanUNVka6aLiOIFwzADr+ESS4Gkbaqtk5zc94AYFTDye46qH43RJahS
92SxKF9j8bnktqw3egtiKw1kS+74aUcw0yoDUG7wha9p7ZxpqBTPjS+dGOIjX9pI5qriYSftB3ZS
KTcc58oOc8QbQse6p0uEXQVP91Z8sv+ftKBRi4gxKS68G3CwIiGdCUUGo4bBZK/kKd40on4LLnOY
Kn/0jphbHdcJYqilVpm4UzbCoS1nzhCeV2pNxBnKsadWjxvXolQuSRzzJ5dACJqBJLjJSBN6LBKQ
msmkIM4Ke9o5Muy68JarYqp/1CJ3qUfUjpvdagFoRAuX4P+ApassoVBrPhbepY0sXJ+Z31bbM+GH
7FUWrjzAP4KMApB/1ZdIEwaw5/0H2D1t/9KPMFrnJBS5opw6PvBuIHacfYgqcVSSDAUXJON/HG4f
X24VbKwBvAvYULiaX9/fawZQdinpWxl96w0JdqOrTvo6WjlmielrsxA8zu31oRUbdiX9wk8ORiMS
CQ2q1uUWOeYWWOe/akAvaanReLTyj9PG+p6xsBfRUUdqFOYfSAHgio1AQSEXYrEqND4gNTrcE1bh
aN9cwSDzvO5NLABh9czDyRyehsKVxCRF6kn/1PJc/f2bjfEsxaPW9JjWf5xGKoTJ52yYHve9Yw7Y
5g5Ykx9LAkW9F+HwSRFRGAtXgMalrup4zhkBwpb9DKDyNpAY2uk+N5O1Dw3MgzN1VjIV00NZv6um
bOqXY6Nhzd/uYWXr8Nn3xuk3M0oVwYuddqFMYmsQ4CdFS3gRM0Yeo3ENWxZrWFLVXeBGZfOi78YR
GKYbNxFuIlzUQkY8j3qT+X6UiV85WU78PIp4rYQ/64aiDUWV3e1AJ+LIFDs3aRjVNv64Bt0HUXZ6
8RUqnq9G6w/gNtDZ3O9dDmS+BRgQQjd+OzUZP9AucEXWWQG+5kP3hFGssIzE1muq7W9QObcm8iQt
RVKFRhtX1nBqI0aqvx2YzRHRsy47ccSM+4KB+crldqwidh6+iReaWBBTHYKeyelVLGwfMctZXP/H
rrT+zqk8kNexQqA7B7bihH3RipBjlJLSXQBVCxmvbm7phVG6OB31MlQ1r6GoAi2cThs8tnVv4dVN
CfOa7UvmGrv9SzQo6T5VRQ6WDR29gDW1FqdRcjq0gevYeBfJmb4D1+xStSIdo4WYtIiUxH3pnu+1
+hA/pEM5aRscnkOTOt84UM5kmSp4ZhBu0hnpBUoWRdtV6de9NJs19bi9o4f7mWTGgjlSDRPSUWQ4
TNF9PH2IP7vPZf4bFvRB/RiJd1TZl7ijX4zx1ZDLpouN4DZNkmOVFq1HA0Sqop9V9WAvfVi1POoj
pju0yFVicrVrbho58d7A7Qk6X7sZ17P1yRTjhDql/4Vj7Txytqlx47YZnhPzF2d8egXwZxxIaUqq
7x/chB85V/vZ+zJGi2/sV662zhWDMCKbIdEa6Vb+NR40L8KZcFCLOVzpzgv6UXyVexSkxBO1db3J
D9qIpledYcT11lk0eFVbTnkXV4xPNtnGN20KzHVQnO/Um6o2bVZ9+BqNdgvsNDIKdsJsBi9cylJH
T097UI5MeUeBiJs1ntI1xAB/wkKtHdd/JC/TkpgaK/Q8tmIu85Qw7bG5QeK2Pb+zD373pd7rpcqr
dxdEcdYHuR8ovCEnY0pu7tRRlw5GLtIeB7t83v0XoVLF3IwgRncYwccD9+LSkr+W+N/V8DZMBfbJ
SVKX360Ihgi3DRAp4rnH1YDUL0SOlo8aOw56bxOjVvg5UJfkvPzywpI6oXPyzgzTo6H7E93vtXsA
1B3u9rQUkJdJqJxEKgrOSk2ImtGX+RJfUYoROoCG8oj8obOVzRt7LG4J631fQ/7qoH/GknsrVEC8
8WEcoZyxBFwOq+42oBFxMMUgBjdLJN+r/L99CYHrUo2QNIpodlo0dBUl+k5ohrGoLj0BObE16gaM
SdFzV5ErjyVmJE3H4zmwn2djVjN3LiEDmDvv1qHgv22mp6GfUwANrpOn7s3lUEt00pOIfF7YOgpl
PTyMGpnvuiBF1b4qJMaIF0TtiLJqQ8VVsdIN3M+ebz0Z86BBkFYnJd93oGjvLEZGS5ZOpndmRg1i
bTqgmrxxB7WsyK8PF/QU/8mIVIO3gz7bCTeGdNxF/20/4BtbBSROtbvmPb6fMieak01GJonxXG9u
WEFI81BsBxKKUpIsrScaPAWQstBKQu3k6ZafdC8Zm7u41JcnMXo0TBMNORsl9RkEubu/glUbKiAo
IseY0vROjEPfTif5Rf8GYRDJOvqdE+y8F0M5lGuY7rOAdxjWgaKrzjco1MCpYKtq8n59H9RwlxTh
6OLE7MCI7FnWs1iIkyDXohwyCSkSoZ48DsEaUApaUWIcgMbD1n3AhV0Mjx0ZPW4e5N8rFgHCEmux
pkogsh/zdddQTDxaD2YTHzqpzHNhTSAHX+xNwDhyMhE8MTD0Jl3T4bzxYEcVyCApIUUStaUEz+tm
k9MmqsNodZ9rLYMolchAFDtpUP0+FTtYwrw84ttvK5h9SS4xyZoLsgduSnyeP0FQfe4pQ3tvxnGe
VhnEPl0MUaekxSBPlkrhy3loeL1q9pmm8k7aa1zlzaleB08HJCD/xb2jJA9ovHtD51YpcUV0hZY/
HX44UeB36V4R1ZxYfVGGbpZWVhgIm3K579HOEMorfMxa11CX9hPa88guABBF3fSTXDplg4vgrULU
T51vboUp+3BstnK8MF4at+exqxDgRg9a2Slfa1PE7wcUwHIEvHP/OH3Yz96uvQbyaI3tp/h7KkX8
cMB1v41GMyYdwOeyp30rSRU/2F7VFqSo0hLWVtpE9T47tb+r1Sv2/86sbX5Tp8Bu0C0ISqOqhHDI
N6Q8paCxSwz0RaEys8g5uh46IclsR6xMW5ALIXpoLRY5tSrqZ4nGdl+2FOs+HJTEKmQeEBYN0nUw
EbCovNwL5fw/kiTSZr0nH3HSL0DzDYEPDS4tx/P/idfFDkH2/Bd7qI1nBKBq5FbpilNDEMohExbo
Ug2Ts68wi2mZeQryok1Vb7QI2QLUZ+CH4+06bVyCyMS8OevvEHQxffiYKvswBPc9oXbZzq9IF6ZM
G5qvLVx3VGOorSxthXPwPKg44BFjkfgvitnmeHW5FoOwOgbPkoy7b7SYW506atMVutirpI7WPZVf
Lk20B5quCFuEhaPAqOQzN75HRw2ypoUzrvvMU+Axow9HTx+ZVVTGBPv0KIS7IkRHa5mCGQBDmWMK
3JpXCpS9ydMjIEm73YcM131ZZ6Hx84GsGDzx7PFYE8+bID0mbg6NHwceh3OhkyH5TMKFdmEWPkTk
cTAdnEKhUwWsHUaWF0BQhJOi5Df8TyziqlooIZsBEIuUWKtMIgmqGVQJRBRGBZah9qhvcuEmZ2fz
vHlas2xtgcRkF4Pi0D++RxEaLZVZuRiHjO09QrAWeTatUXlBRTFihSUaGzXX+smfDWewirZozz7n
5SIgHEliIEgE4OdxcL6uwiIA9FMSKeEoaIU/8A5lN3/HuMUsYhnG/FnaXjBp6iS5dlOr0ZTj5mUd
rh0/FI0hoqZKBvIEo4FQUwLEmTGcPGtJpJITcfke24jTO0xlvJl7ubu/v9sCzIp8B4pL7SUJ0HhR
cfJy1wrbwNqrunmwP9xjhyizwC4eNe5ZcImJIuY53yOFyPaEIQJQtoHpndm2n/gpiTObFBO2Cwot
+irya6aESP6LyyRiNmOv0PTs3tfrUgSpdhq9v/XoeMrsvXRda29j7LEbeIPAKwIUUhay5CePPyw/
ASpFtEnW9BGqsr2kgB8Ly0a2NREOxhejVRYFht7wXfgI+eQ3gSK/nsZXkpDgnRR/vrY3iaaGojAq
RUdMQnfvs821S3UtbMpADs+UL+rWQJFwX1c0FenDeYtWmdQbdl019a1BpXIk6oELqMDRuin9oYPr
uJylsNDcXjSVOXcE45NosWjycZdqGK8cDSAyPDu3GFis/pYmSv/HN3EWzSqK00E7h1pjUK1AsoJC
6QvO8Mi0R9inIueeqRd1irTxYI+yXdol4K4JiWGFrOOc2e+M4+DyPxHdonU+fN3S7GU/1ADi6Lc4
EA2Sc4qtWsDaCjXIc0N9/bGMaqa4c1B18hAHwuye2y6E65esQAstfWwRt2RutACAZ9QtLu7b13OK
f0EACcLs+MPd0ieniNkHLketcOgDkQDkVBiK8FkPyxKu8+uxVhfNufkT/s6hKWLePjMI1quVw0tJ
kg3rSdD1ZWk//rUnnIxAUCfDNddOey5hNa6L+iwJk/+CDflRP5k2i13rjeUzsjxpXPARJBdTQ4rM
7C4pwv3WiCDrEsJTxyTmWS3qdjO9VMnzYvvVP1otbMwUX9D1poQl2uhH9/G4vZxGWe/eOQn7xpqy
gcC5RpeNkw0TCS7zZVbWV6G0kYzwrpfEgPYIs4kE48LgISTOMi/Pf18UG72Bt45sQ7tWurDikvvW
zGR3CEE0UNkgQX+nfMpXYIXYko6cJ9wFSotETPSVAQQJ9zBxgdPKM7I9NIJ7jMcJBHAiwWLIMpiP
Tg+WwlKuuoGbJ7U11XNjDNK20D63CAUJNu4EtaPtjgJjTgxlrc3BG3ea7yR8mzclI0kMgZquuAbu
PQJsy/pwVsGdl6YUuVMkSUmF9M3wCSqzZwAleSTS+iUWuxTSUiUOBEtXV7QllvEfK5zkspe++7UP
U5EXpPmPkuM8K+rMokQUoFE5rKtbyZ7pSfArjcopNrh9cEDiIaSsLAuZSj7I+HakmBZrVsFUD0n+
xRFTx7XeExoNQ/+LOelpNipeNhMjrnbvCHDPPGZ5WjHXBGUlxcVCh0jUyVsIRJNBBSO+qyIJZ379
39cC0mjQqy9A19/v/NWRUl41yzQfm/BTItzDk6cnuTANbqMOU5n1tiercnoOAl/19z9MYoqUUXNZ
6hARb3R7JH8/keJpyJ+p1g5rjrUBhWA0BWFOIOTQkx4pysIqogwVGMJ2aalD5crk7aEi95CPKgwt
D+/DpWl7nh2EiL+5gaLzMm/1neuj8kWfupslIFa673JTiV4Bx8CBSEmm1K0rKbwDmsp/8DqIBWku
39yWBa6CINBloixoTFL4jJiV/tc/y18ifUHOZ+ev+84Du3D4cn9+jcVFJ1FkyLWBme6B5KBlycxu
74s5zutwgZrihI2kzK4Q4U8nA1KcNymIMDn+0ZYqMrD67fDCGiDr0nIiRvsC/CxlxSydDxYeAaSV
ncK520//wbMFLSnoX0RNzBC8T/+VvNMYf8O3tipL43BRQEKrWb+w0ikM71QZOjvu6PwPHI/z+XUz
0JTWUf1lqahQdVRqwMF79C5KABnC7FOlWZjtp1vSSIduvmQNv8lyDVRTykQW2qAhmAZMYvMzoMg5
PaLi9h2oCc16sKg288+oPwxQ5OaG2WowZHmntO8abZGqqPGjPNA30JOg3/vTZtse3GhJIMNwPHyF
U7JL8baT94vh8672sL+Uz/4g9SI3PF+ush8VIiOpD8lEyFHsn2XDS3wdei1aWl53V+nN0ERCctPl
WhT/H26udgjhBBoJ0aCXP0NSVnKMfZ2E+xe5me6tn5GlnWqldZ6OJIBm7pJlfnAR262gQpHyvs8Y
ixhxxZvV9QhjJ4BtpyzzmPyZFoCI++zWN4A7iVlFhHVvQC+xQXRF0T6Tqo0+MUd4+6JYiBqht33h
YqLXv/jYXGbcJ8pL7UsEWkA+RE3jAXjiLdRXZoZATN8zRp0J/tJ6K9IYhc6HzOnFYXSeEBj9PKJ2
uJnvz4ac0qcS5bqGT2CRWYzl6iaUUW5QUogfQDMVXekXrXlJVty5KyDVPMovXLt1KQnfS+vhb5UC
T4K0npVjtWbxsJuUHht24c7GhOMlzRIYrtNfM0s3k+xxi7gb4bLzWm1NIqr3KW0QmyvbwF5tCh5x
4vIQC7lrbrhX0e+TwbC34hiOeIDUDpJryObILt7FSK1f9Q0HBGhUI8GHreeKz6b0WBBoxIRZuqtb
8jXIouahshPv/9xlbdWofUHoxMgc8sWFW9M9wdh5PlHe+QQpKivo51CtRmxXI/jeKxESPjeMQlsi
CCG2QpeUdS7SKpcqb+WQ0tJU4SwTntV7wUDIsKbxO16fPePVjMbr4yoTc6pNk3KQwQNbUxdDDcLU
s2hyzJdJs0BPEAgTf9cuqpcDMDFu5J0JSC47tkjs9ZjSZlyESD86poVP4x0cv9Fwnbgzxx2GKvf1
QLXA88L5Uc/cAkGMm7iGgr3JHkukRk6vwjNJCKAeqFdfrauu0891bXMRFT8HrRBL8TBdn/7sfMqa
6SHjJFxSTLaEdjZ2VNOgpOLtGogdxGi3Hn4rWM7m2yIHalMyTXLX9564utMHBMWFacXglQVqJeGN
qS5+jMXAzdU/3SpcDQFlw4SBOHh9gYmt2pKR+vYjaQRxCbl4dVFkwVRAZImSPoiUGTUT5H9geuhV
hpEz7Jv2U+K8GqRTVIdr/qxJ7L267JHdBw5mDxTZnRd5uP72TCW8a6vEqtFRL8MAwB5KUbSZqsn2
+QYFvGGMcKWkr6XY0DBCzzdoH8h5fSwSGB1X2IA9u73ZRMyIPHKNhZSrNmzwqgS6dL25gXNXBmbG
SqAtumgywpCERtwqNxNl0jzbpJMLBnnBZMlZnkTP5lxU6EVixMqDDMiEg5c++/X4T3kNyogLGjQS
ji98ofQksoX24SeG3PLdSXib+UJYOSwn1HJgD9QdIN3xUT4bJkYa3qCDEhfAQwLu/y0BFxMSn/uS
tw2zx6EOV6R8DQRPMQU/OU4bQKeCZ+xgapDKsNQK0sJ0GBRbeK+ID3jVTSuhk/vKwaHABcSDQBZU
d5YzgsiUHrRadIvZQq6+Mc7zIFMajD2jxBCIE53o1C3zifJNd5tYbdHjErC6D+Zj8Uh2n4vAcF5a
3jiyA3/+wQC3/+aDRd22V7Qu4ovDCALrE/+yJFx8lHde6sRt6pw7ksA4W8AikAVRzSxVyLvNjpla
OeyzXdnoCBSim1f6h+zVE35gAKuZEF0HCGcSmygw+VCgfj4teqtlSnxNKXZ1UNrFIFS2wPB9HSyv
pC+IBzuZP28AvIX5yjm8qgNymtOk7CltcwXuRXugT3K2KJmCuBqAj11gZ93NASZihN7I+NZ4FLTv
xIJKmsXJ9SRnW9RESUn4J4wvC/R1UbxB6el2WgfavXogu3NHSZ1AYMCKz6ua+Q3pt/b+tn1E9ANJ
nAM5G4XZcsPW4L8USb4NQkOyPg161cMgjsy8fGgACykd4nF7yIFSEyO/bF3R2PMVmAAMJHRqGsWI
PhrZnwKa5f9hHy8CDxZDTqp73ZMCbLnWBEemDUQgVEK+MWkNz2s2bq2qxy4DJWjaa7BzYvdz1By/
NENETwSYpY34ZBb5GSKMo9bmA8HIMY8EUPoKWPiweLnTBk4kpNQm95+AwLBbP6UatZG5g7irGBvt
8QSJbvhotqootqK+CiVTxksAQAMgGbL183wHsz7wTlmFlOpjo9wRUooYVlJl7WgH9+9COuECxVv0
3D73knFuNPjEoUBH4Q4op4wi+93wMcWmS2vCxxFSs8rVvtX6x6h/ijn81xSHwt8s2J+5kNvaHVJH
hqfZfMxhcQaAXsvyPa1UkGXhJfhJASPzIwHONAY091JZoIPDhjTeefZSSsHjv2Qwx1DCfpfsI9Fo
tio661qjMSDpQHFKOtvG8S2J041VPUdvsc7zzIA/Dc7JsiGJ8ZGi0mt2PrWbuooxKtWa0Rfkd+k/
/7oQ8eB+B0KnpAl9luaJ4iX9C2eaplNPOiIiPhIA27duTAwgLz8xwovk84/4MG1a+MB9tH51PADl
hP+WSCFKNfnUmJTgRmdjdjJnMl3B5M+LHiqTMbK4Z+hDRuWmJB+VYiQeqJo2ozkEQKfJoEtnleR1
Be1D4re5TE7Hv5M1LAaEPFVMJkbIfSceBaGiuMYm92xvWZXCPfVU45EWsTfwpuT8tNtn/YzRaAdi
Iw8Am86uZ+aAYZmod/9MD/IZbdpAXZCg41VE7miRloL6wiKBoQcV282tBsd8lCAwaGMMFWYAH0f1
z0vOg8Oh78dRXXPIrdMoDzZm0aSPmaUO7I0YbgrYNq21q+cUiXOgR4/Rgu8YtYhN6ZdTQ1y61B1E
JCm+hg3uOooTnMuQ/TASSigWKzn1wxGgLB7YsMrO/w3FYItYTkaLYxB9I7rbp+rajpS9TzndLfpH
Abdv7403Ad+2flrVpPmVrVsWDpIUTxc9QoqUwviVwnRYJHuJejqqiCHjXi9vSCh9i8iHpTPaefP2
1nS6mcSFOYy7qQuJrAcmD/DbTiuKAbw72ttOb1EkLwvQOOUxCpK7ozQlSZaUf6FSsNmF2S9RkAVe
ujzMRmC65cWvEM5Yi6FETAzUpUmF29/rrbHsS3PJkW00k6nU06utvbfSDNRQUCKYh9+CZaRo1ZjW
QY9ejRHO8fYExWQbT+Ct/GLTsn/A6G+aQml7kqN58PLXW/QABejudh9sGKjMUR/lv/Y84mO6vy2e
wUJb/wp6WNvQEJWL0a1MkxO3BwtDkoAyT2DWtARfBOmgdOl0C0cl0eOF2MXsZj3pcuhLCiDbe1Mx
ivtTGiIShXtkk6ahg0winScRWFGu9JAIXnsn/WwMnJW4NLsYvcebzLXnbfXWAOmKUXqw15EZLFc0
Z86Ttukf5SbKFyqLOlnWAdQuvqohRCl9Ah3p6UmRDBdaRjdlpl/G6JieDmUlD/IJ3tvdoC8F9XEY
1d5J9i2CLEUVWaeXFZJO52lwYAiF5ct7xMXc9zaioAXUVqAO6Zm6eTKw1jcP/IYzaWrzYfqYkLw3
WlMQxzPi0uzaz/0j12A57bYPi6L8Md5dJOv3qkgvW4ttZBeM57/MsetBfxNkUtlLyeUGpGrtkvNX
ZoPbEV9TtSCPOF6Qge5jhwvzFhkYsMPh4u4H2xeS+alh2woh05f5tz3HMTCWRHIp6crd1BKQK8Jl
eZlVMIKSpBQLLFnbNtdEMJIXU/vwLRLnhKrNx7Z0ybh0OvOY14pAqSVPbw8qsriEYmR/84qMzYpc
MDamsj52NkcCktBHAwZw0Q7bmBetr7oV0ai5PxJPMSV09LzcehI9A7WHuAC8ZFpLPSHNxBKK6KsM
Nt2X399iFp4TalXsNWeLHevi995ZEdNRNDSnVS8KspkJFAp9OMv7kDL3Cl91FsWcbg6cljrHy428
+yBBat1oPxHZSpIsCIuswMDiiw27yzkyL+pmYmUu/62XBfRK4MQEMEC1EmO31hMUoShhr8POVAPj
DIJUTdXauOEuuw3giZYBRifroDXYWDqboWXOxvOImG+r5xwEO/mbb8OHYqWEnL9A2W7sERkjVnpk
6RRlO4MfsiZ6yFkY1lE2r391rVX+oGhJsPcykbddBk2ftCT4spVgHcfrsCZJvliNgvim0oRvgNgg
+yEHc5aIItFODdm91MrRKWkuSjy00Woyy9bYjLQQTylSmxjtknCnGyCIQaJ2IZ01h0c6J5L/sjlv
IywwljOoj4+BiYgLIsNqkaakAzSsHe4jS0F+piXZJ0XXQDoWNzyihUE0oOSLaIB+cjHhMu4rdcXx
hJuHTYZ8YUYpCHIcSRsT6BfxXTrKY3kBnKs4g7hBFfAORjtLpNE11DClPZgb3NAjq0p1rQ5UFuJH
8e+3rGjoPrsZmZB94NNOcXiUUR9uIYpb3JQ/+M9HSbfmTWZ5QEyYb/b4axT+3IYU1lc3d7kNRmKu
RMnTwDYLmO9jpswNutQicaMnfq5PEZKddZxK82nncfviJH2VQJpFxF2W7N4BEdzWzDAShPclybMf
2AVdBEg8RI5t+/tfRXhjmi3U6X73h4ltZDHhNmBkX3433GLr0p48VkhMy+1zFGArDk3CVjt4ZtxZ
ruh/MyFE4cg+2TDC67NUG8M8rgaKNm6AN8IZHZV6c4pYu+zoQ/rjUY0p0llwRFK1n/iLS2RwxNKc
rISyREyA087bi3r4sNKjDo/x93/0a9YxEExHxTVedPR0VvySNC9R6dIW5L7/UWk+kzMm2a/hY2JM
PELfGLPraJDgvS7Nw2oHnGTyG8WWkoHqEXD2Q4PpeL116lQ50XDTtNFKxegGbKa+KU67xouWv5OE
swfymVqpXOtoogHjzVtA9MSBvkgfMAESI2hv6J2VP3HHmWr7o/BHC8VznkC9A2D9DGBMtmbQfww5
9LMcyey/UXb2hGDDppk7nJkxgKvwgFDXfNUfwVeY8nZR35TeI5da//AKVAjPCqXcOm6ZETfJggBE
kv5rat1a4pLBh56omo5LU894TkF0udh0bDGtXFx+NAmILEdaiZJ0Y0ZJoZLkCHbeKxbi0ofX9VZT
/5JLH6e6XgTjyyJFjV8bdtK3ZFgXaHJR/4RTw3n6kjlHabTLx3FtGlB3iy52P+c3jCNP9lZWNxCq
d2mHN4YOtv1EOpY5bIZvvASBbyVChXIJ0eBKATyBu/QcuhaJBmCX4f4WJDqcJ7xYi7sju1Jp7Wep
9NVRbaU9SHgRCi2BrucqZSqc5XLEC7y7SfeHnDZuY7Vv910SBGx8efIYU+vXEtH4Ss32fdJe04zl
X4BUhlMLTbyWHqDc6Y/I+YoCASpPxWU3b1tkMYS/2G+h4ghNOdHLEztjagmX0Xw9Iaj6qSpMWGy/
q0nCRAcXW+U5Hvxfa9PFKMk/lijdm0HbtoY4h6L8S6bLw9SXqvaKmhz6jgilzfl+pIlsPmI/xN89
wHyFt3y6hQsJNjORZBwxYyK+vhkKIS/oeJXcRsuxSfact9M7QlJJYn8UocLZ9PMdOlOrgpsy06Uv
LMjJ3Bmy24xeZENI2NZyl/xMKlwAf6xMC3TphTasHdpNwaWU8EHGnPfP4vZfEo5oAEgly5naS7Zf
miw4eaEBqWs/nTxCJPVTa+gytvROcYZpUzwCJ39c+R8k2YQBkXlaaKuGIEdF7a0QCz0s85M1p84A
heqZ3X+kGSRtL5RhDkTE4LhrNxJOWaj4cUZhpOTgCj1lDySDnaVcfDk2NdOIaGfG73/SoGMci8xo
9ta+mGmNe5KfNSGxi/H/1iYjvJQneqgbvmd4d+P45aZZd1BCGw2jOYxXtpP3/n9KPeyFt9YFWRk4
CL5bOieihazTkQZDw3mnn6oZP2Dgd+K5xEIJUFFZgUnAnJuhyvGz5+QOM6WTXUNjxaWU+cWNMVtt
OKCjgYjKfdKh6SmoFf9UuVDHOEvA6L/fhWVcBDn8f3JtT1zSu9ApF2YcgRollFDZZTxDqNdRprpf
U08HgsojfSe2yscEg3j30n611ZkD0kIVwzd/zBOdf2YyQJdfxp1ZgvmMV8DMP4xODKuvDmduYSez
RQAa3Qfoe/hYWIzJDd0pt6usaQ31CQbfDz8lw1ujf7Dp0DulduoqnNyuldPmQ+sQw/KQAC214lhw
wt5Io6BxuQK9neu4Y94qz0AHaQmDz/Sz/IXyk9Ja+q7TbG9/YrcQlOxZbUeBf2sF3amwRfWR3ZFT
AQN2GT+oP2xG/Y8NDtl05kjwq+v0HWo/EIhYSVU9h1XXjEzqw8l1VMKLAG9pWpJupOHRtt+tTvUg
AyhD6s3HV8oF85JC1/m0PnWaBxgjYv7TqRR79vY7pAoEeXcetANiRjPR03lDiAVlB0OAm1BC2HiM
mwrf6HfRd17yvGBAdjEwDOGUyMyCyyiNtUfogoihmzGQhq9kcQ58x5OOuDGeBnfXMAPfwwiTzL4z
G58EHUxgOQzP1xv4q8uffnw9IJmQGdAiXhLtTfNHtCdCTAfjnW0u8emcLzLZhggdMiyvBiy8i/+r
FPUwGLZ9w5gSHS7RafCMDeF6u0YARw05J1s3e23ronv0uwpnI5SYXAPz6trSjlYj/hzqMDn218VM
KIXle4LGiYaX5z5v42IBFPhcpH1XRHCi421ESLBaxydv4GVKungX2EjEbx2owkah7ncNEuaAX/EA
aZdTVNGo9hDnRXTdcT88zN/yfVL03ifzjdXtjiybsyVzYio9CrjznXflOHlSzqCO6LoMlneTijPb
8HTETnlVSeJYer81MjkxkSb3I2eBwB36b/m7HmFHp4Iu2YMMOCmPK4kQcuBkrBBbNv3tyE6juTpq
l157NDcRP4oazFwXbFbluZmS07kDaQOjJ3mEhwsQ5u8/rlaa30zFDbSheBY6Py2J+icz97S80OBF
JRUO+v9gjbz3jByZib+YBiYhDziMgWAheFtIe0bQYA8toCz8rSM8k+P7Z7qjyWCKVif7yrta0UXE
77ex5PXBl6ijNewuhrGoqeUQL5llDcWdEpHopAjOuYSHSjlFcnkXPwS2sI6JjS8H/AEGpz3FRTYB
yNwPKC2xSUl+MSSnAZ878sBYxOEdVPY/7VcmnRH8xmAx0xYfudQtr6TLA91QmdQVHIX/HZ8VY5HC
c5b5ImpcdW0/FaL7SwOmwy3pOWIDtBxE63yX/DDF6uS6lRD5dm0YYoXPPVi9wwkEm9grz33CTjcP
JumlpWp19FKkuJX1cO3OvYg24ZP0SyMTaP5Fx+mRukNdF25GGQYnHhJ3fZuSmiU8iCvoGhCiwADh
TWkNGi4+yntwE6y37YOgcC1v6epm3kCB7+y1qqFDTgvPcoWIZgBVH8B5OzOCkFGtpOztf4pVe8Im
YaRjcRsRaTj/LUAVLzRKSGZsE7sIxmu1HGhXIPpBmBFVJwTgo5HVIDOz0T4Cd4LZSa9tw/TsP//Z
7vAgr2qbVeTQSmVFfqse+bBDAw0+Yl7T5JROjEsoMm1GChO1OQs/F6PRsF/CKTqBDbgfKY9FwvEC
oEu4H1s/MSr4ThC6fhRdH0Gs/8Ba8CzTt2VHJx5tVOnXw4QVM4DoTGqPharadoQmn0LGYi4Q8QQp
2UubcZPDJFrMm7w2Lu8oo8Uvu6hHxzoijk1v1BS+OfIk5h2lXLPiXh0lEbXMwZKxU7kHJYCnitng
/2jk7sFPrzEcabDwTilTclik9QoaLKKB3BN+/klxMEFkHl9KS+8v3xRzwd6v88OuIUzdRDQvkpii
fezSz+w9Ukmdvv8CLK88zRmahZoex0hyS6AkmjlJQi7FtS+kyHcdvseD3o0+GO+T3VnrwLcGchDr
G5xv3hcKFgKRMvGNUazdg5jn6c00iw00RaX0x3nOCSsVSLHv24e3iEJQNohCzk32KB4ZxGBL87Wq
uzj2+gsUPeIf4Eer4dPjcYiCL8twBO/eHAH1dHf1JJR3lJvSLnOLVBPkpvBflZp/C3dJdxcb0261
XUV2eGNKw7LMfnWMcVjM8fZtTTBfc1l5VQXWynbz9HsWD93wJHXGvcLPcuJGpHX3YNXkL++Yd/uF
TUro2QtbLPIPdgN8dgFDynIwNvnTht0eGzqDbUeDNj1CqY/Ti+Dfs2nIyxz91KJKgv4Oa0Rvngu1
c8d7gqaIXbx+H3y4RPbhJ7jGo+QjDktN2j4C+gpiizH7nq3CBOP7vq4P6hv4NegIIJsF+nxY+JSb
R5MLhqdmGrKa79r0ZF8iEm7a5krhfyF2dguhDuGYyCIgSS2hFEOocUnhVPfwTnZl/7stqfzSM6VH
YpkvkTcYWhTSM8DvWaYCPMqH2ebNi1ZXkUgZehzqpfyy98KCochqjgNDbmxkElKySXX6x87wcovz
sJgon7PYOcQP8VK7M4RzM6MA/EFSIdvn+nPdqiqPFB2VIOo3xESlXR9PAy3D3qeeNsnFPJ4hmzwb
MnG54DaalziUMp0qtR6vY8ZIbXzWFz7rmutPhzD+pKmgwocKyQhNksnpIJ1QjKvNP3o2p53wF5qc
/NYIHK5dMoTJbzS2LyG/ulYFYqw85URjkOR0faKgVOLAEFFY5Vs4CqJ5U6BayRZzPQCQZuR5q4/N
WphCyk8jBQwvYBHlTYqLlM0eMC/IjrVcOF1zCVfYgmF6xKgyaUyJVFMKbkCfjj41CDKdNYk4JN1S
tlb4t/juHf61J9YmCDfZcPAKhsjfi19+w4eMBCh3puxAhSlVY1LJ50i277NGy0b1VHdLTBIXkloJ
x1UFVUllnnC1s1W++8yKyuuHWO/UOZHin1B2N3/DgLt2O3GbTf18Wz13iNNgzi1UZwglS3zsmpI5
K824GscShIxWY6L5BKfcZTwcXu0kqMxu/kIA/lqA+VUxyP73v8hS8XSkaFwARcNvwMvwNX7l80ZH
nbkqU4f/7L/hHn9bxhvn6I+7sA2fRKFgCIzlgzgXrR3XshOj/0ksty0aPoTP9/VUKBthlsFNmeGs
grMf457kA0+xOAP2bb55wZ5JNRtmy/e0/AZMJRCtkxZnrYcbQxrTZ80xqQAexTqhBDc7BgTkL2YC
okA9ji9AQEeR93EWioUwgRybE300inVZoeWJ8MjkS56o7iW6D+Bd9FBR7acj3Kyq2YT17sKLAxlo
+DLa19lNN2mvan1eFOz7HC2k8FUVnMHzveTh/jzVKyRkr0eto5cweQrz/Ic2Pczi7OrYNPbpt05z
p//cAWWylhqYdj2EdJgXoW0EENawRrkH7pv1txsjnhKMzDmlDtHpyDe5sVswntSrpBKjNye3XlDG
H1uzfSsD58gVyKnslqhP9w9W7MGIHibK/NARdBVcnR6oWfGUJNg+YCd1BpcqgTnWc6XRMSNljV1k
Bsb/5uK4nR7mH+nKNxlBvQyDV2UL/iDwZZBCyAgYODO1q1p4Mya/ClCfo+yxMyyekNl0q9HdG4Xf
486gzAAsqrCoDtylnaIxoNqzj3zFI1NR4TKIkmKEzuxkHmpo/FdAj2QGm/QVjgksOzZyFBEfpNRz
72jpR8KRcV8gv9zo0rs/cN7vhrlpMS8DdEPkdM4rhYGsEBYXdo4luuAxp0F5EREsOYbodBrVpL58
Yxu3FLnSfHrJKuNTw54ANJ1u3vwNePDEc/sN95+i/oqWFTkeGmiKIpHUChFl6G2+ptM2XxIOWGO1
Fz+1t8zPD3FglyDMF2y8MPAK+UoR0h0WrQzD4Sv4nUkPGPaKXJkqttwrhnZo8VUV1szqYcQy+bUi
3c1+1aVOeJVaB/JS7uLrNP+Imk+Z0h3SfOsQMUHwB58JvPdmvIW+7EyBU1t0F9sr+8ctavp4rLdN
ey6KEaO/qDxQWjw4VLvr22gqFLqa3f8Lwy/t/V35mRUIFX2aeOhvX6axcHo/msr8G7V0ypZQVyg9
m1ZMqTo6n4XjLH1N262fYndYynlV/cxnd7Tyc8muNK7wIGEHXZd1rwvuCrhaGIvPjJ4vAGXg34X+
r4hV+B7SV92sK32Zo2m6T8IoXzW3+vOV0lt1wiSEOuk5pJ5vMnJq6yc+AYoDMdiO2I1XD9UC6B8n
VsPS02uJqMS6xxpVx4MucxxopSwdMieHdnqgodGRdsloJVlMRO1TuI4RCQW5JEaZrglYDnBjb08s
UTbXMAgT3cDDT79qfs5MOC07qWNAimNUTwxE2WPg+YyvZpf12aP7DtzgErklJAvwd6lhJFz2/2n/
Ds+T5OoRz8ju6c9R2U2VOoWWhzBHOGjihzUhfMzYELN+EntJv7RLR4nnEdw1611WROcqc2P0Mrg7
6EF9ABQrk0cBDvtcVXMW2Slm3dPVXIXmiwFP6SAaNEqBnaayYqO0wSO2IVTxAIKvnNYIPE9ES4XV
Wwx/a5IRXyALeQ0MxIaVF5lwuxQfrTPZo/UHo1St99mY511w/dhE5GsIBFL65hR/RrofuoNEtei4
XcsAKtDb2Ta/8stW0xyVuddw/Ju02aFWDU6KRFRDxz1Zt6ywsNkPiSN4XTC5fVx1ImE1H0JJVAKV
/oyaB3IyyenYfrXXCLbfZi5/l63R/lU8VfKrfn9Ejpjd0r4PSWkMrZmrRDZujfxRfsFsakcTNvxk
rmDWqVBWch+U5f8X0MHz+sHVlLvC56bS+jDTkesM3f1TDYhNdYMTIvqgXT7CmfkOSG2ZylnS3I3k
GMl9QFCvoBr8lODb2PmDmS4huZ5YBfhTBDCSL8XpugJITzDFSP+rZYdd9KmjJws87FhINc9Ph7Wp
WqzHv+2BNDP7jDMKdzXV/nr0BERDh9GWQl+q8KLdR5eEC+d4XPsPWXAQigoI82RDgxsOYB3aXpLd
1pJ8MPaaZ43NqJdmtPi/6cTVYf/4oVYqTVdkquMFJiYGNfxAYtMKXZpEB1aFxHjMeL/6W74LRuIn
tUdcXDmmyheKPP8iOHPP2nelrE9h9HDJyK/SX2QLvgfM9vlh3pdPEWQzk/W2vFgAh7qVQltpuBwg
qnL29QWPNLblBDq6GqhCN9r5he2lKgJORC2a45KFnolDug/Sdsv8BRhnugxpAe2O1CzEffA3QycH
lLyxZ4qOyZp0yU9MhnfeGPlZr39ivtukckdh6H7dcrL0hjjxjWBmdLg/aXo1PE+GvqHjtTb1fH8n
za31alACV/G+bQ/gr/fd8zTzf2R6FhaVJqKQD9DghdgFh0d+ZmnQl7ApCNuhivQpzUU5WFhFrdgS
aB+Q4xd+1wdw4I8d3Dh+EVlVnHflOrMXCzHUE6WLXMUJufs7uX5C3q/5pMF4bUA8i5013lZWbuoR
R8qOzciB2PfVEVC6Zg8/12vlsBaL10y3vL4qmGwyIZF76A0wiLvpgmYqEKiau4ZR2Bohcoa8Y2FX
vnnt9dAGumH1fPDduuBvk4bKYhzaqRe4gGLFHZp4Yq+0LiSAJP9UWq4+jTpCZSjRnzqq0Qi36+CN
CbCoJhVEXi772lhn8w9bLLTNfWkbyx+3bIjIpM46EepPs0Vy6ZyHAQ5OOLSHjFCcpSCNZ4jjnNtN
kJL2JyQmZeWEUDHG3y/4Zesyn+YwBDVHEuDgWPqQDj5refaWOhJF/G9oZZ8NH5BYog3eWhAi2Z/8
mFtmoTa0eZfl3Csy3kkr9sNHtgcL2G7DgoIZe0qNFK6TqkTjN11ZabHq71bQhGzIIuE/fBt8bBE+
STYnDY5u1hRJnS2D2kugSpfbUvCRvNitz7+mVmg1PL/i0jCCGB3X5UdRzrFucx+5hatK4Wl8iCZm
FiCBWJhwreKmlEa4C+Y71TwAGLj5wx/Qpp0Rv0/smAzjgoVHR7TKiK/9DjbftqXfaLNtuD03RK9D
MBr00GXjjnQHvXJdqRJryIcmJcLF/IfaoVI4kUMOy/QZocC9uiGedvuqtAzCyo0T1a9sS8px5FgR
guyF9LJ+QxNnKLHBYY3v4dqqG2wdO8BygxeINgxK37GV7nYqXMpUnwzZC2gcsua+aJ7YZncpRokf
qhSJQAHKeffrGxfor25+Eb8pBStJoebJg4pLdssyD6HHdzFmM4OFBsrEHNdSMcLtPyN72p20kyFN
fIhlfyOyClz6IsHH8ruXvzN3tAjNKYwYSqJ2Bc0uoWGQWLAyJC6sOPxY477x6kCoUKQozmUg98fB
TCAP0movuW585w83fZKo9sU6qmyafGgAZDEfLB1rFXE3z4av/oHG9uEUVB0URpJpxy+1xA30yQZW
pFWjoel9JxF5sovC0F7+iH1NPXrxW+GmYNCd1m242ppi3xHexJacUkr751C8M21881+9ZYM9+FSn
DC0zBROTpjEW0reolMMNZdOZsuFjICHYh0tHIvrz0B02QgO8AKT45ApXgDppgikJYV9/YeDqed0N
kaDwWji7LD0F2X7Hh2QFyJ4eZHmF7PNsCO+iisKzrsAMNEqqVNuz62QiiSRrQpO3YqYOLTljgth0
1GoZkX76z4T7Y2x6cLMyATDmfk1FgO1LiPn0FPgk9uI1lpjkSWRU6dO+tGT/YGKCrH+n3g6xlq98
wlwHg8q7MqEA2jZN96CiaX+sf+yI27+hBukSmhMYsoPQThD37o8zUc1/JKJnY7NEyyF52ywK2IPH
cUStK+V3y++Atn/UvXRWZsFLlgNsJHe/u9DgOnF4dgQaU4R7oB7Aq21rW3XkxjB57e14jgy5ej1o
d+/DrHcPo6fue60cvz/OodlMmEJ5IiwmtlcLH8Au4vZnAGidzasgu3ZQgiDQLp6nxNUEC0kdd5Gk
u8r78ARMaXNxCWR/0xiLMl4Gmn3Zxor5dYdc74Q8FNIgj68WraGLEMAgru4/9b9wr1gc8A/SVDgU
RKT9RzbX0L1/sx1flADmG1a5hcsliRfz7G4BOjkY8ZG2UUwvm9AtSS+a6geVIy3/1iuWjYXUSz8Z
1h+c9N7lmuwk7XkR5j0FvuRIQpG3sq2pabU65iKLMhoafeOylomWv+5CT7Rbau41h3MJ9NobeIvf
NJbU3XvOouotW6nHdaU5XX5+90q8s/uXOAvwh/Udlgl1YPRRIl7U4S28RnyT3MqeLlff7jIwrATt
7ZVUc35wtWwxCb48L/F5DkX7S81KooTbpPw/AkWwozcot6Ps3b66r9ni9HMwP3DK4lFlOJCYBQez
eB2FtzX+dwvGP8NJQ1ceqO3h78mCsli66mgQN9Mfli2weZEWXzeMXawNmFSJAIERwu9fH+/QmUsj
KG9JeG1CMOcfdEk3Jx8CqHTn84c3R/jh7EdaY40qigEFgd7sjKVA4J9aRuE8g2KNCmrFQ3GPfX27
8AKEkN039ZQCFIdZjbaXvTzs6NtFHHbXjEMCyFw8NKb20lyTQIUpVPvd3MVZc2sWmD76ROeasaj2
dffD1qbJGZ21sQfCplsoGhxphCS+kEH0gR5kwAlZoUBoelTTFLetUHoDDparmuMKbl6PIGPhIbW9
gTuIkDrH8tkbYGNEZCuxT0mUhXYcpRhH3znDTY7ajIRkjRrrle3M/xsL0bYPv7T8+1qfr87pEj4P
mmU1hGRYwfNHF+v8XzZ6RVAaJwfDVC2LAqRw/4r8/PitIZB6qHgi3c2FBFEUjpK0HtRkSO5m1sZC
XFczeRtlx0dRdHdhtEyDvucTKzXXq5jDURlfZ12cMLEsBlLvkg/wPv+3GmblF5X/ifWgBlwmVhtA
itJxu6ju6VbI8VWAiQvlxWIha9L2UZM6fj/FuZZMWJ4OQY8g5pp/8+/Okpe0BaNq289mueOStFHs
MgfVtlTn8gt23JPc+8joStMhD0kEgyw3j6C6j63K6oPmx4l3eZ7DyEGvexqI70fDbHJr6NV8r7qw
cViVEfiqpXKdL1+013/gp0fpAaRKpd8gpuzBVDN9qZOmfdnnrucjzcoX6kGIc8/G33wY9YAxR8Hm
9p0ddVqTRE8YMYRshyjJMVq9S8Ya8wsAXOiXPlTKQ/PlZNiBvaWE+CPjdLuulSEB/NTi9T30IvMq
dT3SwIE2wTRahScC2uwSA2XfzJbXDlY988/6KqnoKvlDhc738obyHUC7dC9TYck+XBEvOXGdF5KJ
fxgUxUKDMYjXuGg7CZjkdVzUOg5B41HTbpYu2eaMGpDidweNHP2Y4IygyMSrcwx9xkAgCx9UemMp
kNFJgzP07mhd0VqxKHYmc6yYPXosUlsBjVqOtgwHmgMHphYS5THjF7EJjou0qJuOjawkjGLhYKtP
3rKvjarZ+/7lOt113KAg40wsBzD4qgqhpfbCbBEu0CMILkkeW0i8diyOowEdRN6vhideR0l+7oe3
ckoQkwb75sOArwwlKskPfTrfW4H4xe3euJe7ZK0vKcxRi2c0jo0+8ymNtOBapnFDwIWCmXz5b5XK
aOxjuqtBaRlP+W0GEZpgEI63id8VxvvzxKkdsqrUdqScJRidmtJdJjCIguvH9fpaEXjxesl3iO+F
l0pJ/fx8XnvWUlf2/mABRZgC/679qbRskPOYwd6gtSvkS3QzNk0PaRhHdMSbgYuyKyrldWfWiDCV
rPu5t/NU6h8YwkxpD3+6kgFcvxMdeCH6iersIPqSRCrLUdCgcJ20KriUgkcaYH8eSquiT/D12h5i
Eeo2CyFoaHG8PREzqeF0B6eLspqNGvxXbHZshHZbz/X5pDc9I9W/yz5K2Lj2fJkRm/VgtBB9dBeN
w91ixAA42orTY3tPt7XkA8C8z6blB7ToeAl5sN+MQs+icYYrzuFkg4qNK96LQZPqmaa4cRz2pA8j
rhXu+18M0rbvd79KRntf1plKpLzkYPtlh/ujqYWKG761ZOZPHw/51qA+kAKm0WlJh7DMPx65iX0o
j/HDbR/h7MVCOjlOzL1ACfB5W8NgUP2USIu3f5cQr7sg1w90TCORe5d7RAdf3GlvIQCVYqOWw+e8
zFDllgyFNgpcQjkDqta9XTu5/RhuKRunPUYyAvSCK/DtXrRmdzRjZJ7gJwqmmLBXwLx0fQjY3Zud
n1sj+lHGRh83L1zTF8R9exg/H6rCq4j6vuGPK0TUgpVTI9UcAqqmpDg9oHOxQv89uQThmt311+3o
lKUOGCJZO0B4lWH26NdOsXPoFi6ldpMeUZBBBYvHtWEGBBFA3ChlrxD04zTrspotUfiNyMosy+Tu
Ilx2LosL8wH9FNIfNuHgYKeYlc8wqUBSzSXv43H1ekqn1+U3Ktk0TVDVMv5eG366ozmOB99vooRw
wHRvlx/Zzg9j8HEYtIBzyCIxIiE9MlmXqUApdtzbZ0M7rkpWPf8OLSMmeJGcO9hzHH/ZV1Lk0/7R
PYJtuI14kXbjfhuwC2WgxcifNkoxnJP6BJfpDtZ8W/NLXOyWpXnPb/oPBqchlK6B3T7kcoNOdiPS
1BdjDZw8W/iWzZ0j6k4csidvah13qaVUyTNb2yg874DzD1t/VvV8FH7yzSXzj+kXZzvPMofJEPeV
7uHtppnMIXYENwzS8q4+ddgvXYjEXt7nE/K9Z7BFnKZCDlKuoLYMFW1tCzeVRUXcSYljAtKVW8Ir
ddxcubumN1bngQ8gBnyUHGNEZuvQJE5ZQ5C9ELJdZYSTb/fVcdYipcSMQHJXbvYwQ1uEi1CQ5RGY
tReRQLMQ+LNqm3+/KarSkoIMqsuJwDS6oV9pfeqxlFOGCAzE7U7o/reJxuWMx8WPYpqIlEOwAXAI
muobLh6g1oTKNjOWM+vz8DQ4EsAtOX0vlryLeLMghEmGl/Nkbt6X2Z/CDBIY3ztBiwWX7hAeStE+
RuC11yhjTIr/R9jTf+kkhoUXFfZqISeCqEU7OlZgEoLL5V1oK/DcPO9uDehlYGfMmk9f3xjthtWd
8eNXN8N9v/HyuIsm3YiOMp0eM6+o/5OS8bs2McCuRNfteiTFByMIigykBOi49Q88FZpbHONaa4Nl
65t6XrfYH9fPgtmi/nyt/ZNL0nYzJ2YqkXRNY76y/aYyB3tGFX4gl0Ra4H0GakbXnpdy4S5RBvQf
Dh7k70KQ6a6GWP+ZMzytC5EdCjCABcpyjwCBse2KxmDcS9t1rxEinR+7ziwJcU6GoMX0YQAg3QYS
twKSeGqzlPjpy8sdjOsc5jNo21Q46p8Ygms/K0ASHUWoip/JbEPDAUhYqhJjJdKMgzs4+X0tuFRH
G15eUdn1eS+sJ7RFhWxvbbP3G1dDp8svnoBtoQyS9hSsZSRkN+bjHuy8GZHbjFJ0B3V6j1UAc9rQ
5JceHyNaJpKp3k9S+xyLi2qWBaT85Regu1bYf7Kw31Ji50nYILY6fFRUR8+94k97cEV7q4CpXmCf
vihUDi7NhABuse54iOLwZ7ApBcnv9ZFLj32V3PV4C6RrBTKCZJmr0IP5Cq5mqOOSOLozcd702LOA
8geXuvVQJlyLmslQU+h+o7xujjbXCjs8LijItEnhmVQYJanrDMtPngnxwFfx7a+dCW3lX9KRDoca
ifABSnyAZa1PCnlNJZkiGNK6Vfo1NDrnmf6E8WqWvFoRnwHPB5rvFvuuBQsZ/KObj2buJT8d5jiZ
WsmTjV07qKBkD6dELJ82jnpp+NQYXZ2A5oCIrvIM9OD/K2jwMojZzUBfRnXRh478yNDNM7s/KeHM
I+zdy3jsy5mpJ76nUVHH/MemGJ2S3WTUlrL+mmvZe++Y7bz15Jkx47gi3e/0xnHQbuX6dcf7MrmE
9Dw6XchhXFRPaAspPbT4CGITk/f1YJDO2FwG766flea13sW7w8z1wjFOYQCQ6K3H98rvKOg37/OW
vyk2o5/DDLNlvZGXYrL42yS9BfbIUknbBMEg8VgPr9gOaEZMAaILi+MQ88sa2vHWVXf1qPzTVVHs
2cficdMKncTQAx0rOATeXfDXxWlVg4eXMwb9uvNbK55+xUn3yo4pSbpFlrrKivnVFiHLdZix2jzp
dV7VgYZpMoxrycTY/q8Hja63bb8klig23lhITljaxg/zQNOq4bEKOlZJAs5k6Ynnc+YeiMYzwabu
bvIZKKI28rIyX7XfIcdsC5wDsxeJgj48twBvVrAYGr11/x3BKSa8zH7MNS5XsS/zW0UmLbDDpSwg
55Msfpp0JyYa8enM/hlGMBvhf4ma/6TfipOWDFKZK7bPp+ZCdHpBK6IiB76EyzvmoQLTehnYfswb
2PJ074B2pYoymVCkYeA68JQNwA9W97NpAIYaV6hosN7kJtdnqo3NuOPaPbiH1P6tFIKJKEWL14cz
8k6iUxj79PDDXnTarR4YyuEakIgw0gmPQwkHM6n0e4/EPDqKvpDo6UHZbxUf2b/6NGOSSCY9+Jji
EhC67OEEpw2raj2efixKoUEvLg3skHJ+5TzJUPYI9k4BBncXjGzfIREJ1Xa4SL6av9WBfiwR/DLE
n5HM54XEciJRUheRxQq0ejCD8OkRTEpFt2j3rSLi36z+1PeEn8nJrsB7rCkc2wmtbGgPe03r9hXe
HKjwTElFRMjN2xmR9b5gXoMIOFXwT112B+PBs3lkLYPBEKt6vr85P+x0Xvl3AwvyPfsD4TV2e6M/
SEo2L5oLgcKJInS21WrRe3hhyHNjzh3ym6Qmnj6Pk3BtN9GD6TdTOrQlmeMNp69lRTc6yghx/WUu
p9DGNs19wXqFhBuZAqFz4N7ud74MFE9Y7hXBB9PrkD2lSqsGqOMO2TXG5rJ7Ai146sqWjQ4yyhvA
iIcVRtN/50ryKl1bs82aBm9SF6INOfVE1uCRXIpNvxY9LXBvBLIE3T+WKezjYNFskU0ztIksuzJu
+G0u5k+b6wvblLHdAw0R84lRmXGpG+RRpiWqOYkx6Jvv/0jXrlg9b/irQm4YUFJP3Y1XxXE/VbC0
ZMuNu3Xut6CtfIUaLQq3t10D+lrfOcgJ4yOp8zIm+QeCYKwmFwFh05Bc4yXWEcLi3b23DYb0SO1H
luQF1GmvhzoiFg5FYv0CQO8gYQZsdPUqr1Kquj4eSF4ndw5Xou24MUzd6RFNtzcnlSrHmxxo/vvK
37ojNpc5E1PEmTwULXKkoen0fm4k/sYB1Jo4jslab3FX+t+0IiPHll56MXYZfB1oCzE0uAjSdd7g
mgVnaXK97wufgVZSyfA4y83iwEFy8IAe5DsjpFP6VBMtn/kChUkkvWyHh9koADQ8QgxaFTmGjNi7
KovTBrHnRfTlmsEO8Y1hF4qPOTQ+KO+nNA5LqiJZW9oR9jAszAdFTcHrDAHrMXtd1WxzhTHNngaZ
GnhUvV8syaWPNEHsK0kOCYxhet1Ee0LEFcqyv3RZ6v6S0e9Yf0OalshzgaYELT6WpxCOlUUTYS1/
CAV5sHXZWkcBL7P6sb9xQOZaySJiybFSRWg1kWCP+IHc+1g9BegtQTfeitQfh+TpZ7Rna1x50sg8
rDtDBFgnPeBsmHgpcrSwJUlrNJjNm7POL5BKtL4CMn9Tff3XcxY//JyFEj48+a3O+muImLrg3AaH
e+a2VziKQlKvcY9RHO3ZjDOK3uGz44hB6z31sCSaP475PNLaKBQbUHWBnplfA0Hladmx2Y543hyL
/XAlG2ipnE5GN2X/+LfR8nl6TwjrswbLdL8XHXXtfRH6dA3CN3OMAKGJqf7tDBNJVXRicuVQDnWu
n/vocYl/h7NwsPhnPLcqxaKF+5sukYYTQAoIyklnQ01D4NhAZ/M58bi9G4AYxKwFXwV5iGA7g5aR
Iqq2QyDd4g3ctz+ZYk3kRehjlF4/PQRHOkBLnoSwS7XWRkk6ordMaQhznQxkyHgUGtSa83YREuIo
QY6UqSM+5LFF346C25zQbNbwECMpkwBJuTkrDWxT6ng0eO9YX1P0w+O/8Z/1ndfDJyq4HSTySnW7
JFjfE3jrPi8pxz90Ks4jo09/J6SabYa8xJ6995BKDg0PYMPrw4a3uuSea3Bu2GWOfZ2lhb3sJHEQ
3kGQz4CV14IU0UtbLgGy4t4hNRoH1QUyELEj3qL4+X5BVLo46qYJXKwKM1tpev03Bek4ZV7h/frW
pwfcgSUjrH23g6X1S3n86+S2e1+siarwyrH8TGcXzD/jsmGTO4WWB484lm++FYvDXnKNk9eGGto+
BfbrqIim32iocYkXBG9R0TQZGf9MQ5GLhb5h48vfYPs9lP8QLeazAZdO9vD/Rn51SR0bbQ4Y9I0m
DBhj6dfBA+clpbomwR66RPCt2Y4E2R/4dJVioDNO0ukFwzmZl4gbFgG6BkDw2+XislUmTAa8+Lyc
qOFiXZ6jM6waGWQcL5I5zlraisiolPf3K77Qe6YLQWTlQjvwS446DUzh8LV2+uHhjnWfRZ1p7qZD
QB3UJxs6gZaSZgLSvKRR2kBA8S3OMSKq1OkA3oaoU5FcWPJVe6iAnQf0eMmQ7cDOq0KtzwLsbBUM
MLup5tNqD5hi1Lp6D34fZOpn/zm+8PwZ7y1P41Pl3ywXLg+IO/cjuSlP6JDUzMPZCbiAxegAF/vm
iWO1GX1Wz4nd/WwP2curv2MyYOjg0N0W7qQTeTFeNqCoyx5YUzC2I3NIfvVs6ZnDk5X6cCL1cwI2
Fmr5+LnrMPSaZY0OVLW1JhBULLxaiFE7JX1SSSOg8wTJCraayVKVfMNvq2mCgc6TnLb/fxX8reoH
F7h/T7xLSNMrPnlEJ9LG7dsoZdxtBzYRDYyLsX2hC6UP9ToizVr6aBSccf8Cwef2tnh2LBdQ+nJ4
UWapXlcpe0v0A0LWa6PSkzc8mo8rCBMtM771lCD8ZHDSm6Y0RUVw+emsGrG3CHPaRNZSs/m3OtsY
0JAqBqFNcbY6k8OgnepqVn38oBkQNPx+0YC5ew1VeCVssydlgDzRppThJMRhHGFO9ITseZraoxM2
C3nn4Ecli/xPzumjGpx1gLKxfuKAs22q0DmufIi8PjJKouJ+U1HdNsON8HlbsMbUaHl6LnFM3xWq
2DsVe1LZiaK1VBR85Qa56xI8i7uRxzc44xrRb19RdV/+FdloiU7yw62Q/z/fymhSN9fFztXsVzS1
gJjO3seD1ZJCXg6SDD0V+lyx4LEa2hLIRO67JAEIbkecIVc8ShdABZG2pM+ohoJKuzN7Hp41YRnW
bVkcdtM5eCLCsqqjrWJVcxYCRMXYVyZUyNJ5oR0a6MY4qBxSwwQJpK77l247qV/HU/TMOtdxHwq0
00DalCQ67+Gs++B0LuQ+Nnm4DAnLEcXbXZJSQhIbv5lxaf5j9tIhGZdXa6liD4dKDaDKWAv2H7I+
7qZQvJM97CAYC0eUCgCu8dVnDCyAlRXcvukPME7ifS4WReoNnUAD9MS6FS2VFTow3dYBFKXb9/Dy
wG7YG5zPKSAVP2FYtG+lzxxNTQLpwcU5SSWYKwagMsnlfn28pmqF2kgat69JBkd0SSDoQi1wTM2v
zZquyYMfNOZ9FzZKcfai6mAQ/8LFhz4IV5gT+cVkhkyq3/GwOLv7xcTtLY108ZaENTsDe89mvdoo
V3r55mMQy/vvVA+UiVBZgOC/hdNaxNynpqCBb/1G1TWMxemA/iA7FPOZZ40aEFiWyroDY5YlgtNw
/DwANbubUZsl6yxB0MdNFmqd75Iuz8zZVIM8qUoIvdlqgEFbXWZZc47aypcwXsWOMwCWrC7LAR/f
7NMpJv4Q5oZBAPgLQ20yF1szQalSl1Ma/noDiI49wSF47sdlAk6A3M1VyfbBfIphT275i2ChvBj1
rx6Yobyrak1DzsdNVBh13cPQ6tRvbyIzd6g1tLYS5dwVp541iehn6SIUOu84eF1WLJc3jfDSVZTK
qe1UpceFzOimiC++UsRRI3HKLVGvQCsj3erWA90yQ6G6+vytYOVin9YLSYUV++zChGSD94bsZ0BH
M9iTkmJ9v52iQkG0VLnplRr1KQBUaAknXxIacZ7fsqmP2ppySC/y2oOY5eD0skaq+c6RjbDz1m79
/gx8YEfU7Xn30gskKvme2g8j+9HMhb7WwU5wDLXqFHmCTIfyrCuXgM5yMilMgbTmiNYbBkvOh7+n
OR/ZP4iCFMRAQF3mE9LNcNDd8AV+33n2iezEjJAizeo2fi6FjIrbVRQEIME9SJehLVfLreRPaSMz
RlbbqXUl3fl8IklQNbFZdCExBJUFC7yjX9k3XpJ2QW3+iDc2JmhdBDSt5ZTAlYwMLJeEbUmzdOBE
iBsQrjNiphytYjgiZPhdDarN4xKEclIHHj8/ey+QKNiT/Xl/SMgtaO1wFYJkr51IA3+5xiGPuvVt
/ATEyFZY6gm5jpr16CSeFY/TQONmr6n4YqwACH9UifbNCw/CDGsRxGJrW3qNCeRlEFxtxD+i2Aj4
xGOscvcK0Gge2/1yjtFzh0klXAQamBXAuVBafNBVQQEnZzdOjGwleP0VGSz1F1QKKL6ccAIJAR4h
qygufLperTgivixPyA3j8siXF1pCwxpowQz6AnMCTkybeTj+0iNhtr6HtZnDGsgvkMXgZA34oFcn
RhfFnDzxU1oV7597InScCBpbM9t+nlM4gKqgoQQuqj15/st5h5vSQHocHsppItI1ZRvj3sejpozv
t/Uktcqa6wbCdtbevhR/8MbKcNA3K+TL5DEEDy2xfl73IMLBA0oJa/oBtEpURm/w/Mf33N53YJiG
lmUydT7ZFf5m18kD3YE+ruLbp50H8F3sJKRWEdfA7VrCJrv0zwxabLoGC7oToWEyH81yK9hvKzNe
eQD3QAOcGQT87URIduYm/QzS/cwnjOhlb4Y0QFSPZRb6F7IpINot6oHTuXPfvdze6qYz01ln8DPu
9/jcg0gpuPnrfsj98wT/tXERUApeXzOt7l6Pf0m3Y7X1tle1YbII77cZ3OAMIDti5lIgd203lVBl
8xLo+UNmBfTnQ+Q5zbM1c3GE82kEw0f+F99S9SPw2nTDFNbrg6CiPX3+cV65TPyK4l82GBytcY6r
eyfjNB2hXalFwudR+FZZ2AELzMasaAYv+XU1sLajFP1ETBX9fckRvdBt3yVXH4OnzqtXUDBcmGMT
IbGcvE2j+hreNhK07MHbFrKxW4VG2bgjslJdGXPafZt0+Rb8R1cqV6/aYWK3EzrMxi2pWpbhMQW3
t9YACmSnexnn6NF0axraRCzgTQ9F2olv89GK4UPDjZPstVsHdEvPMFpSXRaXH2AsasF/Djrsa7FM
QK12FLSWrvuvdNtrbZAQsYLMaxbZTS5V5yp8vUjEF4DFJRdMX4E2SiLnhH7tn1PxdqpoF7LllGYs
WYu5SEomDhzXpKkrmQ1BAvYkWDFYTGG/ja6DDgSJ0G6inqNABCmvYeK3iQVkDPNTse8vQNYEwgi0
rxTPY8mpS0es6PMnyL3AIJznGnuQI350cmEPkmE22dnIFJ1dM4O4Wnw5vLhWHfDGE1pzTjKGWDeP
KuG9HLyYHl1mJ0ICfwC6IrXP1JaCAL9lXSwVIGyDdUzbcAB0WJ7bhdc7SJgTl0jhDfOLgS2wGaNf
5Wopb7jvf7yoRv5kOqV6wVPfVAkghzcKW34UOv47Sqq0P/3I2ZvJHlmi4a8GxSohKQS8/J10lpXA
ha2zUiWzmqhKQTIxyBZNb4Xr91fEh+U6Arj6zMLjSrmeRCnR5gjNUW06/tLo3BS6vAYtJ7xo+98b
Vfoq+v+4rRunNCJeDtiYTsICGTHfQcGdW21E2LXDEWcuyCzfp3RnydbJGhv5HSMMrYqQYZrYdmt8
foKe0aXof06AgGSlGRMSLaTNvq/WpeFNAHPjqT7fxT0fH5lbghFbToYhToR/Svgj4XO/8yJ0f2SU
DQj2TKDjcQRjbNtJv2N2+WdUzWa1d0NcpRGlFSeSgjLBXn2XBtzcfnOEL5v46KCGHa+8sUt5zuKc
ANvc/ADM9BaM1Y9oxC4/p+r65ErrVxAb789kdKHscF7CpAFFB3fh7cQX3+EBiFqP8UGqgQRKpmC5
FDzZwoTIgcnVGfDD0HUOTdFhXilMN5NmIH8fh/1YLUMPK+m/iudz5/sqP65gCPvkimkOLzJzdI4J
CayR95IgBtn6NdOLFEifZ2TUu+tpEo8cuaP4/HlvAiHamIXU0sOjQU1V90mMWajDh2BkIznSk3w/
39qy04N5xswMPoHybvV5LekB8VfxZhpzvypR1OQu9jQpjCDDpkVuYjR1XjCkjCo4UbE2sA2u6d7l
JV6hqi+w40C3HhMTbZqWOPA7L2RABK8EoonfzshpVLPFSsUeh3PzP7J9lEYM7aDEgYwclNpUPRit
NQC8Gx/ceMRYfFAI3Uhs1Z65C9rjHotk3BVrP93xjeawF2dKpI5t83SzVmNtHhrmXYGREUhCFDcI
IFz9M+vH8wyVRsKXyIyUEosd5ZJDw1RkHhB4CJhsOKWekwaq4Y7RAucktqPe4oAGoyjWgYKthuSG
pJ75TWNbPU8iWJ8TKpn5fqGGIWiOoo/p8oEzaMC6V2hqvCVzNSymzsVL1BhSYliuk3J69ojM8r3B
l5xbPVO/uK5jCi6tZxhD/CWxBydq6u+T2vl/7cM8+SFCCFcgLkBWHaZdjnYfZY0f0BkGGURrEKqJ
ix6KptgKyy+77PMBauBzZipHQMeL6h21mxwwULZIgUafMyEGgOF56DceDifesfJzXlAyoizUY91X
onZYbe15Hu1iqNCFQG2VxRyKNsdBtSwNy7M80vo31ZzOgVnLmUnE8jSNBAicj+U8wmh8jzFViuho
+i7jGs+bb4bVfepCBcvyRf1tumlGK1VbGgD/5c4+vduzrO2qzhCmRCqrzgwpuPyRltSYtbtwJy8c
znuExARTXZ/gdHdzsr0bKoBwwmb11Li5Xz7t6r28Pq3YAcQLLQi4AfsJDGWGnAa6EuuqiGFhjW+T
FJOUZzZJmVf+DyhemzRigkq3t9nI0Z4uUKgNMxQQkkb2IMhA+Z+uyxNlvR4egPSTYPHF2mqX+qaM
c6ksM6XHVwKaPG8D7X6uLXbd22zxyWX/EjZ22DDj6vrDQwUUIVx15rCsSNLW+4r5D75qdnvoUyS+
HqjvU7lp/OHa9Y0c56GbqYD1xcsPa1WrE8DWVj3OmqnulDO5HLECC02tiuEbDa8cqLYXkGLbbgjR
l1JclmDv6U/K5wMlaLRKmh843DwcpfLPWylSGW+SfQQPCbCqnRUwSpnVG1zvCUarppHYPxciczAU
7jCHlkdE8G8R+rB4ux0mCPATMLqYC4DDgyBf7HvHlvu/AnYuTt36dCOVNkHjAJS+oqTRLr4boaB0
gU4twjRtyKq7yrGBZXtXPhVVtZFDTXdMbg9W+AXXKxT+IySJON2AYJ7VtYjrusT5xcEpYjS/Y5TM
YxGvz8CO9pzalY6rJ3i2/VBb/GVKSfFr+24ZzKzeT+mrFtKCjAkhapvIoRlc9p5qPvrqvcMwZR8q
OZ9eZHS9cIo0hx29GyNTWjbyiKGyr6r3L5TN+ms4LQic7EFeXbqiJgwA0XvZdK/FnmqdKa6d1ekh
DVn6seC5ML7qTbZvtNu3KHDMM/ORe1p+jb+6prSACJqQDxar4lj3d14R8qTMUta6BM3LJ/LlIBVa
NmXmCDpRHBiA6ttg0sqF3LgS55oXd9CqyHapg/tuVKnYI+QRGCs9cs/deLO8fUuoAhrtEGcP+n0J
IPsQ3t1pC9rNDM0+63xarY/HeCV+6HLQPC91Qt2LMcG7Ug7NpNea/zJ2l615lfZZY+37XKM4BGW1
gFVF+m+jcQX7+wwI8gSjd5DlJBEktd4PsJjOv0ChiMy7Yj+rbowRHTnyKaZwejfAC6iH4ZFOToil
X03RhPA6YK8+q5u1bf8mwTkfdfO5tPvo7KOmfyyq5TKO0iLYjIYtajZQQZrli+RrrCE1wpZybKVZ
Ou+iSQ45zOccqT9l2JYtS6lcmr8EsXP7hIsSlEs5+i9FqcLWTCMRxhm9dqTs60bY2BXx9UYU6X+o
sjtgEbDz/7cafUTsbTCv9Y9c1+sDDVupi75FE0YbywDKCohKXhrs0Rkec1HxldZk07bXUHlm5RLS
NSuuVhPHOwkqZSRKA1PSJI+WkuJ16Pib7zf8O/Jemkw5ZG8pNqg+SUAE0/HujJEaQxrnsURWOAFT
823t+j4m5gI/heaccUfuqaXJMK62n8Cwd3H+Xv4ZsaVjJ5VrlgtDX2LwZmgnXSoBZ75Qx5cZ1nZ3
AliVdLA4lZRE8koQ2fchaGH5kguEqja0C0IQ4VZ+xJkOOPkwSzCSUdokT9XbvsuUG3vtov9AL0CX
0SsrRW4meL5xea3novd5yMNzmlvYWCg+WJWgL0W5LWrs06q8Xwt8eLpwEdpGRuMfbzErXYdfz7H0
HhKNfdB3i0W+UCsyBNeu/8Wh2BPUtPiTpjyXxJ/c8tv0JmES3KQnNyuV30kqkOFsTGWwiNw94ozd
YhaYj0jFdrmLVyVFVz99O2xF78f9bPSaw9L3U3Z6VxGCg0clK+Qi287es3unVTSMSKzAnWATdjiE
YWlw+V83ddQ/WNcuoe1Gp1qohCafD3MwBT1WdCFtZ0PmRdMrAPP0GpTG5GaLwHdn8sy1P/iEPuTD
yssXcR0fKMPfNcIIOZoQDqj7PWApHMWR7jzPNE215JOCr8YD7fyNhstCK2Ux/96uLmTHQ7ywnPDq
9iwA9pj0HNkH5QDS9kAG4S8LPQIpxqqrPGvV0rsPwpUTqIhzYeH2cihCtTSCxT7IiNgDZKB4nQWS
WeU1bTfdMZH8We1scvDWx99L/mCkI2Caf7F50fWasHis3JAmimBpiUpQpGpRbJbnsbnUlv+CaeDO
g4gIzzISW2yoeAsiiYi6Q7JooXmJc94pxOObZyOTczn4oT67mWfqgi9k8mWg9YVAS00Rucd4tJSM
bm7RRq8j5bwlFKrr4/4mshFvoD+2dvQL+S1VUTIvLbbrDpWHhSR6WIm5Hhr/liDs9wl3FKyG3XD2
au1FSmxF0uw+cBCvqRUtDWAHqJ/L0C57xiyk69GDryvtR1fvkjpu9hB3LBX1KJKl7kELGMUIvZTG
ajJuWTCQi1EF+3A1kKmsOe85xgMSKJujzpJbNYpa24E9qidYqlaQWqzPs/zwqNmk9BK6we/lLfID
fx6OPM/FiQkOaT25QHEjlsgPRu8VlYtngJCe9fnvIhYYiOYDbamg1Is2NyDcwLSb7ryhIdkGI+5e
0y9G0zrZZxFtDDDj+84jbdfR8N1d3890UDMOKT6ds8DyXLAa4j/ukPWHiZpFdxzJI3vgd1YQNVh/
a+KbTRcjHpVKjwUYip7IqFstWp4MV8IakBy69SC13m8oMMNk7fLAlxJUBTQ8qZaxZlYXXb95qc/3
KPIRg2J7Q91qsmkkwSQ/5Lj5dp/BeU5x1iQ57WccMWwk8UzBhi2gs8ytVAheAXYS5qM3X8KuIlkr
PGF9lRMvDSRWIkVYMOlag6ncZeN477ZuAg7ykjzL33wgnCrqtmYH9fVXz658Tb53SJBF26oE5bAs
fD28uoL7GSyMMoB6LBJojADzHs4QXqCsn5jCpnb8Zr5skYrTTFvAWEq271wlQqfVYRsBkqJU3NyD
lP/pLnrHHlIv6/8AgPO96PC8NRcLFALfFxdR13il79oOwgZIVgrUJ6hqKc6xnR/LXvWZdcTz+iXN
UC84ORBM0hGxjysPHjoj5rSTKdo+4sAjV2LnniSKlSoPiWRCoZZdoYeuo4NozN7kriwN2UI70yiH
zDVFsP+2/I4PfChxiBHX4DcjOOHyYBvEHkt8lj4aLakL7930BaJoM993pzZ40uLx9v+piD+OF17B
nQFTAu4iGO8OQOIOWUNiSibWd/esWw7ilpLd1fT9oqYlCe3WIAn7oCRs4zgn/NsKjECkLrDngdFP
aeMoK4tXSWGqnqK8LdUAx/R5OD46I5FxsFsA7f3T58VCTO+HFPlJ9In9MTpmLxi59Yxp1+X7TOnZ
UZbY0rbsRWv4gqU3USbnXJVThEK74/UbtJKxThxOw+lkMp1VMKKcDgar8kIhPIIH4eIPNc7DR49d
sY5VPEtlcwV5bTE+QXDn3LlUhBDDCOnQprMjCNC1Mo4MzQHd36mBNQnHPTkkhaapqDOCg9Wk/4bu
a5KUO7Z3cJ2c0ywDvIZRtcK+LMSyEVVatRHmkkvaznAttjyrNQ+dTgGrsvzH+w8dmJ2af2QI8qdC
xtdR65L3qYTMT6lC+6qqSI2JzfnjsSUqvOeS63VUBeeSlpl5zbctrX6xOR5u6a6rFwPQsuQ1v1FS
p2ubAr9i8MOpRCFfr4On/0L4+knTo5HNi4IKxBNKne9cOBTs1u+TDw1FtG0NAEgqsSvka09hrE25
WjiGVj1H9g7xBsaN/OrCMM9IhljBjFlkHAt8bdruGaQniubzik86KDCNK02UeUgvDnYWvgwnOaS6
lVsUoKMfEHFh8g5yWV4gWo6ymay0N+nS/f6mrrpoBBi5Kg4p9gbvwn0209HFBTe6l6E2ZKCpNvDk
31eOghWfQmSB1dsN/NLDYnbjm2uhuIsIrqZrKzMM0MoEaAgOr2gqb2f4yC6gH5gPRIku0jxaW84l
6zMGJpGK97GF8bted5ZagC5qPetgKKwi7dGwnnr3K9+okOhS8x9iGcXP9sOfRt0KYGXIqUftzkNW
vPSgvtRhQUM+0mcgw/yScWIrfric0MGz4yyORytbHCsG0XmugOZQA47oYbfg+MF0K3UgO/kfWjSG
VVwZaMsr5Qcl3kqlu5rtY89YWzpxxye8aqrVpx62OiDjRYeCcfnFStAMqEWRSp8z+S02lZowSa9k
S+DpvmutCliQ9b5+CrJesWddwRZedpxxp1cTIwfPVNpOvnTL1H9FsD2w5CgdaWI3+guRMgqgZahM
bY3ZCWkAbVFQQeVgd9XsuZ44dU7Lvg8ao3rSylVECBrji2vE0QggNVQgvaOYyPLZic8NNQNqphG+
ft95uDubpRyzxiJj/ftZB4QuGiaaru3txRUuT6GgfGpC+VwsRNWdnec9nkAGovz2/xXnaoWvz+Pr
C5ezjlXz5fqBU6odmbDd37Fs8CTc3MhdSyFSFjUfPAFcwbMcbkz6gAaIQOnABvgpXvVWFPslaoXX
isoKGEMSmHac0sGViS4i9OmDdalVik7wq81CChBFSK1dkbjAEAkZ6sEhSbublMgIz0Esi172bmiw
3u6la45Ah0pjTDWNBLp/dEAYqxQNFiw0DH8OtHfbDb02esO8s9RaTWUO6ut5zGMqf7v6Och0FqjC
QdDX6FeYfB1ZwIdMMHqVTVNEv7i0co3c+5APlGxcWSSOvRJEJZP9Zz4pwHLslk1KD9BGwjgZt2nj
s3pzQArGl4XgQfOCHNHhVKUhYqdC/TcCnDMHuD14ZsOS3hNnfYZxgVc2Exuos8mB8rasvOYMYIkM
hc6jb7p8FN2PDvt2OHgeLe+KIsfIX0BjgY2395p40srvEAtjetFx+hPh5KqjlDaKE+ChLG2XYjSB
yiNPBo4xG/+1+355OIwomS0AyiRSo3g7vKfiFeVXgGeb2nnB0zpMk44OB7VkM7vFeMX9NNv5Lv+j
SN6k577QFJtxAyX/mZVHXAPVOsFHF7EthGWLdbXO9vbnrtlOM1sXARvojNUGTBvtaG8Ph7CP8fj/
ed0FneFzfej30cxi7to6jPE0nKzZB5pJEB/MNQyLgopBHE1SWYr51/iGS/5o9uclXJ3gHBvQPCQM
iyPn4UD2YU/o22qxlTq+DeIiZFVO1shEcDsINGkQifm7JTmRFwtTlLhBbY2/9a2YjBnCUavjyzuN
e4dkKbNdDKPNhANum+hg8HbVl6VrYDNDP4mNrVxalBAK4M2Q14N0VR4xKhSWAUdzUoez2Q0nvRrS
PT4ADKcXwCCy3tXuzky26DFJ1lZj+REw7jKESs9MXlFMmO01T9DTrzxYcOK5H7z+3glGr/e+FAOs
csKHSYIQQTiZtIvu/BSnFDAhNuFEV1zdHsLIuaSKxjqnq2kkN3pzcz1c7eipJBHvYisw9WzZ1oCx
oxXD81GnONwAvXqnNDD+6DZH8g0oXDpsSUuI6aolby+1lgugevIA5lmDlVkuZE3srXWsXGG5nT07
EiBZf8oOIdnyOyrcN8eYwwrc8ecoReVrum3GkwMZzx0A3B0ckJBTJKEdX4L5bmj5VxRCKbb4dyTA
Ot8iA5C3fs6rS99rURo9LWbX9tjzxMhysi5EsEWJqrJL360WFwMukhKCSsprSOOgTbIvJNXRmOCG
yPQ1ErZaLPLMahsf3eoC2/BLPHMY9Bp+AskI6Tqn44F8C4s/trey+3oTLHRnzIsP4qyNtpoYaXcK
p4qR7ODQJ8Wrz9xxRrPtnvMNFNN1os/lTHKh9mJHFicCqKoHJ7t3H7gsi2Y1PdWxpFi6L+QT4+N1
G3/yK9C1gPzD9/1bDn8YpUB+bFo5Eyexrkva8iQCMEi3vjxqDgwJCGQRLI1hMM0zJ2/1/mylHZSx
seYep/sJK7iEfMna/JxIXebSyIuayyhlqllePK4n/kB9+LKfwF8+Z6X4gtZvu0LwFHFxZ5FJFWEa
NSScdZJBqWTEtvBUw/HKYHawqmrIZOvl84mE0I6xH6+gVr5Fdvj4TwXWl+jr584W84Rc3ipqYGwc
VBNzaoeqxMK2ge6sd5caPHLhW/r1lnh84+zXO52wBhup2th12JqaOlNSpKuy7yL5H/K4ObvfFRxW
/DoVaoAs+X/Zd7vrn5GpO4Zf0vATa6X6yl3TThVOsXIU94B50hE6nABbaUXTBMESmj7GZ//kSIxi
oV3QWYGLFfsbR4WUKNjO4b117UD4QXZ49Kp8+9qOV2bBpK8MFFBDGN1f/yrk5gBy5wqyhVYhthXM
IXt0FORZu+H/jtV4km6pIAsvSAzc/Rgiuqg6Yrz6xNlrvkLeP2ZpGaoiasSLVPJb5yd5SDB3JGv8
jAENoF72RrBaLssNpAJFwO/0Z1lwQkIGHnZDXFOf7XdcXHrVl2S9zjxS5nIkLhaRJ6rt/Vo5sp+4
VUK+qrPkr8ql+8xfofGKZonhWXOcrhWzxvBIL68Ez7xqM8E3z/fx7oSPnVOuq6YfRrF/vA0OZt7M
vC+h7sO7VlV+k3LDngaNn9LkA4azKFUI8TdVOxskg2jsrBV5w4VIrESZiaZT6M6v3NAI58NnUWF5
gIFz5iz9/T9t+R3nhkIDminlMQf16xFvo93qIKdQfEMNGqywK2g/NtwZ4mH5EL5Fzisa/z/CApaF
yXodDDuBldD9TQBtE1jDG1sJBmWNTH5wdQdwxyoW6QWtj6N5YwXkXKIrplKBg0S8THM9h0/atGKM
pT5q4Y05h7SGRN/fz5JECvy3uofMK8vOAbBQ8ADDeMxpnd9SvfDlQ/kIyikDXe5dyD9dR3PZBr+h
9VOO51hajnQvasNXc+eFhxIiePdFWdK9f3sJ/cEGi9r7nLq6y00FfD/+1n9FbVybbh6g4n7aF8Nk
y5LcNGFBpBHQKh7yRBPTmhKzBAUE2b2bHPT0hdaAJ4BYUHOnu/1CmJ2Os3mtYM26foBBYAdX6m56
P6T9neCnB85OLnjEIDX/rVd3ywNmCxoEyqYjnOJBMSeU5VxjZhpfVw3usqsC6PDKoCTnm+hMMUvl
EuICRVRjimPXOVmKcdzsidlPdUVxHfxDIw+hsTzvK1HJEC92sRYkzC3vi5Z2Dc2+fGnzOd4HiPgN
SOOhHYueiHPycdt3BQgg//tHBI6lvv4INxf90tTKxx2W6zd0w+p2RJhXs7c2fh6b5dkh41CRNchf
eso65lE9GsboEoyBzeNRGOFbPlLiEP4XPdW5+bHUDl0ZlVGiymtGcglRiFMz2b0N8TgkTi8DqpZY
T0NjxvBb66xTubXa0vaOZV4ssRU0cyfV2B85sH2vGSATwX75vQDZRWNSfVd5TBcpyE5mqn1cUzJz
xcy48Z2FO+GUunL5YRL6PUV3Vjb282ky66OIMansAiSPCSUiDHWo2Her80N7ONUyomzPpLK8h4Xc
0R/+HwWF18hlYRQTmp5rb1NFHeDKrdxhwHve79dj6CdXtdbFSGLork/nOCnQwQAGN+Iex+O/fC9O
0rtPczRKNXR5/JYm0VtVOzwOinIFcgbXKv8E695irL90PZZu/K8/ovAvJ8t2r3gRuDLuvstChJmC
DX4oTjjnW/13n5GTmkmHRzOzsYwZ8vB7xi2bVDALXPU7OkqgOtapz43LmB9W+HAJsrGtqLngbCfb
mQmqLkOFMMs0Ke6vlbEVRTp3FN+2L7NVUrt3H7GCf5JsbkirQaNpVI40T4s3fUWseSGKmFpv6rKI
GyLx9PygWQMApTaZ9zkCfSNbZIs4tnIluK0UKZgzAaWp/g5rujRZsDheHHbKnNrYDtSU2/iDfyZ/
oRvx6JKpPKdqbZbuq86L07Pr3r7B2/kBm1s8oZbb6Yw6Hc8mspAZ43pnQSwiCQLFtVpdV4roxKpm
hIC6hH2xwQ1RpE46W38cwb9Rg+33RjUAd0q0qdbJlOvSxtj9xyVItwYIReJnbUVqRCFOveTsJ/Vj
f0z3d5Df7B33uzCjG5+vH/nxAMPz5bgAGS4Mp1sY9U+QYx2IRfK0kGZmM18ZyhtUtcAjAS+2P2j5
B0jhkwTE8NwqGev0kayGcHGjjp4N2Zqctqc6I0D92zy3jbcbgPvSdlO+CPFaqomETirT2bZ6jAvR
k6eeRQvNcKgQPRzq9ivgvyKv3hfCkx1ZCPGzG7ehTu+iKufPo0CxOGExoMAgR9afQnvjDn+dYT4F
kJC+QmoNJIxC/3LhYnrb6QhGERwjVWl6zRFyZ25FzdQPc/jGvNv2FXCLSAxaGUUWWpV7w3TbHK8Y
Woa26SuOaTU3Tafb3wjXCHRAwvQxbpSPRTQ878EaClxllkxU5WzjWeecCeNonuFdfR5WJF4hi+uK
IHyksdi0rmc1AKEf+GCN87oHZhs36IdCeDpHva0nhWAGC8LsxbXs7RnPlFglPM2jeb2AH9FqEQa8
EfNu73tFEcg8yQTk/cxKOOvL+lNyXLokJGzmf7syCe91evFkV+Jahoxtf01Ws+pUWdEa3TAuBEeZ
3FRp0bNL11uSe6TIZ3CqF3k7NU2wyZsro+2v/mLtt3Vbtv5ss3tKOvOLhcMxxV0vs8YvhJXmbAIi
iVgbx/boirMmMvOAlLeSY4yjV4nTH80uzvilf/1thJFcfZsMqjoyuNZsdDWZhtddTmB0VuBSzcnU
JvtvkiK9odrbbx98Gp1LioQ2tPjbxxSeHkz1yBz7L27d8MqiCPfJrkohr0Hi9BH7HnLMkI7qbiNf
m55GskPAynZzPb2agCUThnYYpzUhrw/Z4GjILXLKWmQqidAI0Bzuacyqdw1y5VL0pcDmVrz1zBDh
XNaVzZzYcvniopHiWIQ7H4ASzp9AdqitRv2Y5LkxgUKFW9cG+bvgmbh2AfzWtdmyawXIzGqWJlPF
ELiRPNWoEhh2y+/Vn++w6rsejrTBqBnIqodiF9oCR0QVnuZsDDiD1MLGHGFYIkhMUGSB39lH+y8F
4tS89eNKWgyIKBDcxHHgXoQF5v1HB9gy/3fVwaaaBX4a49q6M+moHdfKXHzzY5ijsb9+uqa8WbvQ
DGkYFGOVqVJzABFpjhUhIUpmVkpQsWa2riMEWYGb0/H+mDiCDPecgEnbBiAsJN+FGunw7i60kd3r
wIDkT146RbRrXh3X8QTDhUdO4O1/K9HBOT0TgUcVsDo9uHt0P5dYs4kX1UrKxCFQyQajpdU2VJJl
Hsknl1BA2DilA1JptXhQPOoIjEyK3AGT4hLLK0ondABjckAknv70MqGdJ3MW16bZnrt9LxBnolzc
VA9hOxwLG/duIwSbWnli0fiMaQl5a35t5m4tfdRj6f/R/8+KvfGEMw3C7+4cq7DQRKl/pDcVi5uU
4ESZZxI7jxlwQg2FdbHWI1JdmGyZ+n4fHV9Ctf6ti2iQhAjUHjfgLCC6EZjPUkXpC/6wZXJJEnW3
Mfk43VAMWhw+MLabFdqqcYwWUsP90BsJXskN45nuGkKPZdMn6R+yOYXp22/wefBbp+BSDES47e4U
tehrdRtJyXaoe8/VOUBZzsoSzG3DdgopaQrNY02ft0n27z9RQvzx0RqOOc5u5iHOAY0c3cFsu0es
/jm/zs5MIIeZ7skspe4mI1VMdRIT0cL5ZvgWvGEGPrjc8w52VraPV3hUERwjxn1myqyx0k7ax6Yx
O+zzbbR2tOg6oIMJ1+SSi9t5LRB8x+BetZsLAVkdib1EtkstGuX5nfSxXVrUeu5kTb4l+y77bEzy
KxWTQ1WnsQRszwj7i2FCfHQKvZKPXzBkTMBXTKOR/0njjACH7B6CQ5mOVZ+B9uEyxOM5AANuMvH2
czVM7l4fJqu9uBlbpTrk+17mKW5r8mbMWESSwGOkue+tJxj9tVGYu+xwoMoa1XTIzsfM+6fCtvgC
mkJDfzlr6b+EC+7uuSdYG8OvegOkP2C2cXNazqEnlMNK1I/RwRX21J6L8aeuVlnHwoU1yfbZJv3x
VYx9Km267b209qu5gf0Vf2fKy0ygGfUHf0VVYegjmg4NBPnEhwrIQmugqtbC7nPqgRDNJWWf7C3K
0vuKbC0TwziGUB2QWC9ktbeM+vGV31Y2jQ9QBBSSaT4LCe7+HQGe1D4uApNv6fG9xCJ0sbpYfb1m
MGTQ4hNuAzraaLD5DCGdNq24lhSZmGT9j2//dJVBDUFEx2ZSFHxWOflTmep5o4TzjhmBsCEXNDYB
pffDifaK4Fx+9a1+6VOd/9e/dchnxPHb7s41CL1Os26LEFLi7ISRhoP54sMkxNlBvy2QPHBszrB4
Na3GUOz0+i8q+VH/BnAi/eXTpSQBdU4dquIPfcs6wVPed4ioG0qE2ODs9QLTyy5N3PkbMdeKojbR
sTzEH1LucXyvVmjG7mbLu6tsELuFPkyd3gfNB2QYpFO1x2d7ZDUwuTC8UwX5Tv350vHqLnhUdc1q
8W2pRTAIFlBQu5P8cIK68bxcu3RV4koLNZpTQjhnKLygsK9vebU3WtiXwe91bQB7/Ey/yOzBuE+n
fKgbU8+0G3ngGFbH//9JDTLMq4EM9naYtlZCj5cc13elzDJPhFyUkjKlt9kOmL056hFTFpudn3Uh
oWx2rxDahf1uBl4ouWN/EN5upFzZ3tzs4U00XdTcXVFCAPKVLIQBsDW67dE6XaZI4t7lRHXcIGiF
UKQ4aE3UGZydAkscx4fJOHgRjmrJOoPisgPBarqlKvj23nkBxuOt5ScLBUmcWk74J8tLc6g7i2ZU
pcH+ugkupSzC6K5delDkVjuRlQnzSib+TJULWUKb0m2Xoe93TWhwBDv/pYwG6tCNiE+uC3d+IDTb
oChuinI5xO2NMtCQFyEoRk8qJS5FX24rWqznwKNjFnEyvsIKx3M8pIEeHvzF66mgs5Wm9rgEMkAp
HWo3ZeC0oYDJg1VBUVQo0hmZwzvIK97frnWvCDv3zsb6228VhLJ6MpoaaLaSMuakPwC1369CiLIT
g0unbtzGsDKIwKrO7NJ7OTj5Kq1fAyiSOEOBTm3L87w/Ti6RLTFZpxNqPpINufvBbcWdK8qJHIxC
yeLnTYLR5mhuLQJWbWZtjvjl5KffF6nYtUaos2kfa5aI2gYEA8VWXTTvbZiXRc7UjEKvCfRDmM6B
4EDiR/a7WqYRlj5a1iIUFqQbkUMDvgb9+sm/J84cmwO7k7HD8UzuOH67I8I1c6LInAUep/nWAKUZ
/X7FZ0ziMCOSc4nudKE3gYjhRkNZsP4iMR4r+26e3WwhOGBf6c2cqt0nWExKES1GTzgkgp8TaQzN
u9UxinS+6RXnP6PlxejMw7twE4FQqW/2yzBdeAKIVCqKwrrFFKpjKLeqKfK3yT3y13hWcl/v5VZl
m2a+26UxxEEAwf71if369aeGZ9BQaikVh5XkIccJtN44cJnu//yC0brTDHmQpBOuc2rRL4Z/dwjS
jnpafnOnghrww2rA19wMPfmuPX4miNrZgi5EslhkC0h4lHflejvnB772Vg6zdzCmDk01PYu2K002
wQecIZogUFYePf3c8lxY5Qp8Bi+EOWssM5ta/beOWsOyv4K4pifcbn9Tt47CsZlX2sq2s5Hay/hs
i/DZGLX20Qv+Qq5GhCrVbzT+YvQPgvukDaSSxXgFYe5U3iAuweoYDhyLUxLotwJsrsn9JtbFfQJo
jCpoBLGL5vcY8WNSm1ji1MxJLZrIGn4cHY8D3Cnt2rPsO54/WAuWW4qqIAoyamDAqWGaV5MkmpI7
Tpy6Mm/QNBeTdknTfT37iahR53A22mFwRrNyC1oU1eB7kvtG/oTrWK+Sr0jMDTVtSuykwxfFFZ6x
LnBhUoFB9n358jlMdDcLi/Fm37Jknw3hvIrdbLDBm6Yr5mz+eSuUIh5f+dT5EAVGOeH+wA6yAmuj
yiLKJzP8X3HR+oNAnMOqZLJMCnjoPmfk2hKtIxKsNVqjks1eeMsrhob/WikT7sA3YUYPeuqWNerW
njxTxhmhzNOyqNN75F84wdQUqWlr6UfDIunFpdtSa//qCwVdndne237sNH0hrwQzuAHm+qaSHoEg
kmqNfU+l3VjjgybtdFGNvPabVhG14jq04ZnOzvtX28hKQmODMxnmmMr8SRyX7lFire2+YN/WHsnD
URO6OLY2py+TAe7bH0Sm+tQypFtp231edYm7cr9mxOLALYdEaMyB9CM3V3OsJ9wNfxtSGVRp2yo9
9RmL5P+imdc3dXm2S30iH7ySYrVMyGn+nqvsz6PRRTjDaJtWiaJhZi6h59pXTW8UKDiotB82lmKo
TOXjMiPtJLpoJDbJM6lKspR5+NcPrCpvrPoCeSyIGsiIcjQWFNOZW3N2ykjqk5Mji7rqHMBBAQ1F
+s3hxwL3jEFEPcR9XdMxnO8O3WkmubDDpM4Z61ASStGNB3irpiAA0DZfgNiOqf4+i8sSa7iHne0N
T+K3WZ5GcOYA/S6W7zw7fWdFlEIE7h+rmmJbTVeH/1f3NEUAriAMlthh23sKG7XcDiba0mfnQlm9
DZeSHJs08FnTcI7k/GtC3DQPcBkEerl2L+xoUkVM0yxiuAKiHHIP6CQLJBejL4iOhRvDV1fCXBM7
G8Y54auNboPwiy2Sygq8hcnL5YC6Q7uhItl27Gn2VOVmKhpcKxVM+p753rk7cVAsdJDVUPs5jp4M
jKX13HZB3dcTvw7c90xDOQmqHVx+eZqPVodoGZgy1FeLqdcqyGKth9kRjhOuxd21LJAm4C75yLqI
g1SfEi8zKxqR0kDA03NNMSizoDIsoyV4o+9RtoXF+z46TgF4F4lHJZHbGAb9PSquLmfLHaLpo2Hm
2HQTCBudVjsI1P3MWGuCUTdonI+gijSF0z+FFRxNzUDazxR6t4mSgTbRgZTna2qyQoo5CsPIpNYI
gwX0S9huHlgm/R6o1LoV9LSn1tuD3UrO8/J90jNutv65+qelk+kafvZxrf8HneYQU/8jNicQfGtX
ThtGsPQmOvitlBjqbY0e0KcBMNbDlCqFhWifnrRyAgzqOO04ls5CVVaPWzJavdtriAYiLcVfNU4Z
p/FJVnjJSziOnviCljDfE1GhI+Agl1+CfzjlBwGaGicm/P4Aw2OyFLDL4JxT099w8ifRh9ioFHmH
tW8/sSn7uhXDVuLWRB9ceXfLWhf5WAysU2tO/V/tNw4hcAJo3V8W2E0BIzFAgu/qCwOi0G5SV7Rc
reGfrCtUaXJchCIVsmfKG2Z8VcKvRkYv++DQjV0sWrXJ5Rz3vKPyDbls5XLFEc48+Fu6VqQU1TMk
avI9KspYVFCtVheesR/9/dTPchkMT4It4CeP/Y5tcNZhgZ6wGlrpBZ5dGKifdAhv7BS3HDQoSxtp
94DgBWceU8CRp6JI0jigM/6ZZ+AQSIzTDRd3v7bBbHSsPxj0VpuNrKJcFH8lMb91vmRlhbft8Jcy
T42q2CVTf5T+tGoBewtR7YGRtIZOQ8G+xehNaWjkLVEVIUW76jw3g5BohBRKm4KyeKPj9S7tT0Wf
A4jSgva0qYm2FJ1ghIp+MIhvMTss/EMeLyLh4lh1hdiM1nzjkDksZWfhXOoG9osaYQqVPNpiAwXm
csKEawA4r07zcdZgCTpHp6NTIEwfhWuKTG6bwrbY5K8AJXE8vW/+n0ArNWDaKu8PdrzsFrO+nym6
tVChkt+GJgQHqrfiEjViDdww69LbYsSa0QdyLA1/Unmw1w/dHgvtr6GkzrNqGOKFZ3UieDIr3b9S
vGQsuU99gsfBjidQ8DwIoC+PLVcie1Mtfel1JLeU1vl+kyYKItod/yDLkcLiq7Freo36LgVhIxK/
NPdaZoRXdv5NOORJ/GaMU49H+MG5EjSOoVMH4HsgqCKfiQ3VomACu/W1xBoqV5w7O/85EcX+QWMm
GZr+oLEP9e6XRMcx5zlZdnWt0CsNx08e/OcBe7AJvztnfVrnBlVtXxA11sqcevHZtwEMZYsT2Rar
/ON/1Huivkr24Xz/Rdk/vH4uY9yzelyOTqpW+W0Jv1uw4HA/FYBhEXfnSY622FCWP2tCBQf4YCty
U3cEVaRUBoxfH7VIcQiJgL1It0X8VtJi6BX3NPqK4kEbfaVs0oPyI2vPb8y2YGpeCJV2Z87p4G/V
JilXusmakOZiUzIs3rRBJW2gKSkp/y4dRKRfM3haf9HlX+zVu2uSR5S/9Eo7ki7HNZti3j5PANQD
+IGt960NfPWT8NYPODYcplLeEeI4ux0H8ySk22Li0YNbe5Fc7yDUtJwkWHkxiSS0C2OLoQCUXVgC
uwHy5MVOIHbocup9vr8LW8FXECCgTzUWvfhD1S6bsmQEAKVb5yaZIj/zSKfDbkdD3UzHaJ/UsVVi
8XIdYrUUbw8Cou75VkxazVgHVJz7kZlh5qIxeFWTfUGSzM/vTGJQqlqi5heaKuufVBDsoTPrEvdw
FQAGGWTjGCrCUBgvIoxDm6eBI1jvU+W59eHHMA2+P2zA0K4JciOpMcKnqdeneGNWj7fgmyoJqlEP
Fv6weVwtKzGNJT8ObQ+PGFM2XYB5RL1lp8B+iseOxm5IyztS6jxJjn0+iMtYi2ZZgtylUiWgYvSl
6+RIRq1hdfkrIxqS1kWzTxknMFu+uTIbSsmbqyZ9F6CascWyGaN3hk93fN1L5mjoQevuvwpcOcfX
r6SD/wdGPiM4b498cc9kJpkYDjvP9/HZnsT/Kqps+t67n0mjTVU+dBm5+6R+Qq15CMPSycQkCHjC
/ta4YbynkzaJ+OdYElBkpeThYGhy1E40TwQLPs352aoexjUXOBGY7n7dkGShQhLRdb6+qD/WycTQ
sGH/4FiJyUHGkfFFqs7M2V1XppkUF7aIIE9zALJPLglSj80yvQtbZNLQiuT/bEvY1hBacflTUmvT
0IhlSC/fNMk3xaMFFavBmnFIZ2N8pheYQyAa3iZfDW+MEpOkSn3oX5A+Mu89IENjX3gG7bOhPcFq
7gZRMVxV3Dz1eLO8smNcIO69pmYX2ILUocU6zLtsZfem+IN5PGt2y104XRtYnLYeScBv9LfV5utT
8V2EMNWja7VZPkipny0DCavB1tT4ca5ki1xcZLnSebJhalw0+AkrDEoZYCF4wCzytutLl0wLRv2R
rQprrZm7FGQYsJ3q+VexBl3sNE3vqZmeCgqUVD0Fi2KM1gcvla6bMlfzaF7mm7jZvCqSvTkfqxxb
WF722k3BB4CEh0YcqfB11PKGNkQGgzuTPWNAKchdyNTGo+DVOlsL+ZFk5M/R+RcrJVbvWALWrPfT
Uf3Vos3Q+TAuD9DkVj3o3SVE3sTUvtMHVQa2TdHwsPz8uuUPmOvWxS6GUWAfA1jeAVl87kU7mZv1
LsZYV7hcFk337cj0iMyfQULK0EOCzeoZfwh2DGMlwHiVUQCHwFTuvVJq7mVQoX6u8l5F5iw1IMuA
DDRUfWUwud4dfB3h+HE0N3dJLiHuzskLE9tlnNouuBWAGQG7tmhS9+SHOOWjL3tZ9xeoI93AuXPz
eaK4G8leVEgtDxCDbJgFAttMGsmVU0N7NdmxUoJbcRWpGgUgAOoXtRkR78yQNk2ct5/HgdNzZH7E
Pddzq9k3XbUulzxPm7NPGaPb66ohxvUacOHfoGUEHof64h/ATZzMA5hhpxCa7m1k7M4fI+ZAAhLX
5s86kh/EubSvlcc9EXOZSrmUphD7JxZ9RsToXNd14suOmAWDTeFb7VPG1mQPx1ACbYeK25TZLvCq
A7HvnhASjhTwgqtZPsvo8ETKeLYHt6g4H63rpQjUt6zTIS1t+++oC/B1XYQFjoWLpmi6iElOxCxb
DYtFyPk8o0sJymW+PazdHAAmiRyO6lGbgbqmnhFzWBthk6DOUA41yP6QpScj1l86y4pZxTA0Pxp1
MzXNEIoNoG6R1pgPSty25nRiKkYrbCI4tQ7oo44v0rKKHMAVKNveJuQZJmBJmMJYLyKi5+5ejGRy
PrnMiAiFPYDbAGLqDWn3wofu9Bx0dokAwJ4avtSH9GJsOmuEeVbSgEB2MLgrt5DMOYpMFJ+2WiA7
9l8eByvsgLSZCn9THQmdECupo1DbYMBe/GZiXTtuWd24Egg+kwazJeLE+jn+ye0QFQI4ScWzmX/7
Ly1db6GS0gC5vy56DAe4FIgEFTm0UGAiwszBfAy3yWpI27iYSp3z0//GCnjZC9CGqfNs9PKWN764
9cYhwBtwcLqQ+ulMx4ctnNBMxWyJCpIMemBhD6RHeGbbeXv5S5RvVoV4VHrXrcvOXteUhUF64gxN
9uVG7yMsds9j+TC179FopsGwAOtrc513w2P6EnGO9NAavr7YaEycJrCK4AJmge0mePVb1KCb8D+a
WrZelhYD2LN2n62Y0RqAr0dSAH7RLBo+K28NNOPH81o8ovt6tnfgNJI/zYUSCHqnlmcXWH774Vb7
gYg/qWuB8HC+/VpZ36wa8YZJIyVgeFr5sU07+HwN1puFdQViiWtfTpn4SFzEgGXaTavvoJ6hiMx8
5J7nJdz3o0rWPaXlmqDDnTO8rBI4tVxsVKXg47TNVw8e0lRYm6f3N+rmopt8nlbQFP2kOw40k96K
0xDLj+ck9s44ssFYAzl7XoGZqI65xl7cl/80hlEinh5BplYjM2vWYVmWOfHZzOJsiCE7+JINhj6/
KCGff5S/sgKXBmQAJcImpQTRV/oFYKusptWFyJvUvR2SUCr9Afg/DeOdtTN61nklEnSVScOTOgZ8
PaTeDhbOmR8krxAf+XEweRDV6EVVyp0Y4PS/HLJSyCqeuOm59gOzQLUiJcOq5wPeyTnnv+2wmf+x
jJjm4wuWUjROMJ8LtNDbYtB4t1F1Gs1nGcEFrOSAKWaUD4JuDaqoS3FitnN/0mBI1dGRUw3EsHbu
VH+6SwnGRDtmTfbjP251FIP+orHj7zilfWFIXbGtgccV3n6/W6VdgJuXSprOFgLIiOlGlZ/2Ybcs
l/PoPWeMXX6iOuKuOBtZ9/L4QycnR1XW08vYIlanj4xNpDn+GiVrAYmwWw6+iLob8ud41yh3Kf9A
WpTqtwqHQTgOAyZzPqAgPypsMMbIrkHVPbHDMZsw8/YSMWNkz5UQ7C5ISbvREWhXnXS81SxrSl3f
7K5NML8rXjkwS7mzuPDZFXw+K06TJg0uBcUGfIAAURbMpL57DVdoZaZ06pFlAjVPivz290x/0oYD
LdDcLounzgfqbGeMp3CVOZmpkkRjCWn9N5ePFsL0cq1t5WvKUuJT0rQsBhAeYC5rPncfbNIdQTI1
tRw2gwMToLb5UbF+XUl8luMC4fXINw04Pv/fvkbh9ELQxfXfwwhdALrFKAgfHKBRnH/vPS1U4yZ/
tLwfG8i9tpJ0V0chLGRzgMYILYvYig12XbqmTQlFF6BrCHSrv+Kf2dEqhdhPc3vD034ciF83mHAA
elfvoZXWdItouFASFgPzO8weluLSCN+SgZOj6foV4poT+LkIQr1SbKzFFncDEtVoAbldQcgKaEGs
CVr+0GkzyA7IjwNaQOGalf7FmGMjm8FvuaQMcdFlmGCG2q2tXUi9nSPGFK+5DM04DAA3IyAq5B+N
vz69OqJDnQrpbcRw/od2LpikoPPXyr9M6LGKBOeP6lnKRGe2b2xtGr2XYPMSnos7sirmMyHf11X7
hCPM5YlM89Lo7lVf2+76LEqwfsiP3z0E3G54BWzuOtPds5CUYKSCDTE/IgYQLSu6CptPYSUfQQtp
5kXQXMlRrUD+KDgWUYXOQ29buAfwt9IlwZUBZUlrE2HMj72WLI7SuzcRMU0O1/ItvYyy5y9gIk9U
YElVWsCp8hhUfB53MbqqcZqopEuoIOShE3HkfwKLM8PYA/vC/u1iucZw2Wn0DotjIeVQL3UTfCJq
Qns8V4/ozw6SPR4+7oj2Qpqff5UwkytQcloqiUKGrNaSaaBiYhYdO4AJoYM8IrTm6+q0lV2JrqMX
B6cEqYDBVOE0/zhomfAqFPEttCX+xvPxgTBKIGiqyZzHKi9juMk6M3smpMKITLbFW3D25BluFt1M
EIKG1LGEIXCMM/s8fW0e6F1wMdXaGmYDueS0hxNXM7jP9dg/Mw9wZQ/GR4py64P9g1blXDgW9gx2
yYmD947mGOJP2CcPnfc1sIqw4cfYBoqssS9TnkKBiu+0dS3y/0j1zkX925K64lTRIsib+nrSLJ2b
T6kZ0tNDQ8jWVEINgrToPqpEZJWa7IOiZ9N/7izOyzpcJt41E788LGGvjovDGp6jlPbDhgB0zVkR
ofP2uc9QVKKeuQO6aW6OOhdjtC3OEUYpJq+3g3wgdxUBbskhiI6lUBXvvlL7qAdWIoP6R1K+oXCR
sZ2IllytZYl4rFBCoGfg6Gf1ut3AtrsA1acHuXGG8LglfZF/fN2NlOcUc92hQYwRyNDj3h6gIo8Y
f9mUxLqFxM5kIiKMzuJKH6wp4Doi6n6mDs7VRPT3KfJw4c0aQ5yAC+amSn+9gNB+rxJsN3ouxygK
OUjz3WXxPQGWFOVfRJMJqsnvLms7PTKv5Y1jBpBbvaxgxmol5RbayizyVqlb8DaygAIRXExToBh0
TMIKQtgvKuNPnad9vzD6zCZyRgVg9Y/zBKR7GCf5WNlkoQ6NsZWQqy8NOUBGCfdrqzPnHt715DWt
M6NKLIO9rXLC1ExV8j+ax9mSSBbnqXM0YXCiuo+3+mtkoLyL8WI9ZYS6N68SVLjg2tanUB0GKDPF
4r9xn1ZR+wegyRs1pS0RA+GIahCLVdhcuEquSlQ0v+3ScIuc6FklLpqUaXAX8eEdG3CsQTa/odS4
w4pi9+1u5moH4TuVwhRZblQGq2kPPkCzkyOGpRJFVtcVss1XbGWaGslQwYoCfuF120RrzuxOOI/d
`protect end_protected
