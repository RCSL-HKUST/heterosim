`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DVgMrbcs+MkP1LOD3iJ9tcYsrnYGUkVfbzQvebZi5iurGgkHv5pQH4BC1MF821ydhW7VL2hjbHMpKjrSZR/VfA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PJUI6kw0amAJDOG9GY6GiRMeLM0NXoltkuT+LS7JaFsvhMV4B8Fb1EK7VQJAAF3Sq55XoRgSE7AHpjk69nC8i0p1p8ftJ6O77bzHZyqLICZf8JSou6ZX0SOhYgI4tFhF5bEanFNXqNCGoryGC2Xe7JGA0ACo5IP5z59wxGjr6y0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sSR783FPRDuDzBYf21pmHiIWni3XGS2HP4CUVHRHCdnsfx2a5ybpcsh9zAtf5X94ckCkttSd/XrCP3mR7YeCR2SthnoZp/lgbFi7n0PYRcXY1BS8wXMK51zzSxTbNAx9sgesS63It8ejejvpeRiLuA3F4/CArOj7URVNJVrRceBDOECSPX0I4C4YfXk4EULQsjnV12Pk4IBIcwB5Fnea185Dpe7W2Di9ck8tf1+MAJwTh80Qw0tY+WtDM7tWZuulZHvEbOzphTZ3+LZjZ8C6+P9NjS2gWei1J1yzvn6/cdoy5S51AOfj7NNE3SkqfpzyOh4KSojTudNUS/om+ntvXg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wBgeQDQp1Z0B9SGtE5zIyv6Nvx6y35BHU4mQwsINSmt08cTR4mv9t0Fm5f7nGo+s/XZFgWeEMl5QPBUJiLKH4eXhCD6fJ/1e8VvA7GjMtuHK+2ETExYAE16e+E+Uelqz46lvxZbdl/H/oOxj2SaY5UtP0cUiaz2o00f6dHdRU1Y=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ne7oXOuL/oLO47NHo1uUbYTGJKpVc/n4b5nMH826v0ve5txeUCQLBXLcPNfnRJHAJv8Upw8OvQTFFvYSL4FX7NbrPjrIAVcmkX0kSsMAHk2OIt2vGrBGcJD3zHAZUG2iabinjVaokCaerXn5O890Xhz+a9i52K9nOUhkW2BHHSfzZl9dShkl5NhffR107Y7hYfMztymOGeJplOKdO6hiExOYAseZsdpvO95of/OQ8UzEJv7CQaDohpPqVQcmBAHgJHPNIDx+ps/zt8393vJvPAXwbT63uUjpMRqoACbHe4hv/N9SqE4h8GZ+55sW73yGdDY0tLdl1MghVjNkyrqFoA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19457)
`protect data_block
YW391t+WmdgV6F4Uv0HCrcOmcugnRDQohR29O5krsq8Dwmuv22iv2z8fjx+Ve5Ma98vlOolsz2nB
VQQjzlNELhZ20BSXRToUh6HpJ3DWdoyyEO1zrERMVEqpZRTdttGsMoQzcqTWvQoWSoB5RmQocA7+
YnAXA9ZZCil8haQNOnnJaL46ydrkgwNguwQrr9tA4Y8z9y4yXTibt0oW7Lz8FvcvpsP7MB7M789e
egATo6t9qhZ2xUqK0pM3kxukOOEo2TTJZCVjNs+yckkOLzsRBeASQq84xm0dfZUQnXeFWGsK/Arg
z0v0nNgvVG/wP7q3rqAA5CC7dJmM37XZVvkw2Aseor4Nm4bJSHhugb6v8I4ipLsahOTLPlwZskZG
wkUNTt4Sh2NQHvHFY+CgsmGG/WOd9ty0RH4FT/sG24wz3EeEJOSs8LaX43tjRw+UzQE6+34IvA5P
03QEyLRQuLoJ6MhzciYuRxZ99vgybnBi8YIBqRbLQfhRtZ3vFmkFrjknrbLvDyqiCxdg5W51upDg
nTkLlgtK9xWJ1rTioQDiB2FA5OteFpMWIdB6W/TKz2ceFY/1v8GXqR1+og6Rpl+HSQgEoaTe9keK
+puzqa34+HIJIJjtKpIyv+IFx8WrkC74zKP5RhUjpYPiR/OuWua/iMnR6s/ch0jg45Bst8xkakA9
P3IXhLG/FQeAtC9rV3IO4GV7+sg3/MK6j4liTf1/pzk9L5XEzBPpcwiuhOxRIT6UsNFF2a317G/s
yiN7SbxEb+YpvBINENPqT6E54Vw3aJCB/36KDDIaF4AbP1oCdWWYkHZf3myCac60f7PU0jzrmxsJ
9ie7LnZd2wOf7toEzf7dp03lr6Uy0FlDOLr9nuyfIBRBHJWkHhA7rpJSrU0UbLtpJdVrUl7+8UeA
WtSdtLY+VvAh/pYoaCiXwaHIvHvahLjV7fkyVRqkwT7pUfOUuXwdXRP+w+GkWCnGxpc4BZedcK6D
jw3yKLLakpY5TfnNOLRivC4NClIgwKh8IYKf+MnFHEP5d2LEq5XIocIbqxTAnyWa2l7s8A1oeDmg
qlqZYgb6wq7D7VXJKkCTrCH6v8Yxyj3b956pYUEgTHI6Rk6IwSPXQz+6W0dmVBVi8cSTIH/a+Vjg
CJjurzwuTCFWeM0nG/S6QFVYP3itfpC/vkrVVTu4vFqYnxZDHQDZ2JXf6F6JCbvkcKjU20jrA52+
9IfHrQWkyYJqhr3s2Wu1pMXfjhjmx3TRX8KxMaXOzEwwhn4+Ydky8BXqRJ95Mrhq/AL9SzudvtDh
vruwBa5Q/+XgohYHQkD1izx2EZLoYi3bzbtyFl8PT293nBFgIaLbYIeMrHrir7TDUR7tfILVUEDJ
4JFz1u4wH5N9MmYLdzraozJNFQz0UZEx6srLIE/VRS9xU09nTdYMWDriGNNIJIMXexo7Q3H9dDMI
H/YPDQQINhHNUWxmc8MAZXjPdZeRWZ0707mtLdFi1DcHe3d91WxH+PPopoP7R6Xp7tGhRuilU5oq
hiOUaAd68bRZijzUzNJ01AGjl1ujR3q4GsTuIST2dcERlnrSig/tPci61mS+FXCWDEE7HfKv0Mc+
4gwV1t0KzbadEh+zB40HBCSB0Ms96Cwkm863I9nS12gGSycYK1NbS1DPFw5In2AmEy7xbREH3eFh
Jn4EbTPTWt6X+8s0W2h6rzgSuQ+rM8Mjru1kYMQI22QNiUhgB0hrTK3LtyS+g1vjCXHu1HeHobLa
seg/W2hR/FjyEnZN9joZpM/3guag8hj8Ym/27LtVuejAxSUlXaOdgBtB+upurhEbbz+4jtNhOuhw
4OLnUmDoB2nS3dpkR2JoiJdn9j3Jpd9ObMXVZLxsN3RhPLta8hxydF90kLebwkEDMZGlYyuDF/1u
4KiqaQgDN5VrvIdTU3PJRb2dxDmmj/8kle09O36rlxDGtaYrvgzZ3tCEId7qL5DkI8DDfhbwYG5O
eUSEjnM9p+9MlqKwWxktvtVhlcA9REyBSD5axpf21/HDBxoPApVec6EjFpJIhU03o6/VmJwWR7no
0KasKbQ+1px6P7Aqp44q2q62/J06p2JOlOozSbW0fBBZm/VLNwQgwfPZlkX7V9UXsfysPrc5BLrI
buSUlCKP7vzZ8o74YFE/ha/YY2G5FgZ++fYzXtsElVoMDKG5f/zKyuVs5RFXDXydlldx4EAGPsvi
joaTV1EfjQVCKn9PVaOzBL96GIQF0zvSkt7HUe9xUCHdCUfGrFCc4iw66dmL6nbcdo79Hv6GXIiG
ycj6PwpMJtsfQcsIqYeUL0ncxIX+MF/D6UL/3spLl+kdWRvEI22Swi6Rn3w4RLgWsLHy0eiShY60
WkOmjNgmZNB+9Te+ok+9o9u2PbEI/8IiTZAptrwVWAVA3CAU/aA5AXGvswx8iSLLmIZTOMmUMs4n
ciuP0KjVupxF73r4AbETM34U4aqlGRq+vSuqBZJzO+hRTsbPRRiTWmEBJ8KkuW9g1P9uvMtoXqnm
T0IdX7FkB7oeXe+c6Rb0FmbqweO+C6bx3gGEUXl+Phir/HV4BXpouKyP1r/oNAB1ZfsRRMA7XKmT
DMYNTXbHSzfPAAetcU8wL9yWWJu62Usq+NCAKjSZ1CIqyU6MiCWXDGdoRk5DAkalZaxgfMNLa7AE
Sk8UEppbEQNJ0R1OvLUfU7+W/UeZtkmdZ80uud2jD91Vbl0fmzkAs9taMfIfNEzpa89UGbwWuhVS
xRSxRSgVwKMv61Pp6aLkdr+rmT+s7M41UCuLxwHMQgVXvb9FziQPx10hmMvhCu7m5onP/ELSRJdT
VdbyGgnzqyumaY11I4nVGVAUodjG/C6Fdf9JYJ6LIEI3cBWR0tLZ3XQ9m6/fMBayBEGhhcl8VLMF
GTVjppeMXb5VFq4Z+I95P8QZgdwbizD/4i+F5SVVxFP2TuMaoQsftcxGvvwMs9QjGhd87vzJSZbZ
pawLlc04tZWDI2KAigVXduYV4YqzdnC/abJvXtuQ0+HNHyXZsb+V6PXywpkjIKCVY/yicjy7ODEk
dbBPPTzRtdFPw4lpbBsaGP6Wz3xrVY9xjScTsKdKQHFDAL6tocAexSJMk7PlibZUeeaepsog2hia
l2iF8rlkG7jMh5xB3bE5Asrj/lLlkooFBu71oEP+Es4X/o7BlXqj6x4qYcJarggRX87RvX35P4IZ
AKr3UUvKRD3c5gbVcu186kmsgFxlDjGVhSEqYUQSz2BA33yIAjMHDu/XIBrv6uehZxMex5fpCR/f
1lvwYeG3TUIMKiS5hs3f7O9/MejpAVemQ7S49qSGr7col+DVGh7gyYDvl/wi3bntoSxr1qpX37ht
BvC8FS5ke9ZPaNqTdA3ctZUMKpbxlhxUGK6SUZ4zhJrH/qm1i8KApsTlaD3Ci2YKpOUM4LHDcSZ9
klPngwTj3q9RIE0dQlR9N12wzd7ctu66R5gw5KNmjqPDAm4lOZJDSrWy4w8aBDBZxrgk752oP6Jz
sFQQd4HRo3WIo5CDV47nG83fvIgXc9nW9UzOruDx7R4LYdW1aPt3KODw2btF0+c+n1nWnVFdpNem
sFRbWTWCG/S7IflHjJ+qh4XsST5YJOBmTnL9MPxHXzn+QDk6Z35obzyOW4GavwKRAeUbBuQC7hIh
9l+i31HV2w8GoK9LJCn13GS0ykYllHwRZZLz5L3dVKvId6t3vQSgghVu9LYiPqQyAbbagR/GUAid
mS8msizAHNcS2xbf7zU+RKhA6Cqd3j663XD3//EVuHjD6kCQkq17E4248awIKLV3d0YTdHy8CBFy
hu2xOox3LESW7dnuVLW2JRTCqIsf11+cSE/dIfxNZIwF24Q3+GrCSqvJje/nOl8XVBPt4ZL+eJOy
BdTq/n0TGIH4qpoPwyi4fGFnC95mzbU96NePuKkgtgzJ24fL1tqWUIjxLSlEhtfJV/a1wmyRHvRw
RBmbRj4c7kLhTm4tcXHNeJBLFNVlTaYrapL9D7R66SThehXYdyhp3zSIxAiFq8N+k689BLdMOU2v
4jWou908Nm99IPpjrNHDcOzhwECU5QU9/Phf+1wgxYK9buAvejolro7C4PBj3KDhFIruZ0uwgAv+
nRq7LRRuIW85m3sjDBkH49vG0vga/J2I4qy/A3GSQB8xP2vpfYv6xWv81rOMQoMxjIdpvhrBx+9d
nVqj/1DUPG8j3QEwGo22W+HiPUjqIx2pB2eIf387lIb4018y4TkiscIi1MKVLup8BkH1mz733Xy3
K04zUTdTmivNI1uTS0Tq0zKr60eedT8c+ABIxRGuzvV1WxTV8G1oYYW3DBDNORdSX9MdJ0sxv35k
SOwwNmL5ssYOiFRGbuvQSjok8QnrYuJBO6iRwM9j3OcS0QXcIjDnHqnWCYAz4T1DWQlA4H+zrQ4i
VdOWH4amq1ehS2TUmS3g/hohdW0E3dRyxoKypLGvSe+X2UkFUytlooKpWCo7VQzMngz9yQzSbJH5
kF3bybjATEMK4MPGf3Sp29YJviTNQR1kXTCJlR8RarKhZ1u4cza1naFbJXOwJbc16ckpL9m4yOlL
TVQQXXia8wFGydUARtPOYEhZ+l0DXBeTsLowc/BHWRYnMZqdtHZy+12xzMSYqF1U7Anbv7ieQC8R
MHQzfCHrWjVyFXBvHRIqMfkCUZKVbOp9syw9Xabn1nYMT0kQ1sZPzClrOglG082m2oEkCjj5SLSh
bu3mjQm7/YGX8MQ+mSaE8NV9us6NzMUj/RzNwKaTLQv0E0Dv6QjqVcTPnd3g29rcc+2GBAbnt7er
JRNQNkHEuS22s2225DPIFGGhRxFMWdknpFgt5YfNECA6rg1m9ttrEkDPxXHt0t+B/GoLb68RiYUy
MNowj05fwjY6JJBGJf8JWOeeyMXYPsqgXaVWmvbqZ+mAx/sDIRW4oIjJSH4uvpmCQFnOj+IeAk5B
WFsCOmBzF+NzgggxPj/DmJhN6BK0Stazkm9E2Y1s96ctdb0gTP9bVrENpdQfoIIvRWn46YbxVjsB
hxwPZvWf4Fha5tLYmG7y+aE1PleFJMvkYZU2HjX4euTWJzTn0AGY77UgTszFvrHctuzjeC2xjeN+
0qqMEFKnjUTCu00skHiVBNCPvtvAmCR8qKeysF62/mXGQbXs4MxrBec+CglTUil4YVl0BzejuCSS
oB8PsnLZO7vkCn4tAVJb96prix2pm6rFsnGOqMb3fv0ZPiufbd3rT5w+yFeC+E1bof+RObYZVf99
T+tWZimJpFPRLm07TqF3weANaD4xxUdua9BkhIT3vCNMdnzI6ESw318ffMclIgBrLMGaluYa/OTO
RJvMIrF1MsLqbCbDMetqLsi28qhXBZXB0JbEaNZYluHv6dJLajM/IeUBDJhVCxLRdSjSCw659+Rg
JyrawvpHt/1QcWjyw4OUAvt9YvCu9yBmpd+d5+Q5flrf6pQO75lGTegQctfRbJXW7SsJWg1uOrhx
NZjirxeYu0bxddN+hPl0KRNBQSiAGjumqrLCbH1DtIVhEKa+INUt7rPLefqo8iOh0LZoZd2GncH0
9o4SEgaE0KT98CWy2sNd87hFtQWkvqH3rjMa27ociZJBUqaacjZLYOZLzdtQGn4YNEjBaU9eEQc4
6pfs9kHLFnGv55ynnWaR4QvjoYWxjGcEhtxEd8XDYIYsve6ZsiMs3+C6MFC73ExTjnYiQKsV1MYP
MtKYUwcLcPLcSC/oUETJu/oIEsVsGOon2/rxmZ/sdyk05k0nace8mX7HlcUnJoVUgkgdXCnkcCrT
wMqSR+e4ebBvBy088gds1WYX47c0xLcZwOZU8R3RoHencRvRAFZUOLKUqj8vvgzUomQfR0+zPYc1
bm9nTCP4dEmsbBpGYfopCFZHzuBtBxnqetBBPhvafpSGSdYRBPkW9pnvQFtbGBAvdaEZNAmw9JPm
FiO8lkBleGucOKMVozvNWNMtCI3lqbTNVKVVGn9LX4IdKH5jGgzCAZz04hTUVdT5x+dZ7bEYhSCX
L3YdohJyY3FTcE3u6xvAE2fBvUyCymcOL7hcUE7StZknzuRCB00xTXnZsIHv63vaLPv8Biq9HGU1
w0Jp/wFC7NHKRAPd+Hk+esGHHv+0N6mXUGZjvBliNTz7qvwzKx0pKts9kgw4ESHrugu5Vc8I4zhx
LFGvqXZmst9cncm25+cQ73afuZDmoNauO4lBchKm7t9cSOOZ8XVnRvGKTXrjVy8DO+85ytHqS/24
4PJyaQV+fouTFHm/tGcKo5kEVxa9QCO6MtbyV05thcTFz3tGGI0iUDvyKYCi0sinNrZ0a31S4gRn
AhMvKNWU1RrxQr3jaoFv4RITeKrZjJqVYMMGeXF4toHHWgZrEdP+uWYl6hKxNiIyJqI+22soCQoT
ChNUZHTy7IcVoxWVZ/mXARnv3OC9w9FynQvAuwHwuzZkkd1+Or0bopVGTsvpbvX162irSuJ+OpIt
ysezNpdFbIYja+5qfMnTJCPZoVyjMOnlfulEGdYIieqF8ouiE2nxAEjBp/Ea0x1Wz7Kt0ilK337R
jOlbZ2/necYKUU3uUjRwWpR8H7ENTTZwELa6EoDLgmHra/mxfV4P4szFz68gIRNCGemAxNOIKJdg
6GepQVvBgqeen/L2Mfn9jy3AiySuuhDAjRwuG9ZHugRkPHQtulrQKIXd7Yf6chkZdWXQ9YVy875V
jgtS5k0Bn0gWcgMzeeYYfzqix47DASeCGvimG39Y/NSZ9aRDf0UP3AthmvGoHk9of1Pd/QvUopgk
Zid9yQEQH3UjEi5Ue0rDR7nuLH2IaHTj0vW4F8pyUFXZtTSG8Ih47pVnqJ7Z8FbwUTbBLqBcAvYJ
YYoVRrhDFTcvHRAABWx8Pu9WgMkHoCxjVpp6i+tfucqzU/GhxCWE0hqhsVSo8QJvxXJII2w09Fyu
WhLpw7Kd52JF6O53M7MObDN1RNssP72pdIly1cRwKN0pTGmzc4aTXdM4auoBgZ4VEUoFQ4Cv/yJ4
BS0OclFtxsi6UyTuGQhBt7oKw8dWJCWd8JFlXxIn+EeisItuGjMBzTvq9/5XiRtltC7wVmIT0J+X
tMRjCzjuMSGuyMOXH/stv2jq8Q7ZM8FRU9wjhtB2tRJANUyxGO9ahcCDfoTyUNker49CXjL+1HMe
W4b9/2qzUfZtF/Qg2cayJe4Lvbilq+2G3/DtFo2H1KKa3VFl2iCywFJo1FFxiz3wQGsfVDo6JPUl
5tEwP/w5DFy5QLHVNsVOLagBRaulpUZksq+af9dXUwsJomWlCMsMDDnBBeQYIiC7JHX6yPDHtvxr
1BXIc+LJIBMi7Tu+fiEthLzLXp13LqU9AwWo6uZzifCv+iFvWeaLT5rEgZu0C3+yGoG8S1wvk+NH
UxgH8F5AmXyTmQt3+izglrSbRWT1uz63b/KLRyhT+0YhMt7E2wxwyGB7cahBPx8gzaiC4Kzu/Ma7
Y+dpu0IoesUNcOjhMCzyGpC7QsKcvJ3V8BgMgbwYCM1t7cgAQ8EZFlMKVxiBJcZJlQvwL3uDqXga
EjfcSQs9uDi/pH64p/WLINNJqIbVngspo6fvRfIg1U1LjwMUHMqRtGrAbMlQU8K1UcogtntoUn5w
lgXsbxdtpR2NlVxWvO2v9F0iTFPiY9gMFQCTRk9TMTTOPAtLSVPe7BsqDKn28lxMyNy6uxOTaVb0
RtISzdGL1qhQnKNwvVsyMD2X8seo+fHi3AJfF0MVXhx1wJic0MrOMl2GWQCmcPg6MQdMmPwipbDY
B0P2J9vKbk5Eo5UyPKT6HQDRR7BHq8xS52BB6BSVr5smgm0pIgeTLQuPN04wv+11uP41jN6rG9+f
jlPubiYeoQZMA1mO8S/zLSRIHH2QxNjgWWmletrP4XiQ9a5bTBY+3XfF8GBsIMMzPuPJFjD9g0El
cBpN02pF92OpCl0/l3SBlk2Wcd45FW6+H6vwtf9pVez1NlIyuEcwUErW1MLpQcJ9Y+KuE2Sp5DRc
IVYLZzxg/fCGO+y49M+0AqT1pixw1RlWph0+PSdg2iMPW13KhbAkdiPp1k4o7iX24uq3jmMnR8iJ
utz7vmmUPsfTl9Vmd5zx9KqGwTBFn8ktMMEbVxhtDqnE6UQe+TBGoRSRmfig1LhZYTAj320KgRhh
Ti6I4KTU/w7tMxyofMpOzMMoU118AT51KtGhuVZfg3mQpICjXGE54hZRLUdNdsZmQ2vCe2+qvi4/
ikRNaDoD8cfqGhqqG04mgdXRO84CSQMGf6TaGENx29WxjylVjfIEjk6BzVccEt96i9SkupkfAJgi
wtUgkGp0S8WTnBW+qiGf7P4oEV+WYrrqScOfwmmaCn+V4+U4qLD7B9IEVhsHj3b7We6tR1/n4w3R
9Fq2bn2DYIfCU/MkR/nSaBzTKZzWzDkD30Rc6713HxPvaNU3cSCYKvmIRGsp/yOTQXUqzETuUtXN
ThYw2plyLqqk02KK0gPAfTNQIFMEhLKfuVGwryLyWYMcEpHzruSU6bETCh4XL6Uly07rCETYMsXF
eh/wt8SgYoTtAE5J+spxHzP06jrtO03GS52CDeftR90KTEy+UboMOR2/pEYttAIijRLzN8SSWhOC
290otufCNxwX7SI9aFtseq1qYgcXGQw56RBbRgjAad6rf+wPpYOD4f1GlX+9Drb0KyUmrZL4neCf
EAiGYILpBZ6X7S9wE8TpTFySDaPp6mJuzlg9c7L7Vz0gATgN9V9u4i2qUqLwzkgHOllvglT4+J6L
CCYsz77bNuSPX+MLQWWgGL8/z1y5MHYq+q8czQEX+W7t/Uu+gcGL/ripZVoIg6sYesNQN4iiHfrq
NVwrgIfbS8XPaCpxxPBSts9inl6USL0qOtVRJXW4qxbChZQ1sGRDEpkZXIMBicXXnzbPluJlW6WB
J0PEvgcuwcjas0+9ionFMRDmhvAiUvKQsIWKeOrX+Jc5OPYrOMSOK6wuxd7CoiOr8gfC8SL0uYDI
fr7qSZ2IFYc5PT4WKlAEmAqIt8Gmy/vN1a7u00Io6nZpW2+pcNA0sQVqh8h9XZ+0+D2XQOSk99pw
1D3wTGQFemnLRCqG76mkwyiOADfs2bZyj/I9Y85SdEFgQd+oPkULA96I1vcP7KsuYY2TaX1IRAJX
DjH99HIaVT/4t382NXBOIEkVW4aBHYtm0riJ9I6jd0ppkmHCu3TbAIgYNLeJZ6nL78KAoSeljoTz
BQbnxWmUcvNaPGwbJfQROD7iytFTtkR28JWwZnOTj0ho0Ez8Z+u3bCR0ku155QhEDAtI8CFdFHG+
+qbJoR8sggI6DO4euVcHrTz9WX+i1xc1D/ZFJczyFSsLExBUBN2BBu3QfsfuC+gs4gepZJQf9wXs
OfRCBL+ps3kel3CBzKzk/KOsShAz/9Jn+arLdItF2Y4ASzxyMUCh3Vr6K9RhTlVJk4Ff64WOsD+k
NBWw2dbvwPHs1NdWEaKeWIsgD7123RXZ9eT8td72r7gkiyWj/XgS2PHFyLvtJT9R7E4iopOnOq16
pFfSlY5AAG+TawnrL2z3geTaN+EVtILWZXsmNPaTGcu4yhHnRRl7an5h/p6xOfEhWBpuoPgH1S1V
zyd3B1j+Ue+tomvE8hLpudiASZGnKOah2vjCnuVS9MJKb8QoVj7Obb0F5VV0d5B7RjikGpSNGfS+
kKwP3wd66gSlDcyD1ZIW4mykBCzrvVNAPqYRbwCY5VF28YyOvN0QXLlZ1n1j6Pmp65+N6l8FIN+D
W5VkPLMjdrNKoM06JiaWY91CuaE8dZ5Z7Ai5N31oicY7juHq8NY57IbhjP/Z1oF7LGyrnc65hUuq
QdDRU3Jc+h9t0ELs5oeZeiPnXjI6c0vl+owVUjH3aVQLniKR6mBa2XCfPyPtRq3SoOcHKAfWfJtg
l5xqQvujG2jvRmzQvqgi3H861LNm50sDLtRfNH/S2XyCHbQlF2SSLOKyzGiLTQGVj8PX6tt9ToKn
5j+BqBd1seMFVyNkQI3O0wY5awavxplwoSbVXPsS8sPtRuNNFWZXomeHVIrKF+FGS6fJiwIQUIQn
Af4x5Yueq1DOvQMedNxgv1dZhi5zA8J5+09IwGMJ6n5M3sWF/EaIv0l85xUaHvp0YWriTAC0m0XF
2QiYdYzIiBmiEJOIW5HhXWmX309DAZF4/eri23+rd+T6BSr39CW9d2HlL25VGNN6dmsmg4dNTPbZ
FkvQhCdXDBlC+pym0Fqyud2fiRcAU+/n8F81b9TPYf3B1boG8lqgLKHnvSJOaItw10X6vHO2f2lW
vDvSewh9tdTnLg7bS9+vh87VuTDVUia15mOm5NrfxIP1B3nPYSE8xQ00RjLlt+lLdPaNhZFg71km
GV4nfhpKJBJePZGq9LSjqEBg4+CNPcFuAsluL84nQPCZ1Bdeov363iJMO1Qkm0eIub6nVIlzjWe+
sNanB55HCgaQ7i+gM5jOhZmYlSgM5PpGLMnocbgIX6vJqrDhQsLPqKYb5XdPlb/FbOCUufwQb7Ow
KOXgbWUi7R5LhQLlGdNZ/6xLxIR26273783W151EUwK3YkmHWJ2saRb1Ij/Vf6MycEzuoAdo9P8+
WYX0WwoCLKNVM5nGNEfhJxaFRw8itWh2rNWIubXDXuxsAnqh7wjA5RGZx4AWvoMj88wn5k7J7hv7
z0rPUOUSNa66bIfJWQ5klUrJjp/oWDs+aatBmjJ7oEiZlZuKBTk8NKEIAxsT6h+2q9Cx9jVGcEFi
T2w5KUE9W/oT+d0P18r9L6a/nwUF8cqekg3vdE7sFilueKhFoPvSZZP0rhG3y0oJhNSmz8JIpYta
w7gLKBpaBH9Q9bQzzYGt14kOUSFcnRnIAGFC9QqV6cXXMMH6BoHDANIljc5ftNLZNlMnuu5Rtb9l
uDTyR9EnZwRTZwCrGRZKVdW2gND3lQoSJO2LluiOtrJhHqcRgdGWzktpUUcnkQ66DDww5iqavla5
NrNdWgU9mRfblng40sAvKJQ698M2Q3nT5aQsHH+KLxhtDN5ioMe0WVzA2M7tryPs2DOX/cbMGKrs
IGO+jVDyZ5zSXje7bKLW5Czxev9uKkgYFocoIRH0mbbym4VIluyDE2WDXBt2Loc2GdOG1WPirUp+
trVTYHa/LLc9PTIrW0UgT4YL280E4VkIV2XKpc5K/KyTQ4jvFyQxf1grjAAIPN70iqzbWjHtV4eA
TD2/w1HF4JptK7m7PkOU/ky5iLr/DW6tclWIrygbUS2xeYOdeQf/EYrnKDawSxw0eaH0WJxJMKTG
z/qHKh5L6lQBMStLctnhfqfF41z9Bs+QMM3H+rRGbrnLeCnwNq9kwGyQBcgcRNCLOsymcECjNbxA
neQKtcrbsfSlVQleWVNmwIL5TJCd8v5POo3gPtppy1LdrR3qC5HmgH7hdb8iliqElyfKnoqBkucg
l7+hc7kuGFKchV+W1wLOBriazN3HrCj4E17V/HMPhguszUXbdiSIRoCfyk37r4x8tcEMzT58rhMC
xM1u+qWcTJ59nhfZKu//0lPLV1jACirukb5+QtrbTwfqFhmnfaOit3DOQPwShAs+kgSg2ibfqzWN
s7GI/6UYRa/cpCGJwRWyam3TfDHK+JNCGLfJFvxQNtBmXAQr3kwZSeQ8guAUwjQzDV0QXTg70OOS
wH1PBbPpbw18IMp19+wEStxM4mhpaYmFUC9TQfscYRNRx9zot1pEIUWg2Rz79kIR80NgO0eMqa7V
OOw6VqBbIvz5DTuAstKxqnhm1l3XAE/lWj8glEvcYT0hoHZ1u3tM+5iTQwQrzuozC8gVzz2Th1kg
MPdBnCPJDbyHbPFjuWl9rDP+KNXTQ/1xQ2CL86LyDwgouJvAjIOoBheSlDaOTmFm2z8P0b4/gVIC
aPOvIyMutqZRnPcUuGWVSDJF4WzUrRNwNbpJmAHYkw32QsqsL7cTZqqdjuumK7bQkE9aA8xKUp9t
zURevlkJQnFQ/ElDGo6Mau+OiMxyOaOYy0RJpsoiYNT6WCOT2Hj9ypZltbzNv9Qf1n+xIYbhijOs
mLRHXC4ZbgpQC5XhWDi5RtZEVw2k+etkspOpKRwW2aHPpmRU4mrb3HsXQlkjdrYhx6x+fxKqSoO7
BC4WWaaLv9uOtwIYwS3snOeJqXW+rLCG1frFsY5hgVcS6PBwkCeOFFWDZe8QOutEiFyCwN9IXMHB
z8HltFTTJx5W/p71EwGQCvWNhyaNrmv2tbm5TeGNtPQwF5pxoNZuAozdTbXCfedofA3RDorEqbLL
QdBlU2pXQMfgXsACr8J/oDt8+6C52tz609BVbpBzAQM2nvZKUQgRHpD5L7TAWRlRgtQ6pG5xrWsD
MfNjN/hfCCq2EMbYUltGWLpx7Qa9bs6wjSkCSzt6tQw1th4XidCJHDbCyLxkyroE2Fyi99jBjz2X
sl6Y3lBmnsuRbMeiVe/zftWnaffaU/ZIPq2wnXRQUBg3RQd1fALHPZv+yGpMCst/GsxAkyeInKXq
B4HutPFJQbyyo7du0RXDWLkk+y/Dzc3NX+oYn9C0Ruy/5rsOKEuLHBoDyQjSsM7p6vjM5X/XMGwK
UjqpMKFZlVtK8HNC/wD4G3dmO9DF4l+HZGsJCyzic211M7sTTIl0G7nUVOl0j4AZodF8WiRyKnyJ
GvM6Jb7TPUMXGkNQZRytTTlOKRJIZsvkRxsowoEa9C4p+QtvBchk9Qeu8AEt+HC37yIWNlaSMg+Q
eFqn1EpxoMdKmOanWx75vB1D1YQZmsBpKcXAZPbi6AYiIRg9O/lmaYagpvDGR+sAq5sibq4xsMon
h1fGIe2u8Oox+2yP0VbYWcGV6B8z1heABNXnZAjmrI3MKC7bHhQXWs0kNLw5NXtXsOUcc4bAQSkv
YFPB8PyDTvLRlQ4mINKpp8nz6KAC5pk6JTQatDKClCVevRZTArMjkUX0O1QjXnvGEVrHYcYtmU6Q
Dib68jGdfZNpu6y/UiIHl47vI9VbzMV+p/EEHhHIT0xz7P/g6TzJb+7wlRjiyaWzOgMF3QmFms33
aukj519XZQroVcaKnuSgZ26sie0JtCTUlyPHGGa+rVoLNTn5e3F7hIcDWZxAcWuelKaADUeMGIXp
jJzuTOpQ9V3Ke1Vx86HuDbo4l3da9Tlz+LqYyhox8RAbP6TplZuz/VReAIFKaQmQbTxZN79G3Ukc
5650abZMiFOeKmq5YSRnhrndPtOROcbWSfX1qWWvCJBGZLwXK1CBMwP/Y9xD9a42s7qGclKEj9aZ
i+58fchbvWtoqMO96Ygfpwb6i8stQ7yw/IZntiBMKYvL5qYRzo92dnftisldQ+Kh9Nl1s1od65SI
VzY86ZfKdx7e3OL8G/Wsvk0xlNsxujLu+DR6KI34EysDJ+ZJyQ+7sqFjjmgsE9brKk75NFJMq/aQ
D3QNdcKJfeD4DUpdRo55zkI/kRzJ9XGuFVkNeQBuRNwQPdXImvRyVj3CIQDWM/rI0nh6eibhdAsA
V8mIlcBvXF7q1+WdvEnIK+x3AcN0KkbEne9wqmbciuNwgNQS2xBg3ldkv9Pl/JNYTSbJ3zUuSDVN
npB29f9pKNzo27EuCK3Dgld/5eiZ1d7HunOYKnVEdmYd2BJA88Y8lLCHsYeKircerBarYl1mHZXz
3ObKWDUMrtteXUNUyjiiQJNQ1selOXDDlpd0x4cd8o0+mvFEqfXlpxUjUkm6jZPreRuc/KOtI1O8
YuNt5Oa4qhEFcPKhtMjwOMmp9pZM+KAOlosSuxQI8IDMMgt7/NZd8suPehIBWCiNRhU0f3W49Wkd
t9TgyvznPIK0Bk1TdE8xv5JYvjQgTa/YO/adwthtidpQPWtsA6GcZ042dCUe4HRqWGqFdEyPpojU
ZiYFjiEuYgqvpXzibVIvDO+lPj0HukGY/f6CFg5dPVZ9vloEVmASjbi8P/ErrGghMcm97Ex6/KuT
XQ2kAs0D9EhdjRM2dpE+nJG3rGnNaCu7wQCmFKc1XTjaVhH9beQaAX7i7+ppBeMhWAEPQlCqCvG8
xaofaKrEOFPNuaqIHZ8APvfb9gAMtydn3UE+K1aZGrxzoyaEqn0QQzSUWfHl64X+KFMyu7PIwzOh
ymbKUy1VeRlOW6sA6RVHlnbmXcWgpEC7MQKwokBtboRtcK6IaxDWiLyKGQzTpNeNqLqwvqkKhbbC
mhSbu2jV/TNUNxtD960uMHGL1mdwdphNVE2b9j5n9WJA7dqyoMKfJSGorbkylw1veYOCRgc437nh
aycMCEfBlDAPVP8hqsm/tOB5Kb3TVLQb1KczKE8as4XQLE2i635bNX6v2AlX86YCJySmGh+ZWu33
JKcP52ZMmmCDwifaRmGU4tZZwZyOpzqFHxRfLn5wYdT6fI4fFQnRRJbhsa6PJeNB/0Wn6pciFfax
3I7+s5avp8zCUYc3Jpc4cXh+dIyfIkd1B8WIf3+B4KXZXiXFrj7Y9xExrSJP7qTLVzDH14QbQS5l
S0d+9i3SHBdpUaepg79Linko6F/BQvCcj5P56j9kw5eWjfTJ7H3P77dHnaOQmMQoUy3/bNLaLTAB
54kuQ20ns6nXQEl3b98bvqGNGugkkalbpLIDWruoqPAXa0reR17DjktmBTI0MYabj4fle14590Pe
tnRISUMwpRg+lRVtAM4wpdSXK1otAyvPU64RO3RPilUtIOFzNdz+BGw06URrVJSzLIhb6T9HujgD
tjizhlZ9i3PvpAhG7SDSMpedMHkM1CuUzT9rw8laYzc4w+CyicpAQSh7qJE1LsP+P/msRPXYuZJ8
rdqyodgeVlmc7QBlrzHgBJCSWtZw+2d1HdyyvtrMtbMCVk3Byh4wHQesyCPzLeTBXdF+YZR50NOK
M/JhSbBKPinp6kRU8o6Im2Xe+XY0579/p17UC/kWbsuXIXtiBbNe3sbeyfOgTRn5xnZsfWPhnmsx
zkjM183GBctAraNf69ofQdYGSZavWoWPyT21BYMxHi32DdFuddjUC2Xu37DsKCv9QkHGRSgq/oPz
PnfInCwpc2JUxG31G15DRaEzsEYMFRiWzm9hFz78v/gGjHz2GVcOIkITrvnyFFx0KEOnYPSf2iqD
HSQoh0b4R8wgxGaHtXLxuGwfY2Ouq82BDsBume+npIs0v/Dl5jipVQ4Y8FsZ8jA8ufXrCCuf8IoH
4b5llwZNv2Y5kEGqxEeeo29absWYyrLVrybpCMjebMZdWzYz2ne/b3eqgeD4Y7ITz9khwlScU/04
z+pSJnL7MK0MNJRmlaO2N84c+Jhg2KlyJ2hTqYOZhZiNRBTOOLe4gObxkhi55HlrNZSDBjP7Cr+6
MdPy0TSVIhtx3lAhAsQX4NKCgyb3dk5WpIt/CecWhMNxyg3xU36GN5rWOJEa/v2nPQEc+njOYw4q
OddQv5G55tAKWl3+tpGtLzymQzKc10L6EW1SkfbKmBGOlqS0SdVvM/9kGXeieRji8Fxjqs4Jdxe6
Q+DhqIo0gj3zQ4wQ1YS0FLPBkXnAoRNYDZR2V5/LHLr8iHbeqVkGSVpgyPfrLU1Q6LX4LEtbXFOb
zz8HdBGYU++XDApa+e0dkBJNkFcMGni3HET5AGk4exmMdcgV1boxkxvBz9qYM98Xyn6LslkEGgk2
CirB4h1QD1bUtTroqryTT4toc3wYNvzpCfeJTAXa2SkMx1KLuhbTuxAqPNYHTNupycx8lFpPId+F
2iryOS2Z9m3ZBdBfq+K2qrBP+lihZSIeSRP7gO1HQkwQQ6tEryPfQEXfB4ifs+MTTOaX2Mcr9+lq
R6Vx6E3banFmTAHJjpb3iG90kUXd4Wsw5RRm01QGwudNiTlOK5M64PoVyEsrG208e0/yK8dTznUZ
oWT+TvSULuqc2QwXXlLOu30V05hAAMGXNsNAGtlZak5DSVbYzgWQVxOsIo0wBI93ypz+TuTB++HH
29/4mBsom+KaTMJPB4oUBsQpc+FpPgY7sF88vXUxnwvYs5xdq5Hayiv4o9bt65F8byxHZgXE087F
yT50H5+CmS/moMdHDw9bX4nywCtzlkMMD0YBzQSlZnqizLMxRKhyzRg3L/85g5rKG439HIuOQ+Em
F2G9ONp2SlmChLIHfH7q02HV67eQzwgHys7dgaKbfvFSjfnAdvFQXC4148INqA1VFxeXPZjTTPVD
Eo982JDMpQwG+RyEyFnK2vtfbo3tNi24tvMRA+FjmjtlqWp3ufSIUdQ++Mo5DiMm5CwTzumIm7l7
ZOi+xahY1x/qiYFWXVmd8owwtkT2ysUzsPkqzARl902dyqo7e241z0+wBRb9S1BrcekDyKlq0RAv
5npK2tKveEdaASUls0s/mhcpvg+hdeiy50nJUfQNO8WCBEiLUKHHD2K9awGDfVaKUqk+LnmvYx2h
tvzZuVt/SDFXuRF06VeYAvyQ+vfgOVEUX7TbwYd5TaLpEGvmOYZ6xeZ57tmniaUQwDOQ+sMIUaar
6dw8k4T7gdlIiRn7kBeH4zQ126e4dYYHkQn+/6GPdQbZB9ZU2ABsxzMovbsjaJ4zK+gi4L0Oty5J
EMXj9nBfxErl/uxIYpyspy8Uj629azMHC5gUIa5QGT0fMR2kRDMkiCaKP6oa4jSx9ePU3KbTj87B
YbZrcoRUnShluJYoB+bD7x+yOO0qsm/Jly2nr5x3e7ZhvNIlZlRjY9ZNZMRNwmnCD4U6S23MHuNs
XugNv4uMu7cQDv3JBlPe2XVuA8tOdz9mCqXKhNXtSi4MytmDksFh16uyGgSOzrGtmwuJhVkDNY+c
fNmhCk78EsZofF0Nou0r+6fWFKNdOWykf98l5MgWRJWq5BtV49XXg2sLLGY9UOwdCr8vUmPbP7ZH
6ijUyGmRtmW78hg6rIwL6lYXLuOWQXeYEeO9hK1sDENjz/NN/JVUYicEVDcuxoAId1II5Y7eIFnF
rWOf6/5L1i57t0tls8lREgrRHd67oppCvnEQ/Ps0gltGWNjyvG6vjxN9nvQIbszHLj6nWZ+G++55
0rPwpyGZilxMMg1rWFFWjMfTvD2vFAICVQWd+epJoI816t2HK70AH2oZ7dS9dRhgWBgSjj+0PHDA
HmHhegor5z26a/+ueYsOtFApeZhzvlINSd+zRUEDVV857knBxNqbjdZAP2Zh47054hxPWF/6E8nP
gYtEsC8sAEJmGjQLAxPyPpncmC0e4rCRm2LZknqROgs7eYIG/XhhIe6u9N24jfwuHkGuhbfaBQFG
vGEhez5pQODo2l00acB5MbCnu5fktp5QhXYstnt2RCVBvqirE+RadlVkRFzpmK+eM0fyHMVBG4I/
seTzC0aUQtswXo+3ccFMfIfEzhfWe0DGEEEAkNAY11n38ry/bjEPZcM8xediCZLsoFCbAqJGFpu9
y28QykjOOCHbguLynxC11mVnXFfdjN4/pvoCeuyptXo/eU6VYfvk2PCC6iLB74BinBZDqzNds77H
IdNfcyf8GoZ4aFrUcITsBKSZ5TA9N9uibOzR9w0Z9I1v9xkueOHoKqzI5IwrvWClcL5iYredL+JC
4i/6xmk9rJVMGyfQPN9uUJ0xmQG7wfEkC2VQf6W0cC4i1HKLseDsuYU7Fk1l96JbLjcR7nFaeMYC
0j0anSXFeykyY+eoD1HxPoQ1vV0bDtRFvGmaPQPBkiwuwY+ptExxI5oMxmGEjVqgoR0ErX5BFB9D
x1BOkrgtyJLWpk4YyPBkBuE6yqVaTOn+aoYAagq2GMXaN2nKjIl9gKm5JTdeNqHEybyf9c//lNbN
f65yPyZgFPj+z7ZpxjnPEidnCw2qwUnFrVq+4hh9/y9k6OhohW0hxVvvwxnJoC95BwE4c1f5oaTw
tRMVKgSqOWzo4itqb2dh3vSbOEoC6nokCJvID4Ppd1OQYftO8RoMXZBBoBbbxGNe8eWdV+yk1tYG
m3FwRPLZn9YaVwQ13SktCLg/QqfhuAaTwLd+6LUOaUF1qTitUB9JmQoU+39+KJY3y72CLv/Fo9G6
LG/iS/94URvkkzLM8MP09bdpyvFM7X3iEiAgBpjgGGPtUZcXh38YetOjtyb6dXKPEA0hKW/+julA
N5EIrbuS7lTqCqP8pOSzYNsiE1MS0PyDApXKWilM2PH0RZxEhzkYXdR/2TJyyqH/V2f2FOqDLenb
BLLhtWlWcCNeWiWILMBF04JX0G2zYWI1Qw4mV0+iBTfnHy6bfhZy5+1jKAwFeSfH0wzxhHL92ytL
VKhdP9pjLPkPjFJtY9Dpv7kspeBuGKLCViKvzvbiYNNgXtg53gKWHvjJDwrDR9cZbz/uzrHdRQQa
36oQH90DuFbpfLOZTtJbrNAJ1aXI3u1NUi9rvFJTa/dCKYeGvpCQsFbrdcbYf1PDw/3PIuRxtqDD
Y2Tz7TrQ34Vb4EAtH83l/ZuNZTlsI23h3MJzBQsBSPbiRy6adVpKlXY3UCvPohePsQDNO6Bz7LBD
Qo+r2v7f9hIhoNWnUQsEnXqpFvMEcjGdaPK81DwlBuORP+0yXZOi8VaIzhdmDcnyk2uPJWtt1xMo
KxOvT3/6ndBOL/McvQu1JP/Kv+sRe7QPrfONONgP7DIOfGDhbPpOOFYN0c+rmSBxBSmXC3BpRTIv
yhnkoxaSsQUXfEczDDHiqN2wW4UTgRN037L3XQZSuH53ybvqS7fmP+Hx+qPJnYD6I9ILvkSC2d2o
fdW1TSBnKntSJwLkqLlbnT27kxvDghgMdGfXY7JoaselE9ZtwsIpY0FFCmwWXqts1FLkiqG1iXiu
HfWPPvUFHWQy3keVMbGrFakYYPAjWx48H+ogY/zEu0taLkzhW63e6ScroMppkRbqdXFGrXGpMOQH
aqWlY0uDkSrvcsVqSLy0C0zlnP9Fw0xJcmbXU8Acw6S70hkkX1Ie0T9sqWyho3LH4nLVukJwvtYc
/AIhxyDeNZzaCVq7jFTNufvC8PiqimlMUh9QjXrYBbe7R7DUM31VmeWKxnIXgCEFJ9aL49q9OhCO
iVo5d5WTE1BTHUJ0U6nr3xx8jVgX/o01WyRNKRImFxJQKyLjVDiGMsz7a0EjgT1oPA6846ahM/7z
u3CWQKO8wUsezb5m+XOQ7xTEnRagbGRHNWw6s5AZst0wHop3TqW61ATQXn9IaJNVRGTQdT/SPf2/
YnrGlRUGAnXBlTrYeuo9kDNVD5/BeD8rkhnekG/IUa2XXbReaGWp4O24v3e8j9mUKAE3eikmuVa4
GYIWzpED3sLdCFIJqioXFFqMBfn4Q65dnPQStdMMkNNfEIUj07MHgbqlLpllTFAUKOzm5aYesHN+
RffutTD7wqFEJYTRfaWA1WF6aN+4iYm1qXjUg1t12bM4KCuliCONAyCiW4dJ1fZ1bb2HWo8H9H/l
pY+RLytlaZRJU/cmWBhCb0yK+Ca1gO9ZsbY5azzreE6fyd225YZTPpR7DSFCCy7+rUgBUe/4mp2K
RjNTfJ7njP38Q1w0vxNaTDpS7N44NKXRAogoC2tULldYsUULtxC/sWLmPI6qv0FfVIRt3z2zi4Ta
6j006q3GEFOTLQt8xi9k3uOSzD//ekr3Vm7zcydfvKQcFzOuSA20pqVeAm7yUXx8hnZwm++ACDvF
L0zzDwrWNb1HznLu40GNiZksp8x77U/2VbOfqU1hjMBrGupV6dCF6A1BvC7A1oL2EhUWjWfjHlz0
JXsh0OWe1e1obbWAv3kYWbZlnxDG6H+Pzjj+JqbYmSps6Q5/lfW5CxnEDWQ+PaK3aaieKhVaLfiL
Qls98jCf7hOPhE4UY1szR7W6NNF4Hu7Qd99zfp8jJMhVva1oB8oh8moFfwfH75mg4eV4IAd7QBY6
1CmIricNP8Wqh7s9mJwX9ECHM2oErBDZF73Zdj80u0HLx560BYiuX2Nf9oTf3j6A2wulMF0wI2Hc
5bbPXGSInW9TF7aXV1rutcPzbMSm9VDFU7D0OnjB2dIbeoIgwkdo+DHYZQ0qzRgROrgajYmYeTMH
OB4N4cCjPplevoBJLNalh8mIdJC7tukPXIfH1nvsNmmllh4ijQ2bh/hcG4a658CSpfK9rhiamiph
LX1MkoYlrZElFGBefPfg0oL+aKY9cZUikcimLFIZlb+IqGy5VfbRXWMXDXDFcrVxThdsLKwmfkem
1xErXxKdzgQqi8wKaJicXGCv4CMhdcmWNpS8cQ6ehBz5G8Anjfq6Cdze627OrhjqSBi+XuPwoIU6
ObdlIULs4+vlx9CykVMMQhaj7S8sDYQ3NZObYI7OcoblD8NBcJxWFG1W7iY1q9myHjLFcM68ZOPC
XOm1fK6jQAeuyo6CnRjpVpZoCjd7+Gq4Vzszjb93EaI/oAh/0CWp/s+vgbZkzYy7VbJ82HnR3/Ni
lOmvFjPWn2hvoe8sI+PIWqvCBZ0wlOMPRM1bK+GrFkyvduTE7hjnoqZ0KS8T6TPG+a3frjz+CrH/
3vuBsAU0c6qnqzHJnNMNooq75HsoNdnXXR2+XgIm8Xx6eLAX8NMa/plaVOcyndYYsHkBGJRvdxQf
BIt4nVW3+4QkjrivAlRZftNu224/BoL1N5dIrIlDweZGttdhjEj7bc4fg/uPjM+wqg/4Qp3aVlPV
fU+Wk/6mZdt30bG2sbESYvX6SFzNNmrmrzOp8RCw9Smu26IdwOet9PLVCY3wJ9VyAbU3roboOWm4
rOeJ2Ix8UKe9/DDepbHO/0gDJoTW3se04/pkbzrjoVF/WH1iEdegqcjBsd1y8LXb9bgC4t0x5dem
d+em7OUO0Vh1wV8Zy8E8nxlseAoGv/o3AtXj9hxAUbjIXXNJWgJ2iudt4ymPcwc3iBAS+BY0JQzL
Wjj59QBt6PABt9UwzrEfzYaCK3R+5lABu8Gd4Ask/h13WB9/EnP/MCVbBZNX7NLUdzMvF0jOPDli
SLK77mPtJJnCb+ZvXet8irpYn7csKcnGR/wvbMFf8CmvR5GcQa6/hnGc4kpSmyk99tz4mMcPMQP9
jJyzwKg1jVRg52i+SprAKijmz2p0fB65xdV+Wu4VQCzgWpoPjgoP4BvsMiJbKp1vKuVuqypqKhmH
u0L9TiF8B4U5z0DlgUsfsbJbj1CgtQxUlntZBiMEKTqNtmzoTIWAZMpVTPtTn2g8GQCWdn/qRk1W
fIn8/9aKSvVfqSMOcj32UFlx6X8LsBQbPvE18KV6fRAma8boBZ/5qE1IhMzdeoiug04NsjQGDMfC
Is5J5wBNHyPc2rQPApD2K+UWjqcXPkOl/Iv1zGDTl9TbbEguxgoqrl5gJ73IDHQiV4W4Me/cG+UU
TgIS6CfvRxhgP4yYUInVKw88u+Ki3Grbu/GPXYp1wRdgfhAFfvWBwppovNiql54lk7r0LkaIAK/+
FzzYfhMNti2t9gGHUQ2s3jCdR+3R2grhEshb9BL71P07CZBgpbvV6DPlY6CG178VkezsT4t7gqCJ
tll7qE1PSRdNIC/KUEjevHK796VG9yAEdUIbnQIOORstp83RnLuqU3QRYPnuejoDsh75QK4gbAB+
oCLFjj2xngdFzyYnPy9304vsQwR1lKj69ewp62uVpibUZ6ZEGpigjUdzeOSz5eUPklNUBwUpDNP1
f4zBOelsJ/REczorsgYscEjzkhXJJ4hQmxS+irZIZjRYtfP0WiDkyr/vqK7uOIBjJZ//DvQMUr2m
Piru5k/UySZR3oLHkNUwey+XEWIqIlAL+5L08NWGkgEUPulHsW8Ezbik/DPjYcdpQBWa24Ut38hG
yD8vaSEZgykmCGYkDZnZU0rrneWHQbNQDrLbqzp1jxRIX9VNjyYBV4xLf4qvcT1zJAVExrMkTquu
O1sl6hpRpIfRG0PGlwyTo6HXYmpdnYmrjeNixz2gstx9PC8T8S9mTOQLsDuDOvvG+yI2BIJBiVyS
KtEi839dBdIC1AbsicJ8GtX/X1tNa11kReainNZAgk5fg5mUz0xfcTDJZ5yqwYUyQEiZLFh2MMsm
2sba4LrrBiQPN82G4RPEuykDc3VakhzZucrokEnnYRZv38Ci5bm1pCCMLFh93seUoRYeGfwgAJs3
WhRSLiXr2SUVqwIb+bggE5U98V9EALHVHMCxCkqG61gBXDV9ViBlAWfkm1avkXmqLROXWXgUzDOU
bQ123dDmW11Q5I9dUs78DypRBpsDgn/lFtqEKji0/QIJNT4FxGG/jtnyuesSg+M+fBsnUwMISHXX
M0XCKV5YzUU8FeWIpsgcmaULFHejZvBK/E/2jdlDYUTUPTEqWPPcBMT7nzJa98OVlzqLMeaG1u+U
OOL5z4NazNGD8rIfYQmVa0pIjH74P4uy/RXtIJHuGLlKR0r2z5L/uTxJUFH8EUzkcpq11h61LsRu
cwke/opBTtx8jBYO/cJymshjasw5sB9Zw2Z/I8Rz5Rbkld2UpEkO+QcPFPF3fRBa08dHkalGJQJI
ZriGCujgFeb5bD7RoH4RWwi4LQqkg0DzK41/CUg6aOB7JXNghEWxNpeUQLqj4akFc/lfJpYORqK9
ZRLvcDzKOTkMuTKXH/1Qnyaf/y9ir7mTkYuXSuGfl/n+/vbYpLm93UDaeTFsgzy4w5Iq9j1Cjkf/
jhdbEiK+pIM+bmDogDHyn9WIJ49LCa9iCAuYFbuRxGU8LOS5WbCsfts73iDaqm+LjR8RN6c0P73d
YfjHShl045yqLPU0YoIuIBWbPj5xGto3Xi59iRRE0fF42fLmtZFb/I6pEvbniAK4V9AqEpT2CRSZ
zu/NcKqgPv/6HAJ693EyJKG1NHBMvsgLYTWM77y0QZGXnVanDgk76R9ihnMU6OejVOyjjnqv6GHX
yNjQMtNijuSxfdrTjQjdl8Szc6UBm4I9Nq+PFdAqW5mEmlxw969TYvb38chh/1D9xlQR8n01LaiN
2tDTLzBv4NTdyyN46cbyv3iBp3Bw+W1FuedSUmpwqO1zoVOvKWVAoLNefNTTWgTL6kgO1Ebj8DJR
BKOMFZL7gyHs2fORUWsgBIh2GDmks6pMkI6NhjSsw88znoxV9AsIMesQ6xab6EgJHz5g1/hGa0xa
zhOs8jcz/x2JhxMz671Wo04V42XXUSDxeVeSp0UtgeGA+CLl7zjtFwtfLg4R0lveNcG17fcU43SJ
k71FEjQmKcpjjv75aE4rBsFoTE4SRNLKr0pG3l+2UaYM0UammNP6Bo0zeo593Sh3WY3PMCsuzTXt
+xIdwVQYA7oPmbIfe/FckjDc6aJQsDimONVzYB1HHPJb+eqWTeBqBoskpdL0+pHLtpeHYggFld5e
kmYrLRByzgcYX14Ub2gixLqOVu4mJsLIJLsB1vFYg+ZG+ZBc9rde2iaLTLzBqhR+wNfsPZOyHU9D
bps8ZYvAT9lloSYNYkqzADDQbpQ8TfpZ/1TM3lCY8efoqWMjWORPBDu2leYosjEN5zyI7hykMA6E
boNclPG1HrV6BS6yLiZ3B++yJ2mfp6jCWwr3SkjQLfsPdW3Cz743ik47Qj5zGMVQP9dv5G7EFCWn
3ybe7XSojBfw2ZhmX0GdKBQ5bl3a8ViyCI6ZP/PuxJAd8VeRMmanZ9UUXB8lDZROC7PvpY8iACgw
bjRrCcVcY932kpLrH4xaOA9Nj4qWImDZzWJVXzlmNs2p0rwxrFTF40b59tfrxGC7I7ynGJwujJkz
D0yHRg1FgJuPd7dnwZ0VfJKC/jXN5knefRKbdrS/6WMqv7Pk7+yTLCQvqWC7dAMfiXzgM14BEnhC
Nd1jQHKDIOBOA3LcoW+7dIrUemTp7IcVvDQu5S8bNLmM8n4OKkRHIvzNWVrKjVHMgowCD1zm4DqW
a9fcT1sW2f1OD2moFTaJ7lQot2AjFjrv6KN1jHV6K5kxUxtUDptkfepO9fjTGB4t44WUPk/mzP0B
DXcLpTwtCYqHuiwEgAfFRJmjRNpmqfiYO8v2hcrGwz9KABLKQZnJWLAxjxLdDlVvIS358WfYRpiW
B8bazCNXGywMgh5/BOvfVo/FmA5YcKT+hG+e4c9CX8mKoCJHFvmqbUkiJ1WN9FnXKfHdkVz0M546
CXdknz/h+KiePEcx6nR8eI7sH9UllFl37jurtxe7RECvdaOXD5y8ADjGW83LS6jN7Be84dTpHLZD
HrbFqmww/5LcgNEs4FT7sUWIvkrKmj2ujQLTF6IrAZAQmj5yBx8HEk3zg8p7uOcwZGk2hCqZ9dB/
LpSh+J3MkbayNBsBhwCFWKdbrdqNtgWxZJ/XWb7fFwD4KIi73PWlHkboVdTBywQK5Ll/LZE5dgIk
GOayHkcuP/9+BeGH3FOr5YLkzv3AwPrCjDcRpGGs0Cnl5olwIM+3n7rT87WH71CvNox0HWwxiqac
/Fub4DuLkirYME0lPT2rGuW1v3JaDU5joOICdFjnaqC/d/0sWImRTfAw/n2fTHzEbRaseLrXAOr+
19khSo71C2wtzKR1B6Qqwk7c/TkyDX2lD018pU7yAIsLM8WSlPdytVUy0MDm07m3vCZ51glNVxeW
9lUVQhYpsnkBkWPS1+DnQvKSIDUfN2R3uuuQq4CuQqTrWqFKl2DEqkmZram7gcvfk4P5WCT+W9A7
UzhOIbB1wewYbxR4kohTSmv7KS71j5gIDUHZ7uJ0tKtEGvHbFou/EVCY4gxnta6/fcSgrmU6CM8k
UZ3UhJf5x1or/IIVbEq89tywgIcVG0llR0CCI0LDICkGvihyHsm+ebEFtCN1abDgWoWLDkAOWsn3
Iu/cbQOh9YPsGpsC5gMTcudhoxYXuRDp4ipY5w3J1XVgFguxPuSrxpd+2gW1EtEV7kwghZTezyqA
EkMiEvWOBZkWk9RW05H8ShS2Nwp087q5Cyf5YOCdTdfjByjW8PCsqNLb3LJ0Gqrur1ATjJ2KujKA
UCeGwedeIXdeZKgAsTbUF8A10VnXxaxUcB8QOEqNCRc+AQ/TT0SDGNsyQhV1R/Am8Q36AOS1vW50
9wsVqmQItYldy/sDaPuLl0PHFzu11ZVTM+fmDr38BQw100ymAK8zS35IERFBG1o+t0k5OZR7sSKW
Dug4wv17TLPH5RC45Udm/Byu58AO4CIIKrRDuL4F34PtL9/swHqDzCkxE3uaYJNKJUtAivXCINBd
cNP+5wOq1yYmPNhR9uM/PAM2qybaUUlrAq48kQr2TXdgJKVEwZI1ajyxj33hbwrCzOhRuF8MFtnw
6OCQtYy2XsGFn3MRWj58nt1vOrQ0yrP2IYtnQPs9CPHcqkNcAbHVD/pvEw5vdFPVE4DLTDiLe0Ri
8WLgHp1vyZCmdwtoSJ5lzRNDjp8aS78WGVF8oHqSCYL+wGa1tOhuHrLmpX1tUD7uNtGbWnqR8aK8
q609MGp13rVbE5R9b7VTME6gfi45xOsjq/X+GuNpMi/jTreqe/hPAj6tWnaAhw4nATB30Qf70KNq
UdOYUnKA09KNurR7mMzmI7slK98jqlW9veGg3t0WXTWbOkaTxQEaf5boUQnTvvMa0CC2RlCIH4Qd
jWvevXlZ0/vopOx3k8ee3Z82lqZMK2PGdQ5VEp9gB24ODxWd36Km5zDAont6HlNLLW4uNim8lbI5
gKFG9fWhMKR2zyXhR9HIHXcXbK6NPjqH2D/TkQRK4lo2s41n8lvhmWTDLNClGwFDmvALAhdCLOH+
YP9j1VlxMN+Hx6MO1cf3+4yQAZzLk8c5ePxJhHNS3PGGRokaOkxiCySUMZG5X2js17K4iJHzqBr8
qCwNNmSmqstFsPE5nCsqhCeLHI7v0hq+avqjS7k7oE0gnMqmkksqrRBNtl58WNU1XGhR+G/p8K6R
Ho0hfMWcNuiujU9nLmY0rZEVCqr86sQAKgcQ9BjMv7r6+GY5WpvP1LZbns+GqBZEAGkLfI88wEF3
PjE7/GfHenqaWQdVjdc4ykU4Qv1JmAjLac5pBZRXl8eX7DQnmRUt68CV5te8e3Re9wWN4TGTjHbC
lYWcPCFnQwY5ws6hWhozvgyCAZiGtqu2KUTiGdDNZgBjGfVbdUB/0iuryf49b5pOBkr7jEshHex/
Rttx33m4xdUcuNoEsRL9dDBKZ35dis6T2YoR0ObIMnvO0CjSaRq46OQ2y6hyAPe9
UL2u
`protect end_protected
