`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dqWL8s0zCsvkYc/RdnpjQyDXYRC8lujJjrHpNSVmtATlwxlOs5Yro0UwCkl4Vq26+qKPWB7TmoHRx2FfYujV9Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EkYzeVdR9Oem7GC/HzcZBK7DGkdeHD3rkVaBiMVCdBei+GlL9pcEs+jRfMrRFVjQe2fgri1rD+N+Vg/GS4/sFcD72PNFSHuWQu4PHWnU5of/LYuG54P/fwuaIQPJbcYCEyIyv/Ycf5d/m6YNV37W8X+jL0JZF/LVWRIvaQ/HQ0c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oX5GRu9/NJZKAZSzddunNoyk7MggDO43bu6CdEFtAOE6yxEDpe0kCoHvQHWlK1pCnaP86+WukiBhD/D+AvjmylMJcI1tJH+4pk6jyjL6ASuo7uoga+6R/L1T2EVAaYJ8lIM4e7Ft4n3ToJKILQhhKn7+nO3AhFCvorN6+ACIBC1Vo7/M9p+KoeShXQf0Z5rqdX2iRsCXtD50RIXC3kA/E9RNlqaRLr3zOfhU9pgSXhjBirLFtTx9lIbD5/qhPlQr9psBRrSvTFzdgLRAXsJ7Cz4h6rX/blkLqXgmws8CCQquzWs9Y0YZvtHZb7sFa7iSjXQb7ZFSVdrJ5dtk5mWP1Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RUSF6VP5U4f5oUDsg+FV3bApHlbehnfBekn5eYstX7rNcJ/VmPbr3XjFCcoiVeTG1DfboJv5bKJt/a4gJOASfPla+YavBwMAvdMRjcHBBAOicbdvv0v9G+Cq9sZBGViHT4+zjIcCqZtNtsp/BPH5hWIgT5IqkAC7wQ4ZT3HUAvE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o0RTekKMcuhesyB1xGOlWP8fTlhWCtcOd6zoUXkPWp+5KLFOKiJ91/Q9AJasEUhjy0Xq+7SOxqXKbzta/4r+bXsfZjvaor51Z3aNhwr7gBlDR7zfqzflo1vLhY80eTjksHIk8s3BClaAscOGTjcBiI2X0JdD6+/dcDiSAOtZyOd3TAY4se9cVLA0pBBVMFg0/JDNisfC67Med15SBrfqbPy47isuLjnxNqckDjWB8Zn0tiyvKUjleZouqtBqtzDTCBjguixSnFMKPP1UqJ/06R1qZSzpa4h+IvxLjAUUwv+rVdK8fvHiiiyqUeCp422ukCl5yZ7iQ+6S1yA+Wf/W/Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 427849)
`protect data_block
7TSF+wNXEg7yFV8LbmjkFzs1Wr7It/H6DffHpjS0hyUYYqLryAiejOvsUzPvRkBEO1o5dkAX5Tdq
bVrMoQW3Il5UgknVBNHDYw9EXDuh55Nv5QZe341IuJ8mbIf5HH0ij1HwFTf2gIbuXGw0o2EG1zs8
pzqY2eBvGNvANfpK98xfV3irbkIEs0EMnvc7SUgocYn3Ni0ZfheECW7VZyikYbonP9OjrxCTGlG7
oVd4xLX1CfOOl974W3Q/lIEgjZPBZThwO8gKmnnoDryLZd8gJF7k7IxbufE4vW5y8kHM++pZ0wZn
htFMWmXRXn79ipyaZxXSCxOBg2z0Po7CTpujQKSwn7IdcvvsnH3UOX74y42mvk0J5O8bB1GUl6BJ
sAVEQonYVzOo9q3ZoTQNynFiTEVPruW6kdUoxbiX5FwvMcSFUTDU9B9xtWo/CKVWJ1Ji7vMPDQ/W
CFvhilpnuL2MPvYcj7rxuNXK8UBsQWXo9cdX2vyzC2yujrxzX09GEDZV+uKtnyegkU9KWAZI7+PZ
n+efqIRTvckkOaOqC9KrNArqgbOmcXT/x/9pce6naDwar+Td58nfbVWIHE9YmclwTlhHc20lQ7Ih
GLvtw9UBj+Y0lYhL8rynlK5CymVhQO6P6W8YG3tq7HjhnKypyP/iMddWAE5UvZ0cMEZZxSu/XKAL
cmWO3jnfJLR7Rk5thq9ZBMZfusQAW+3OY68vdDj1Zkum+EuG2mti+LAFeig/E7aALPJ7U9mESCvc
l5wZk61PXtN0dtvHeGTkETgS+oUeIjTwctc5NWz/oFOk7gazracAntPnJKjvKZQM5wARsbO0t8cO
UOCYMJeIiE/nOrVf0CgS8LnovRQNNI5B6YHe4Wx3jyhVI9dwGy8ugaAyoVWn/RRrsIQBTceFqzxY
aRz7jfihGknU1moqmlBnWpbr8n8dYfWfHoM1bTLGimFCgc1f2KzN5q7fM3+H2xVAxp9WWfl4DoMv
ErB3j+wRpstxZIgE3OzQXNFicAzGRZt2Ef2C3wz7DuYOZ+KJejbw88HCO/vWDBHN0FKkzVT062Og
EvHe5/vbyDYtpxK3np4Wa2ZlGhVGdEtYG6+wIT9lhMXFWt2jD8quGHQykurw4i2GM+2JypmDR4RH
9drsrjKAIIBx7EmhMgdScyjWmmGL+lvZ8eNvXYbpPzAMqAAHVVWrz0ttkCOPdZF4k9dZ1ginmZIt
wW54ySbQg/1U5AndeWDBFani5OhNQ1J718uIj2Dm57Ztn3/WuWqUnh6By/UErIXTJOsuMo2w6g0h
nBABTP5a4NoRuJcy7vPC8Ng34bVixoaoymD9gaT2HZK67rBbnFjVcSZ1X9XhIzy4KB13L/D76NBO
NKl3yWgE6pk5wrtjbfbTylJ0w/+aSr9gu7Aj7UjIHqICjvCxeRKAeLVJkOxnaktGaGelTuA1R6Kn
A4v7MjJHpyqweV+SG0o/wJMdBtTikVkusz6ZMqiv5HBAkwq3IdmWSo07EhRBZPgXOYjEo0GcXhNP
UaCv2j+df4b6e5gwSVlXq/BRF+D/cFrXYorgBFHiZic+RyqoocUXDtjBZxNBaBi7G4jalUDNeczs
Z4a97Vfp+ExCkRAUVeSPwNC94+yI/8Z6gM0mPy76uhuNDZNCVeMsz9CxxUFAUdgOdDMHPIaNn8yw
oervBBfxpbx2A0+5cikTNEH5TN+Zcl9NjXuC0SF/dUux8cLEAt2AKX+fWsIf0ON8Lzq0rfhMkhw9
d7uG/hJZvT6t7OfOrI/OGUELR3dFh+5ZRlJN3+3/oJR8kiquwZx99FwvHfVyCqDUpMhEQO01Y78b
wCUeIkzm9MwCt62kH7HO5bS0ln1bhUGmgs+1/yoD3AxkLicHiN8VxPnoAS78XQhq8/HX7sdrfQMT
JInJiEg0EzETJXMDzkAYhCsG6YoAFm/OidBu2mOsW40zYNpbs+8Fy59PVAmjojLNbo+oKOLIY30o
hUzk528uBhw58tM4IzKfXmtzVKvK8P39XsFBtT4O5cE69oLx3H3io8bcH7AYxbmz6iMv0qiQQjBh
09IujMPZgGQ/yDDalctoithgcBt1QEE1E69kp8wZ/BedRWciqn4Pd8EVbWMKp8KDHabKau+i3U1H
QXGZl/FFTc+quowEBM2mNeMBVzisEWXUy6Kr4EEZuTireruOo0joBpYsiha90nYHW8P+gYlNWX9l
MbJF1YkbL9RLUvBAHP9a8zfnRu8z/rxIGcRXf9El3eXiEbaRLTAxXtBq1Os2IDw1JuMKCo+6KdrU
xDHMFxBd7lTVel7EHbLTSYDAm2Z+jhmHlj1ZKYTgvaTIllq8XJ/1sRUIKNCSfl0kDW6q9HIvTBB+
C5QlFclv5OujS+IA6pk50DENB9TP2hhWkkw8C1R6ANzDeMihtsZNE1Q0UoQHNMOOlKR/wUzwrDTf
qz3dGYQXt8FRufopk+pk74MxLMALnKKBL/M3yNYGYcZGtvsMias+9657JuGK9nFD5oczC0CwhCy+
yQCE0Fj2AkYEgyjHK2hTtbMGIlVF2Q2L/1524D0iy3LMTPvxD3yJouxtvbROGyvnBwkUEdDkxxcr
EYhlvBJUR9Ps8LjcalfdSJq1tDwXEZnB3CtEhEmmcwQO7MT8E6eSQYcNKol0epkaTIKNkp5OEwVD
d6T62PUoB5vTzeGerqRN7HcaQvoKLCiZUZ1n90u43+USEye4omNWULVVKK+y3jsBgvlddTBChh3q
Fo7X3FuXeY/LlIZ3TvOGUsgSP+ykAOOFrTItprKMWiE18PdaRyddqfH/dVZ2b1b9+6pF9LfUBnGw
Bw6FRPwyuL1MeS1g7HduwkStvZ5QwUu7sCSQPigDZ5I7trhOUC1xqajYTpmA7Veyc+6075+bzDZh
OLreEMoSuyVyehoydsY3sxCpM4rZRezt6fRLLnwq4dFQhpNmdLroI2IljATc2FndrocGlIpgX+yB
XaezcVbpDuQJvgqnG4fwnXRKneZ7K4AWkt66eNf6QuWDzkfMbYmfwK7UChUlXcLhPEA0umsQQrYA
WiQ9I5Q5jQh5TwLIkrDNihM4HM/5k7RdMLxdtjOOQGpaLR8WVenLogV6Vlg6RQCeE5yJ72YUhtZJ
Nl1zqSeJx/Mxvq3wcJYl1sunpoTaMZuY/rL4ma1vPghS5jW3nK3sWGHrNAgbGOtsawGIBoOHIgCA
ceYtM7x8kaczDJ5EYmoeLRcE50VpVsiUs88LlW7C5WSvEaS68Hx9GZIa5Wv3v1G2DlyYmCQ05Bb0
48CmvVKR9MT9pQCQIqfTBd/Tyb6q+05fpokqrauHFBWK+NpX2ljdXrUwdhrZT/9rA9r/IupBD0UD
yjacrhlWuBZMOUVSAZgiJVA0HYQJl0FFLPBcWWtIljqXMY0EUfmxX2EkSRampZ5xkIf+pxIFauVu
BcuBbKcTfBjFETvuhvWSimROFel+Q7JktJX79AOYriycfKRBsQ825omET2hL5+ACxfUjOiCzX0Dk
fGUBFMpoa+K9Xw61WA/yN52kATHQlF94I8tj4MXKGEpkcrm/wNyrsXw3KQaXfnPpkG/c95Y/4f4l
GfcAnh+Bk3VMHoxAQt/EOVHFsDvMMV1Q0wWGdwCQCYQZ1YYOalqC/J2Vz+FinKjaZEVgWvk+1r0C
DeTtk78lXXQZ6WoagFHzmUCCzwblaH7VPCyZDNKmSiGTh27bkJdkKTssTIzn5jhBPo59UqXUeie7
TF05kcX7CGEn9UdaJXgW4Di6ldlsHDkVzcF6GA2x/qwt3mifW/Ifxetc7odvLHy+pPP6r/mBPED5
fQIlsKoDQtaLJbBSQjCSGajq4N9PtwG3H5RSjppEJMvRBZ38csVemGtE9eykDk0UURBYXJOpSDHA
HBtKG+CqYTUrTL7cLoT9uWrHsKY31KHqx0YrE5wbd+ljZjYbLAoXlzyzDt/xtPHw/JLak+0fjH9I
QuugB2web/YoUEQfQZ4uE6ki5bW/+lGXgTL2VSk+IaIoMQ3NsnFKj+ffV/YDYaLPqDnqx7FfB7qw
xbe+3ptZCipWImGz+bjyOC9UfHgoAUMCQXzNlReoBivsJdaSwnspUEjV2eylrQVUlBwCjbJozZUZ
1gueQc8AhqyRxVDbBEeHDoHfTVs6xrNTW9UF51fDfJ0wxDBohDvR4QxsD5206MWlJYffvC0GzaIA
BFIM3KO+vLpLbTDkme7Zh4cfMSRvFy7+cJC2fsl3sd5WDSUixVr83h6jZHkiH4H8UUBH6P0Mmfr9
bQ6N86gYgiys3e0RtA7CeAyK7h2wP3hYAfTkVec9LbWqI0tr9akFeXMXMPnXo8suFPSSTkKUGf2L
TjDnU+R3YD/MtqANhtoXAOXLNT9LT1zJ7hQKvmcw9H5Z1qRqQGxQsyFVuQqg2Lns7dFdiFKQDOYn
kvSt6mDwizNUdYUu5EEh9FhhOPxHJBWBXC29N0Jnps/8vZNsxnM1UO+eO+ZtMaXgGu2PRc6Nfg4D
CUmRXaegZv6TCAQ2CWX/VRG7InPdfctdU6Zi5HOr3I/8hxcgcqiYXmQl4YBpRqvgouUoylUmtVMb
CjDBkfrNgJCa10TD9hZu6yGO5PtUwAS1LjAd2xV2H5zngJlWZFPtsee8k11S4Gf4xRv+VZlMcdZy
INegTaj6PxyEQ8cFZ5mdgTA6+L3EhPfpNXnrG1N/leEwisXrbpBa6jSBsNLRRgOgBpwpO16EWh5X
Q/sKw+OMCw88bOb5NylsBp4UPeE3uRb4pM67HhF8W1mHqED224l3FmYdicfMQSOXfBA4kjXH5gOv
HMxfem1PK36Ws5KnJJuo/E04DjqSSVPu5YBuC1T+Jz3Rc4dAeyBKeDpUp8+0iAe8X/DCqa/x1rYM
kOEs3X16CLgmYs3auOTn/gwITzUQ/OFO3EA1VSS0Y2RlFYLorvYkv8E5SkGv7/3omfJYJ7DeRONU
Y5nb3kfqrMEqop7Mo5L4h0b4hzUiGvMEekfq8vI5HE9hb+GV+RZCX6XeFlx33lbrC6GPtg2gxmWU
gy/mWxpIGyC7P/5BgcAVXV3Y2saUOnXMdM4+SYpRXoGH9QftB7nQ2NsM9UmUHgxSuiU+uGSvL4Dj
vyedoW+AmJWpXC1tjCiUdQtpg3KezZB2vMgzBczO7t6o28qRSTQg1jZM1yCOhJLkFw9rxZKGskEH
x78YINKhwzayv/e2pdu21RlybKjImnko3RJlEamyhDaO+NtVY+bjBOsf9qVE+scYDnL606dEsHVB
TRaEYcH3gGkUTb3TSTu050vqksYeGbF5zotBuHsl0luB7jD89TT9Tqzqq1JDFOOLaeSN7FcBH69L
GuiZedjvQu3/VG6DkOOykDkC6HImFJ/yqK1Gb7CH0WE7Y/AOUPFXX/u4v5WtBBjedAM0FQwnwFXc
Ugu/NqAVevQUXBmqQaMRU/+xQ1d3QbSw4B1vaZMab/+c9MgzWI2lfjrr5hNu5MzAF7NmMcx53Mht
z2Nvh/JCwxpA6/27NOWllF4ws6ruTgw21yhKVPg1eWzKhZ1QCJrld2mM1ctdt+O+7R06Unn95Ti6
pafCXlSJ9sRsAwBJLbDTXR5KZFhfD1JVSUaLB9HQprcsPdri4ouykmj9BcKHoO8mfZjE/sFUQNwT
Y73Z3//EEv1YTVQrgtJJkDVxpBHUotsSGZE4dCED3RnfnE9T/x5q0iy16vLtBsB8qJjWBIH3cqYd
i7myP/eK++OyfqQkhYPvVO1YWZFWqMwPvs2/GI1LjXW+zMU0IdnCw2PmHA8uv6StbYUSfNvQZ9sO
KBSl7t/D1yXm65f9vxss6DGHmTvi+JuWHaNmXjktGtmZpsmeWaLdQyHJ032m8AYqgi5NpMZTTMN8
7FN+KMxIOphT2kDwuDFm52QY6GDl7DjkDg/mTSSn5Dv5NBd31vwM0P2LsqgR5k9eP+HjB4iPU4JT
o5sngNdBnCoNynJmGE2ooYe+q3ERAIcZ5xaSunD7VpBGgGwuCruH2W7QIVJ0+rfwvuDQHARsIArA
Tvt3cpX/6MD5GnA/yPrgfh+pxvW9Tbj/wsDiOvj7K5eG3DxbZaaBNgd8ORJ90ioce62ALNG9QNUP
nazO3q424k/kj8Ye0oc1OxzYwrqB6uJIMcpzuj5KI6GWKnyTDMS7eLFKwmrpB+ZbZohPmjc4AlEK
rR3y0LpFyux+/tFHZw6HyzyYSaG0BZ1vIH6g/gKrHBqFixOMELKJHH6QeUmpz6QiPYnHy9ez8KJu
We55FGj9OjcLEcWKwqk3hooo5C6/Rs82gAv1QT988hRICl8ipM0nnQ9rLU0tSJ8+FumpPamsQE8y
zBeHFshW7USegAL61vSmoZfWYSNiRQ6DeTDJCPA61njOmdVsiW03Nyi85WGVlA61fG8DzTGMVFV9
SjovnwFr3+NmxGU/y1rT11BbT5gE8HgJUH671B/vO+ZbJ09iiGxzEsOEGnyx6ymmODQpdqjvIwuV
04AMe6/tvKRSPL8G1euXYU3Re/d6KLh7Rx8DSsrBHaCrraYXtQA34HiTr4StuoXrpTwxVx9I89R3
VdlHZSe0oyCREQBvL04dUYO7EsVLaHbckSFps4J937VelkjW6pqGHwgaIkH+SLtpPysI0y5pmRJZ
IW7qYILYRoog7kux4rAGoB/9boyD4JMRT3b4Lm33pDf5Cs+9DY2AMumaDCSjt32ebBqgNpGwNDNl
5siWWsJJg8rXgPJaeCmaQbJMmhMdvqccDgnJixoLw/ve7XH9es4Qx+G31S9SlmQcgIb05ITb66Fa
kN8Py1tvcYuAhQS4FIIFx8hmMnVUKWI3UCHiLSWsqUOdKDM+SZ7bpcVLj+GhyDCgIQ99knWRlexx
GM2rqkWLiv7JWPP6rYNMY3HBFbTUtPuFhb9RPVQY9Ub5f5jm4fxmU97yBj5GSzh+7z6ts/o4CCfp
HIqqq9LWk7L/Xehl5rWZeOTKskoN4IVaguTktE9bGmdGJkOS//9yrAj+L8MTu5yt32a44GZ20Hbb
nqoFaHHcI4ju7P+MdqQxNHorhbRREOunt6cKKUMg8Yd1QUVynsPyzONQLh7A217VhZwRJHBxhwti
eNRbkTDVK/aSgFB4UrLX2aYuuwQgOrgZX5GFP+HL8o1yQikruv91w1wTbWmatA4HdvhNCXmzEvdl
sGdvgubevGS3XQGWuehMFWXck/Q/uiJjNOBl7YSPWKFCntw856zNvNyPXTJ4lOy/R8YuG7Gj4H4q
4D82ul+BioPp/z8k+uYI92ID2WGLmpG++s/ofJG+nSTlDuV/sMwCxTaVCahus+fw7+P1Ih8rGCRU
Bu6Hq9Vq9oiU9hah2Th2EBkD+HnTTbqWchdWX+8AF828Q4YSDH7JkQCQZc9RKMDF0K94u6DD8hqX
y/5t+ZcmzetB70brune01k/GMY1TxUsoENT1mA7ChUnaJTcmM82wIq/29+FrGW0VoBLvh7NDUcg0
7OWsBoApx7EgT+3jeank+fivNebnczFebED2QQWG0pmIt5ekN/4Rhwzi8PuYOnbYkeXQERpYbr3+
A2fGBq8yBwDfzdiF0lE9I6DlxgtdqBy8+nhnHZbX1K3tD/RiCDbQPnv5/yrao6AMB59aoqZlqnqk
+jx4IvjiQfHk4LqDMc42a1Yy6sAseZadixE0oTzYwAfG32lEOVLM6fWxYlYeNv/OOzusJ+SrdhKJ
A/0yhG89GZeHyZ55lY+M1bsn6duRfINVgENrNs7pCLaOkSp6IxnkLIFfsGyizqos9bGjEz+7iRCA
vj33QRbUeDQTAftirLIQiFDEBLu2lrDTTwXDNTd/iKlw007rajgd7vv7W7nZ1+EdMU3hDzWOzbjs
rdxMhTfUGyAXewn2Ex6X4e8bt9juVF0nUW7PU13xY0TVwxKaUNDHtEK+527r6xkAwOVY1XApHBpb
ajnQBrhNZkU70GdpKM9/2/IHsEsauwrEmH20KTvOSAqF3e7lk60KYeXPXahxyc8u/kZkW0XDtVX1
lshvT8xJRTeA0lFIW/iENi2MxK1bIe7+phr/3nNfBScgQJHYOOYQFbKBKeGEOX8a5ZDpznyQYuI+
7y8+9bYW/kfpNlYgazXxoxjkqnWUQWNYXlM3vTjcFhw5LBBn0CamKbQeSvP/b8NvlCMZIJdX/3B8
KGJnmB2D9poC5MX5JuhIHDkttYZqdPsUl02nLo7npHnGHOdM1lZSn8m/71X8WocJAkXuPmn/UN2R
dNr6zK5YKSdu6zHDy/2+HI51asvw3VSSIZ69Nkp1cCh0g/j1bypAa3sSpCqOcwrAC8ZCxI2X45SQ
krGYZppF5Fr7lLWkqwemyMGXoIlVcw+1m2MR29ZWt/MkEyBThv8bpYGRMe0jzIKg3e9IzN8usrKQ
yqg/IHnkPBbKhaZ84RAWJ03XGlNvjxnp8EXj/TG7rWKrj6vbD7gZTVjY7FLI/louiEXaeziRElLd
uAEQaSe/7g2vYn8WwCs20Nqu/rAns6PdCTQKwujmdLID0uUaDhhTIKgxbkZd6TnwGn91cy4YZuqJ
ocL/Al9G7QU0Me6jSG3NimoKNWu4hGwOXtEC5+ICoB5a8PhPDSEDlBOMzjgfh72Q2UnR0ZrO2oct
Zc6Hz+DDhFrWaaGNh2QAvgmuYLQIHS8kTSG3fD1qPRuHOhMmu3fkrQDkrIKpG19Cnq0WJTlRR0oW
CqaWYhfTDiwlNg8QkKDtibQrcjMrHHeM3LhcKccZ0LsPCOsSZGhd3+ZYxqLxDEW9lp0x96+B//jw
fynPdUHI7YtKvvv+jeW9bLn9X0CGv0la03u2gr6SEKuzNA6DyjY0pk9zoBTv1hP4TMqJR/sNs4fT
iKi09j1vb4Qttm6YYrhgiBNAMcUZXjGBoKmzGH+Bc5APb5ITXIc7cLNVq7fFnFrMmg6Bl9JwHetG
qiI9DIiAwwjejNLunGO+Yv1T0w26NxlFDcHoIjkkD+kM3sFcT9vSwtCdSHeerisMPU+cpPmDf7q3
J9Pw0ynifuFGB9z0z3FOu27kZVspLPGMEAoEfSaMgOJnXIhLhaR5eOU2+I/qAdUaoDcdPH/B7sWR
IWGeJ07D5FIwyLIDyroxhkqVwrPFomg+fJY+WloWjWEuf5Si0GYHc+TylHKn4/TYvHgl0DVWMXuK
wh8PrlNx1GqefgecTfNuYs8Px9GGQ6mCDNMCBwM2xJHGzluf4I9IGMq8xS3qwe650TPP6rImDhn2
XvCoYnMemJjuiWr7qSCs+7wN9Z513ZHYeOcAgFWkqneLssw2kJbc7sVACiVeAg8TByQHCZMm5Gqn
LffE0XjHNRRdl9TEP4v6xlOd76LsGWrF4vqYoZ+ioGIUhNq/KNQ0Kzd4pvImQHqMsJLUZ0f7/iz4
xYCSM3pHj/LS9eFresTTZUWqTwzc4ljvzTcTklh8xScPvFuK78ej15D20lINXsRK1zxz10+DW0yX
7GaBKv+wesaZiI/c87z6IzbMiNfQ52++YovCCQfjzTaQN3ZfLv149Q5AZQN8WcgPPyQCUOZGwVDY
dfqjfxmi4fZ64xxeFz8e2Q1uKv/aRMpJwph+qOncEjG0dOQHGLYwMOApw9VtEbB6EspqUdyiPR+x
cD1xjR4qAT0dc1pPBoN1tf+F56b9WHwusBuA0nRQze5mmF19gJ7oz80iH08CpK37Yxh9ZIE7VLyx
iz+kMktz3ztGPcCT30oxl9CV05p9egigQnjJbQfm7BIc4Rd/3HehaYj06+hVZ6J50b0OytnK+UoA
cnK9RgBgMA9/5jn3RUCXxAG6rAb1RsPpbmokcKQ6r7jwl9YtpyRARdpTNPU5O18yV67eXRmkrQTd
ZwJPkFAGu8H8NXz8Ik18UeOmpgnUk7Ta0W3GyHoUe3cteDPIl//T2g9xn8goxeKLamcOWIsi8gZq
ceZveeQwLCSVDxfRoNOGKUMd1mjfBTHmNvfuHdQphiy8xXVvotD+1UBb2VsyUM8xGEFJcJTu4Ahs
0tYALupE8rdrOoe2jb1WDDiqyKe1iWTG74KMdXPiIKgY2uMWpc3s7h1NQJu3kmTz+A8EE6ecDRxC
mfNa3+emK9N7lSIaw8jjwRGyVcsyhscCNIbOijCLXZE8EFqZ81w6wEsXTDIjGkNsmOnkzSL2rC+d
V4YjBRbJsyEe/JNmTwasKUr6UCTnr7o4z85yK8rECjv9XiQUJCMH6yH2yD2pAN8vGc4yB1L6+aU9
Z31hoD8fIzqkSp1+Pl+9ppCrWRS/J85isx1gYVoYHZIk9UEb6wbl1ScvRYLDTx0tdsib8yp41G9h
GO/np4DnjNPwusnNDGZk+XYXjega4L/v/Vj3l9fx2QO/qA7I7f9ymBDPoIkQvmvskr+y8nNMIkEF
3+x9dhG1oOzxyce3VweA3qLLILRj8QI+m1Oqo1Bno8c3FaaX6/LnQp7fiO1Q9L/B9aPLdcEA+atM
K16Rt/RkJ5x/TFQkWhQh2ZKtKn4Ty/ttv8S1LkA9/8X40XlQOUR9Vq1CI7cIDTq0KOWo2S1lOTop
U9uvP8k9FgOKwsgYkDT8ERWHqVGDSijKgTI7i++eN5GOl5NTFxeWO0AQDJvlM90p8K197D7Abl2M
1kVS3/u3BGYQIqk6aGBhTvejXVu5cXAf8g9qytzkOE2ZbBvaj6dgDkD+zmnyuV7mCfzWCz1t8s90
KYGswooOT9YWr+HdzVtFwo58bYl22+lNRaOOufQyuVfS3GmFMpp6mdNRlFgg/HjV1ucR4CgWQLoA
dqtNvOTedn5VzeJBSd0B5OpPtS8r+0n57iPA7EPR4QMNK3e1kVg8oKvv793/kgAp53/9wvd58BIA
wsiwSn7lVpjE7EMEl5s5SRahoOKKToXPEubMuw73MDVWc+8gCNAn8rwiXwZZ35pHMyG8SsvQdlWz
wkCDlfp1qSkb79kc77OHOWBOuO4Fp6wHrHrud3lABcoQZ4U/xwe3VHedl+woL2nyOD3CR1uZ9mgQ
xxeUV+HUKLwuHiaLBij3gPpDJOwEmkBkf1imXuwfzCWkqI/T7anEozVtM8an0gl6kPkVGfWjuDQd
jX1MheI06+/sy95jvrRJjjb7+I9EECiap65BaRSDuLHDprg/B73uy2ovK1+dgiohOGyBGKixxo1g
zN9S0A+GjAkUSTW1fKWdh0SEOUCeq/l/oYt9QPGLGfAUGS7e+S0I7dt/CCSs8O6Ut6VIeMq+nwaU
r7tHnl4+VXE8ejK/7KvkhDap6jJZ/WdhPLx4HTJEOHxNRlC/1w409H68+ihYQ2rdAXaHwz6Gu+1m
3gj5YcEDSv5cpcBrTESszy7yk6fiyeiTH8kErXsPkiz83Qd9jdXOTT54UGMjkl5Bz4NHMHD/5gqz
09PlYoWXpG8+2bAuAIAbPQ9mjGqMkzUDLRU9j8+zp0k7+AfeJ6OAgIxqudlhmP6eYkG3nDgHODlY
6EfN8AtPRjzkpM2MoauzUluKTVbHwEbqjSzMmaqBMZxqo6XGpXk4YJctDmqWsOIFXobXiyHyzHHq
PKaNbvKOtZil/UiY//qSYvnJhSoXTz/FD1CThVdqJOXKHo2RA/Py7eeEmhN4jYrzPuh31NHXjmZv
G0WY9SJ3BRq4+iblS9TRLlH5OzG3t90rTSq9inHqqxUbtIeb5k5swd97v6Rgzo75HNGJAUpWNGqq
AeT3T2A0JvUKFLw75MFB0B3PTnSutWmBelnU15tOq2VEraGfTqGEuOI9HhDcnZfelSukqThodm2z
VAa8i4zcgC4h8YJb+JHFkc8OBcLRuHCQ5d76CB2Alc7YXA0UWA7sXcGPy1qqFWX0rPLlGl3nR5Cp
1xbAHDgTNY9/7gSjpUVmEs/Whpn48U3RhakQSlzoERq2OoT7tcL+kOxjYrgThVAxklUMIQ9POMVj
FU8CSVhhqZb4BX9XOMGgzoTZI/FIN2Z5SaMZMp5AJWwoZtsRyfwboHC69EG1z318PiIapbevfIJP
fv+k95vI2Y8Bd+zrrKPBiV9UbHFCuVZMVp55+XhEbnTaxO8nLYLHrCFZixiyI0QWWNUe6iz67RJe
24OPYxKyw1+Tu1xaLh+NwaRu8QyTcLocvGVbPg93/6GoeiW1+7FcqmXr1U6EDXuXNejdEobrZNJF
PMW6a1M7NotVQQyUhG1ykCJ7qPXGf8XQ21UIjRoTn+l71qkaDm+1fkeDi6lpfr/bkAtoVJLYYYkM
do96VCrB3LCUUVmhx/lWZwWcwGyGLW+7/z6vBcgC9w1ccksctAsuuNYrOQBS6fVctzZ8zFsdKdxV
G+4RBxAJiGx5Gr/f8qFofFgOuF598T3jLkNP/M3Da3SRYxpBq9whkZWJPN7kPN9dG5Q8INuROqAc
WsdJnP9AyDcsJg6PAj3ADBl6Rk+XLo9+Wm+95c0nEnqIXXDFbDrf2wr3ISsw2E95thz5ulzi79y2
xPiSO/NSPVp2AA57w8URHAZ0FC3LU65W1FXbLNgO4XG4YOpd0ZW3YikliVKmWBkvUH08uMmxcLgz
xldNMHAxG4IUm5iVW+zE/OE0Fg66sQpjJTIETBMLMZ2uz/V6SsnI2LRmspdziilNSndNmrXSao47
Wr7UmZ8ZCKgMQn9HcX2H/sLXuUheMfcBvHS+l07nMrQuJ7jELeF48P24b+0Y7kCXAZO5JbkCzicH
8CMHGwrIyAUOVnoZc5T8Pc9V75WsuJBFFJJenXLZjUaBZyQosKK/WOekh08AXCJdxsiyQKP6IM7F
N20zh2CwBEDQ0p2rc1m2pPWKKGcT8WSnehVi/Shv604qkL2JcMGHhE3tijcjuwN/037JoBfzQkHa
b7Cq3MxG3ftBxsCo/DgljQahZcKkVFfF3bKwGVviNooCxzDo1UY7eVpcqFjRTAjS5R8iZoHsu7b9
xPd+zc4UZb6uIf5j/KgoRs28mBp0I+mB2RwRhn+EAMaP+0xpZux0kn3UiURKdgn2DkphaiUMbMhL
Oofd95JRJAfqgGKrs1GYZCdcp3pz4CMksQxZg2DeoZ6FV8HKNksyu6DH3+dU5W67b5SGfWkw31xR
7ZCNa6foqcdWp4wzrAGaIkGPClrc/UXY9XHe7wQU3vpS+XcQGed4+1La/tE8XBOrM1iBjJKrRt9l
vMjx7Bx0u1eb2xToSgqBT78Bf6aPPzIQsl2dGCeW5zTKYvR+MfnKeVSRohl8pO/9rG9KB6f/sltG
hyqfqAaVf0YbHzAYlmQoa89CLwSrVNzgTHeDnbYhXrkX7fTX/eyCdbQW1i5SuE0F7xwMwZo1Nvo5
Db5oqLi+g0F2Jnngfz+v7gua4BC7blXyRRmDvNPlDfgowESCVMZzYMwP7sxz257yWWo+BeHp9O/S
TqXKUfUvTNIvtM8LibVebfKd1LSTulG560pLlgPi17WW3kSZp/L44VJt6Ap5QPhWPjq7rqSW2nIX
W1t0VfC3X8iyYpfLzxGN5AUYw4VoygCRi5vtlujw+CFDw0uiWlMQaeh8rY4LOCRGglq0LgoeSnOl
vN48VCo/H8x3oX5h4piVFql/rebV0JKeaIP5XKeRvdLtYDkxBF3o6spadfM9liayBVJyfwSwWS+7
1xP4FHRp5kVAJoF11KcXXp3k3NZUhUe8Xkf0QNU1fiJEodLCTIiXsj5+i13yYZV98MiFK7Yor8qU
zQ2RvtIG8k5uKTl8wK/Qk5z9p30TIH31eo4mCOQA3mif3/OPwj1E6pqWz6vcM+W8KliR+eouWugJ
eiWZbpQMaQQJaDiG7UxLYae0Fxq3e+x9ktYH39+mbf0wXysp1q1OMmtvTLC8WXNiycYRQfAivb6N
G4TePdTmdvaHS6WAL7AckzasYHZ8TJnTUVtLxefpOG3VyOc/uTBVRzs5wTf+E9spSshCx/QMsWAF
Tpfo+cjNBI3pSFxzQNx5W4WWssjnOPaCl0zRmZQgMJt8Jaq0yvr49q4h42PYGlPezl5Brt0wcL5q
EACqfV+SygjbV7tK7g5mm+3Y1NXZchwn9BqM36xXO5bLBHSeS862yRGpc+T0q5vWcR2hTLsjtYk5
i46grBsZR+j9ccdKsvpm8HxMv/UeCoBfPk82/h4luz2jc0R/7JVaHjYmVLU6/G/zVSSzgnTlYDTI
cl+f20FcPMqnTBF7uIA7tCxlyn1SBYC1wcTJRmRotCwZUTJlYNXoxY5HdCF7pbJXB95QNjbWSVYg
ZFV5N+m1dFPbv5Ph1cc6fM/Z0dDTfIk5G/s5zu17saXTlVe0gQHBg1bVN5ALyQXDjaLvvZ31oRyH
1DDlnOdRz8z0Lyn0LAdo3iOPhHUzPbxK0k62FlQAGuPgG6S9b6aH1O3N66m10KrXCvkciRMhsIY9
1YjTKKsMeJRlk7QDLtF5+U06WXFrvfF3uH7ophze2e/Pqnm/JDM9zNoJmkmGBTWq/AHOVevYZ+sZ
c8/SzhcvRty+XenzSlmozCqzUpQblV6RrGVIjnHLwegQE7IYqOWb1zKH5Ow/oSKrhXDl7kV81M2L
LScRH6CkGvTsSCxkAVtc9Jvp6fl7P6hdX3eW9bj7T6EFK8zObY1jzqNNklRml9M7HNBCksCoXOoV
Jz/7JqKhOrMxA+hcC8hsGofdVEqTfVVYsm1MN/Fved+ksedD5MfmH4IHFcgeSXdqx6LQwiX1wLB9
cxns3YFh+5ZNe3UI+uFZgvmKRQ0XvtV2UKI8VC5r5POFuEGAlJJqpZNBgoHRg/U/t1wpA/2wIWzy
c1qwP/Dmjyo9s32mxXnKXuOy4kKKMOCNcuAlI6iORsztSOguuSVxBpr8sn0FHViytVl4b2UIaxIB
TuDelBI3QD7b8Vigb3K58TBiUsKe9WGs+DV9L7RN4inCv0XRvxD31yDfwVgmwnhrNGPfcJsX+Q8m
yvjIuE440s4bCMkyL3PxmylQnjSoGYcsdZRiTTPeSDCgtdlZkq6CTDkv2nUiY2UwnK6YHs0t/w/u
JB9TxBFT7I0iaM3BCySy3qy0yvM6auFF18itz4/pmdJFFk1goL11lto+boSHEeVmsjF7kTYCzOAo
4qeNl/YorixdzN96mRkAUmem+V7u7cPxG0Pgsu1tnXBZLGNixwdo0Vs6Qx6lUh6aOXCZlsycXxqR
KjbFTC9Fb24PJy7DYgQwowA2JAHwUsKJISlU6Zx96/pIJr1P9SGQvVD+vRNXGPvUmsArf8enyrTT
gAQp3MOTaAQzJaYZ5La1A6cfblbnOuihcSWwI34m66LDxGO4gaEwDza3iFvsvOlrWe2yyZsfXHYa
1Yg9uThGJZ8beZxP3jDeodgza1kmkdI6e/7tY/wtxnlD9E0y+MjZOt55b7ewURkaYWsNOitoECBE
QcfVMKtZmC3wF3HBjIbJVUNQ02BFXkN1AD7fPIJwyG+XI2lojdJ4exOx9sUA9pWiOpry4BA3Mq7S
4fB9r9SoGYQbufkDVj5qBGs8GELF56HFFiwNb5WB2fqa8SL7nLI+e/VPSNASqpXPvtC+uJxzM5WQ
lr3gxZrGQRGZaxKjCHi2XFVVr+YbQBuF3l5YFeAH8PGtAQ0yaXwXuPqlx+eOux1Ff3wpU627JwWf
Scy1yh4s51gattIDO59UGz4fHoNZizdZGd9co1fIUQpy7ekKur9PlyE5AQqSmakNlcyeAG/rDg48
xdl0dRr5UfrYOZbs2JmZitulQ8eKMnG4oSHK3ZhBeOy9RakGYyzhh5eNP2jssaIGPuustQ3yNr+2
ut+hdGHqRHOel0y/251ptbz34mC8xDbga/h2WBHdpJNMvbcLqkv78v+6w77ZLevKi2cWUIYGVujP
msuabs0klVzbKsG1OMDjxnZgveBKdWxP4lI7zMvjkCy8/MghBvRMRtCTg/6Rr4ze/ehJXvXRlbtO
PXatjTQWiMLgpyMbNRdpwumeEtukbb/IaqNWXJIwC8WD6F9rn7/wvb/fDzqOhOv1ulgDRxlC2/Hb
2paDkAGvKFQllHYQL0tMgmqfzaeoC/m8JUA+BJ+L72JVi72rlUnLyE1I/x0yn4+McKhGRQWgtgQo
m41S4ybwSms1tEwYyzxPiTDYBGi03Fn38fcPEecqPSUHbjGHWayqUwHBEkmy7GGJlrz3l7ySLfwF
yhZTreUJPVlvSCzYBNfSdNwtNibxCB7+0hXGRIifxkW1RtvqT8+xo0IjQ33LEk64fQbrJUVY8KNq
Iiq48EZqcRxa037VQ1GCJ+C9+/TIVxJGaLZa7t91OTUO3OQxv03aqVUaIuuLX6wq0DJXS5D6IKQi
l+0v5KfnTT9AHJUUHGzugOuDZO0dglBbCF35BkClvwZtevgW5kUDU+SANM4jNSuM2CSVr0Ou8Yen
mQfhMuH7QZ7kECiLAsrrOB4bi9zpRWfkH2/rnSSdbuJhzzzFPicSg5LBJRrWvesPBOIpEpLQi9KI
JFn2pUQ0EirA21xmWMGcaw6UvIDtMqi+Q/SMn1ZA8hb8Ke1IdHD4e2VvuBtgjwe89+NkPIOxxGUP
cPdRfDRyWGprtLI2Gf618kZWwanm3Mjzo7AX9Kie3bExbCaYGTdpdGZm7MzKsU1jX+sjyA1vYma1
nygvOXxo5P5r78PNURK+DfBClhVMuyWczPxeV5o6k6NcWTupYrQ7BIGsWjIEeffJhNcF9BvTw1Ei
IRi0TK5BfcB7bwbuKnMmuefr47TOf2o+X12EWc4+226DiAen3xIBVyDUnfwwxcAMuWBSwd4k+hSD
qeFIdL5k40PNlhFZxAWhnCZ/tH6aZGu1khl2iOuKnjuw5CegHS4aJ/B8UZJfvCa2u4Pk/Gs4d26f
by8ytar8BQfR4BF6yOEuIhxXyc+1LPoTcecP4b/xBzcEyprfa+gJtvvkwkWK9+SNL6Ghf/XDzcV3
jCkQQEDuNNkwMB/fejN79Nkc0Cq1s00ThqXLHjc6Wio1W/E+HMjPUxzVWLGTzCxnmEd9KzCBElqT
3Nm2G+wdzpX7pALI7JjqYYPhnz4baDU5ie3naG1Bi8yooJMFlCqBBW7xQ+AT5f8oJC5GxCOctHie
Oq4Xuaa8gL1b6RPC0TJYTs94OBJZFSInAtYbsosSFzYY+Y5Yx+LFCpv8LN6Wgq9P/qRNQc+/O5Wu
qqruz6czyhCVlJqfcDwMOcyHlMh4V0No7MM7oclLS8HK022AZX/OUjfokSnuXWhSFX4Rpg1S264+
ZvERAdVCEWNmYonVs2zXAFBnLFi9u84hF3/q/e8w9cPUFiPgLMAz8u/5aTa98grH/yaTf9mgQEKk
yqh7dsqyqtDhak+OyK4zrDofL9lJdFdkr+kgNKNZ5gf7+Zjvb3DGWcA+tGHOv0MJKT+WdvRMQtLz
dv5AcfEPjfXITqfV8w4CCq24QpZWGyVwYQfMS7/lWarW7+EQp0twEJCyrSEJPq3/D3yWKUujtVS+
r/tCDb7SdvPilaGVxHuT/U0GoXoV+l/7sptyZ9DhGMDeKcKF8r0tyj0lT9srTQEL4fZOkG2qpaur
9nH9GCAlzMFAicFK2PWdK+Ta2/PlYkijK2OJhu5NBYp3S3MV7KolPYzXOwQ41SdJ7wkQ7bYgMumY
ONjDplDfwOfFv4qQrOpKE2qc+XU04JKha2Umv5zSP9STcjSyFwMqPATzNfhFsRl+2UnVhGBbuSOv
Wjp58Lf1dBro3sZnxMCg2xoJg5fpzUpIVyrUjKMlDsgkRT5wZ2e2UA27OxZzw9qQTulDQFOgLfyk
R1rog+ZmkgRREab2y9fYGXFg4jmDnfBjz46BHLMwyvQEXG00+EKv1uSdVf3hh8J6vCY3NNLmIHcC
9Lc+92tbntsIbKSOg/XfBRdyUCOzOCmuh9Q/75o/pR0r1REbTggeheF9zDQ0qBVFoQijxtCkcNrX
r9WNDvfNh3DXKMju+r7gp0PqRXvWZelesEWr62IuUSMrXayZzB5gDCFjBKDSuEyTEv3eredX+9Vr
sNzLNxhjquekjLkxzHssvlEn8AFeIHzekwSk/ljXC+IBz3DAdl0ms4n3kS/IoFIUvtghx7haN8CK
8S6zJfNDEHr7326JMcVDpnEB9XqeFDkr1ujJWztMwkOfh8XlTqcIwZcUHdk7CrFK2RGGV///rSuC
uG5iRiQ1TFEfbkliS9urdbqv9PQAo2t50JLR7w8BkkAOWXfFJ+M3hy/2Q7b5Qx4x2tQYqVn0ptLX
m6Hor3Xy5+BlbAP4DeC9tOvpiDUwIrM4pIviNq2Kvbpsm/Ty3mbfC6UgldTYwZqmxt0yMkzNfH45
cn9Ryrba+bVdqedOjHbdK7z17NV0EtxFBRXybWP1lKgxRLvrgt5AUyWcS0TI5TVfPtJs/oZYNATJ
pvWyqBOzHPCkir0EPc3N7NCwwoqoXmspxq0fsk9/RpuNT904Niy6jX7gXuPKh1JMmoBNhelB9UyP
j8R8jxWd4+a4AO4TL4/yqMCj7CPPWM3+JgbhVd1F0kNcdy5nrZVDkmxDbWff+7wbA/jBRQ/z8bQT
zDsH82uQjo/KOz9pl4Y3OgkP76oprGqLK48ZwVLt84wZo4bIMrd38pX5BWPPLHtj1JEGZG0ALU89
JSVC6H1x9fsY+KMt9DF4c6F7vKuMt9qUVDj6TZrnbymt5ec0N7V7HD6fFbvLAUGsVVDwIJuQnFb1
0Tgs3frPVetNImS2HXoKjzeoZRyMy4TPLpHTf1r7DX6TFd803ajMf1afaFgqzS2NJahUnWnnCH50
9DvyVs/rOprON5QTVcUbmQozgpQlsid8nRVOj2P1XOiRGWI3fmOWADS7n/X8a3We+KhD3KaewOP3
8TIbDPHMLgoyOXEIrONl4RIgixrDAc3ICCXwU7eaqeXubsSAeLxIViwJbJ4ixDV8xMyMkS+wW5pU
xdfljgHxTAISx0x3rVUjV+4P07DbnjOeJx3meXO7r1vPm5FBftxIKLsxR7u2ofYYOe41EnW2qL1x
wB+qBVYy6ciLbTcXF6AVBQj0sAdAOvJxsAvDiv/26igMoAUp9U+8cU7+IsDtB7X6SLQITUQ+bb4B
4aZSjCRYOu4ksWRLGraX7Eiue/SEiyDuRzgObwDDRuEpXeXiRaGRLKbQyI+mGMfm7vqg+mdxxL7E
nP77AJujfZcHtpW9s+n1W2v2ua47/xU8zkRikRE+JUINuAMT5rTNgBofZb2qiiDD8sPw8Co8Dif1
Vz5S2blFgMY6+2dlSCbxhuSdDGU6BgDb/aMWkEvSWsr2XBQSZJ/AxfjYJpi6mlqZsoY8aNDV48Mf
gTcGCZSYm7P+InA50YD4W2iy/KxFQ4zqcZ1gFmug74CDshURssKK34RogfbIYojuXaLdRB0ey2MD
Bjt7OZeg2tJxIDIf4Bvs0G+N/pQ4E4bw8WNlINl5vxYNmNJUN5LEuIi99ms85JNWT/lczLqgBIAq
khcsTOq2Ed2JteIG1qcznM2MFGUE24ngr22po2sVs/TqeBtwWf7956xOJa5npbOPUdOSM5tXbCb2
sJccYm1a8iW4osPzBHxU9Jr3d+catGqqhyuWAqh2gW4GRNASWR2MhA6MxhS8nIFmjgwIB1L1WU3T
gqFldIqskh7YJHWAZ/QEh6SIAu5XynTrOzCYTWk8Hiy0NzprTgGyzCotI3uFf4/s6uqiycJeF9wG
umw6ebQriQ+pe2s5tTrTpoK2ptLltKiwV/BNpxIdyNCzW2XSaaG7lP/RushTvLuwXJo+EugHiePi
W1YI69V6P2Yv+or4y9P4zjYJp5YTnexqyFAUMB5l9OxsWis7eR7YfW8vckULmPZoPaE+28maOkn0
2wOBo2Hgv9fL+06Z2zfa90UIFipPzuQR5885jP9UpsrsnJ1sezeIs1rnRlw4uqPf3GGwpLLs94L/
BpGvSQbWOwCgjeclcTflk++zcHkJ8QdgrXaoZJB4dh+QIrhIyyTX/1eDCLsswzD34RM4MYMk1TCV
9V/RBqUvLiym+PZGRDHiH/25S+9pc8UunfzXW97z9hm3qBOetcfZTCxtDI2kzjUL/ynvZFNdJctq
Lbuw9xTDTIebPtYj4NUvPo5sZLlhs9L8DIhUtOgu11oazuCE7Dtg5p6g+bHkI9WPHpFKcNLOEZ9x
aWg+w9LcVotUMc1zEkrwaRClCZIvxDuFO3sVSisiq2AHm5YZBE5xWYPvO2mhU/F68z0e/jYgLiGh
Fm/Nz6DSTKTM+aP7iqKUxdElCHF1A81URTxzkR8DNco+CKX5LsWxmuoN3WC1R7JKRHkf8eV/Kg3g
KnzjT0h4MLwzHEJdiENTGxA/d+SZmA679SIcHALkCEbfVFr34njYoEQ13IMXqyGg+pRPW1tw4PsL
fo8OeoR237IPRIbrDd0NYaRz4N4gWAnqeKVTurg0awZavCuG+IVGolq8EkgRNLNBP5H0sJzrrxx3
AS/pb9lCdXEjcqu84e6LCHu31EiMmyuMCUiIgAogaPIJD7BThI55igREQocsC+qivHWRrgC7hsGm
vTkDIAmKOW3LsMDohhjmSmt8TFJ/9/dPQawTCBZusslQDMboqCL3mwWVbHiHkqOssIOxLVTIus0z
m+5h0K2qdcxIeES9rTTUAzTJxopaLWA055z0VspQXo6vP0S0gfWwWsdqRB7ul2IXTrBcytbAK0NI
jn4upOom8yMDP6K3HU9kCZPF3xZeHIXYQ2Zx9ylgditbVIEBlYcaSlhrXcmDRGIWgZCXI4NPFq6K
VC3Fmafs78iL0QRQsdV4KwDRAbvG+sonApyR8iwau909ecnVTv+05awVUMGpxMZaXvCiiTguY01T
3TmLCChH8QXksGExlRP6VjmW8wqUUvZh+7Yie2gKI/cdvNEfILnfWuBZYMmKKSy7dp1kEv4Df32T
Q0OrGKYUKuAeB1DWJKI6WFqwsusX8BhQ1VOUy6wMFZ4mL5IrCvoyKgOql5wipcJkOJI+Zf3bpkWG
49voHAYzcRmI0D1q201KgOPbYdWDLHAv27V2fFsJjU1K6ixKIbdJI9chhRPeGw8jngIBfRCW3gIr
cEFwo+0e3sVMqqYlf+W6SQy4PC8DSrp/YPXoCkh5X0rPG0xwi6h11muzWLT4kqo4HcSIDie+qYVZ
UJcgZZGnKpIi36RHPFeJhq687fNV1pKDxLh0/EMqEzrisR+Cwi0rIP9Dy5L2NdvebbNUMS1XustT
fBvK51uV+Dj49JbplCrSwUSuBNJu8XMOnxrdY1OwEO5sC99P8e1kyFUOe1xFeYgzEXVoNhLcwyuW
b8qR4pypEcBbyoBlfsgTuEIQRG1+AOuJkQd8r6zU85yBQ1p+SdR4InqLaPUx7+94XFxnzNiAOi0Q
ADPrEI2NnTNMSv7SSseZMv/RdeQ1Yqyp5+njyahN0EuQYc4HxvONmlO+CjV9Yt/Xzqyhc71LK30z
lJcNikh87jLT290+4fQXCfNeMAC3LwzQiWs0my/FFVYeZ9XFCAxLU0Fw+CFnKJFQ6pInukYgQPOf
Xb8zNS/bfj4kxXIUQ3yXZ+72mnZS7oBF4b+vL1ylgssodFdP35UHMSl41fyamAC6ao2fIZrZSghp
BEb/gZQaGD2kdMUKvMtlXMaMkD9TpxGZSCLHOZRayNMS3U/tIMTZOlejIBTAlQV7RgO2O68jxNLn
i2Dmp9Won0ihVVjOt3PHiyWI/BWFmXKRq4m69nyyIjXvfdC+G3NsA5Rb1bkElY2e9tfOrqHvh1wy
LHwUhhqIWTvwdk3ihtZHPYzHwal+hN+sQ/8Wa5KuZaHHekNOlUj3bDoXsBrn+gnlcEkVUP2MhLo6
odCbuX8hgxR2zfuQFFUzmYFMNUI9If6qMLE8mzZ0U4L6uXtBoNUIBuXIabZryytIh7+OE/fpaHIr
s6utQlrOJFLTih+m4qlAgeJVgXVehvpgdTy8MvCp/8xIqXi+hKaIYuU9dT8bqdAU3zsXiG289K60
xM/lnLHp/gCrlJerliOCuNdx7z1Becq8L1EtWVcYxMuVBTPzFrL7or4JdyyURsDEOJSDbRz6gRru
L14oCLVigVef1BFCE0ubAdZtNsKRyf1FHzDQn50Q+Ui7iZ1LMC4oHFkwwcNKtKSpXh0UxML2nKaP
FpWcscIvylE7ajAZWbxEaQ+WO4ww6WhcnClzWX71HoyuABKn+bToos7ErU+l/DNA6aSCbXyQ3EIq
3WAdrmeoLY+Q2OVA5FiuGiN8yDUwo1i+FV5MgqyWhrlN/8BQbrl0zPAX/xYg7il3R8EY5flyZ/Xj
ef5LRyLqHDd8BphvczbxqPonhZc+uLqNyH0LM2pSl8sRUVa3+HPeNpLzgriEid9Wx4HuFYPimbQv
FYbmyxRYaiBVpc43MUKKBArxVg9dHgL32YxJgDR6K0J6GTeHnfnV+f9eHbzXi68aN6q687VMJh9Q
aBCkRuwrOONzZrN1tCGw/81EkF7IkYz7wHX7Hj5BYOIvEfatAvyzNMuHKbX8u0n6xXDp09WTElYM
epuVK0z3rAIoxbfvRz9l/r8nZ7yGzPxLzdBNsTa6wkQ5By4zaG/VvLgtVDy81wSMKKQ4bMVTsQep
oKoBVHsW9SthjN32BHYBeTDuAFkphYuKpHj6TN9KEV/cfUW//8CocA0ovH53sIfgEhc8WAsGnNl6
zXUQYv2i0L47OqehZ6ubjjNdOeL20kAl0fxy291RepF+C42DzfLIEncO3TVfx5DUCChYVHJhpmnk
lNa+46FFqsWjzn/bf6U1bFguY2fjAO++bDoGbItgMl7YPglr8Dv6k/nOR4/gjQHVe07So7iHNOP7
S3S7IQp5MpVegwrE8/hb0R9a1BI2ejObdKRyJs+Fr5jsNYD3g4QI9tXnB8AjZMAiW+aiZZxu+34R
ZosePeEUIyXD3TEvr/3cTyZ0gVfV4TDTprl3cAy5rEmtoXtE0id3qt/4BPc1pg9ZHxhA2GKqiu0j
njaqovDXv63c+CYvP+X+NQ/o5dsmD7yOcsTYeO4oQGCsxiX5TO8xvpHqxE70XHSmU9cSDrf//scT
73FEJxYOXLQHF9SRmOKSYvyYKG+du/iryFZ1L9WtZHZUa2i7dCTABTy6JlaUcx75W/iBg29HTZ+m
WpAb+cKWOVZfnvjLhAiLY6rr4tjgabaXgP1ym6Yo5FQBWn5ZR5VcTogCwDjvXFnK5kEHpRkNiZBR
Y32rqFScv9aF4isOOAGZdTlVymIcar1K7JbokOIo8z3skTfeqrmpWmzw2Q4heYoB/gJ081vlTzvY
Kf1GcO327yPEbaAsM/+bpshWzJeOS2AZrzjk+xihZk8KqdRl9yrFgE5jwFz7HJ/P8cNUgiOYVyox
/1ievjMDPIQphmXcdo5QguFjfG50HW0xs3pV+fqeJTd4mXr+ZXAR72KFvRs//QBIxd/IK1ln1/Oh
p1O2/ACjycUTj+RYFVuqIEAeeFIKm2bOVdsgFRAB8VwKhsuTEGrtP+3jBxU63wsU9u9QVi94dd/C
FWVUUNTA2o22kwL2YiYaFb5r1/S+2qB3dqvDfZ879t/Q2908ITORV5o59BEQ/rowtX9vzY740y+4
JW9xZ58psFrSiSXfc+WB6V0oxjWd1hubZmf1gqSU2uzHIduf4TpnHqpMVY8YmubyRwoF9yweszTB
IKuDp0l3UmS/FhtMjfTxnrK48YHNhPQioirK4BVKdqXHQEkPy8OT26HF9WPJnV8As05L3Xz7tNIV
Fu04Hf2A39hitEd8ZllguICxnGfm0QwHHsTWJgUGnrSWggNcL+XHDNyjQons0WIIecVgQrShy/0E
t1JQ0wvcISfQXuR0v0XlCMy58jP74CoWPnalic6f3w0TQlwJLV7FWb8YQPeGnyx5/M3cOmZZKSyE
r0T+52JoiERVU/MxomAW7RrgjrvH9V1Ug+uGv1J3nFX8VTIXQcaeSKB5KhsyS2Nwcdw68J6Nw81u
U1Cm/20ky0lWijClZ6sh8daKMWmnaskgljpshNoxkPiGJAJLBj18G4NIANhOK3O32Pm3ga+2p6w3
TV1mWeBjr1HDLiMB3u8kVCJWyvG7g9vuHkQ/PbIOrJHtqSNUMcOI81U6Kqs58hFXzouAgtwdOL+e
vInZTFGkZFcMxutLlmUAaJS3QNIOWrAIZmymTZlUMhCEA6P8gdmZ32sRUmEBjp6nyVHxJGubIzEu
EsMHwuJRRlRWzns4myKLdMp4np3Gu5SGV7J5hETD3dSJpD+Hr2w44/gq8fg8fZ3ACGTIUvWjwUmE
LWU2Oh8Py2aqiIQhi2/d3wu+MCI7gTwXao41nhew7yURObJKeIqTHdkCaiIcAOsVeuP6+LVkQ6iO
VZ8VvVR1sFGyRzd54EnO3+d8RwMs7iJj9sx7Pm7bqRaZbCvJXAP30TMbJRjrQQOUdT51fwt/0Oww
RjNNKo1rVj3A0bMuiLzzvAD1dtTtGQ8gsx/8nv8TxlZ9uSJjVkMRNBxF8jgDm7Mm1DKzOT5d0y2r
LcnCDnp5irYJ6t2JddcyPvVidNUslfOpScdWBUSixXfoJEvA1QqMWe6P1nuyQNB8wx+rbS9l8LXp
VrUBOTtJCsELVetsubRx9/LZgb9G5kDvo1UH7vgh27cOSth7qidw71fw9IneifBbxf0Kd2iBpfQh
KfJBaxNPjyF82HWkhF+gLC4EaWFanMCjBJt/H2jQQXRKFr3+b+7U2GvYhZArzHb5LahghKF7ieoD
iIKziqtfrBiGy10e7GTabbop9FSDcT4bT+PsKexHSY4vtSBtpy2mpciuboRydnTLF50grT0UaRAp
0bRzoYlUnz/a8oC4STBJgtb58BeT+4eKRWE1vmKXOfoBZ1B5jAKV/2eFMdR+6L2zIrzYS4KV6jrZ
jkROZL+sb1zFJWKgeppvxZpwutMzcOHkgIV2m1udQQA9EMblyzp8j2N2TeXcHfviUyajizMOZCa9
7OVB149bHVFpKEGlhLXO+ndyAWwC+5xBtfXLWRzWAmMMFiooRd2waf0fYtnngCC51AOWXw958m44
TS79Zhd8Jsd7SbghWLNCU9HH2VGQejlqy7xjzLYvIGpnCn1fnGaMm0AjQDsYm6CCxusw/2y7/NA2
Lc1id91TnZGCI9GBuSGMnCp9e1tVVv66/9CiZnSTa/TwVNQBv9vLlBqOSYFzhBIqOTgCDwVnSr/M
exH2+YMleAdgYizw2X/ISwI3J9m6mrpqj95vIvJIdG3nRLiLBet4lt2SuZrJSDJn34Nh9yNA8lMK
FV/oiMwpPIVn1rYF7TuUqxPKbPgvCdQ5A/cRiOENoUCC3sysX2YgFqtgFHcsGo1/UWzy7RuRTkXg
tnCxRVtreRegLE/ChlnsodpVLlORMv5gHalnwPKRUu/TY775mzsc6Ce3VXHFfBlbMSICGTpWwgRR
1w0a4ihRLsUn6Mt7K9sLSkDCTU6k4v3MOr/9KwzKDxMQpGkYG3kWdP7vxxAezd7hFdaXVpwWOpjL
jC2Mqas9ZTQJ3Z4BzR5uAR4ek7gKj5VT9vZUs3T5TXZ/x/TyaKDY3yh7bnDRxE+U5UcuB+OBH5Ao
LHfJHl66SY2R2ZJpnMBye6Vpj2lcg3jaRyRvtSBeWiEtjbcUKYrHv6/uey5Uq24wM1527NWaBMOn
M3LIAV7lop2gaf45NWQD/+F1s4Tzmcd9uXimGEdWFabR8htbc7J1Agi+zt6Ew3Dt0CliF49doyGX
XlsNKB/im7L1dMlGcCb39rKeg3JKgjxEg6Lltqq2yZTcLUcJowtGJLn12W6tsP+kiD3acJM5Be4p
tceN5IzwfNZJWS+gp//5/kP1WOFW0YKoGbSTzfSAbO9/1fic9KD4vxDqBeogVg550Ud5bMRIN58X
v/d8eIQ42/cKEWuyyVH0tejuRC1YVlaMX3YUxGSLetxZV4ASMDH9NqixniyjrQ+dGSRnsq18LIxE
bMiw5CVBqjNupPtXmEWGlvI0GH6jzfcGNZxdSbp93lfTHBK9JxqAtkXV8f6BoBWAxDO8l/NHp5tM
lj6jBP2Jkdn1DlAznThKu2cUiTUGPvpjjsDwn3FafcJmsluhGrQCtq1+QXwl3Q1oPMdr6znPcaXn
exN1oHiHvd2JRzxAOMgMAHHg273SnFtwTbREtQJ1jmlgYL2jv2FvAkVPNYGbe9cku84rCk6Hbvov
TKqAT4piypjC0wBNe/3E+UtLky8cxvBO+sS4ubqT31HBGnkovQ3y68dDT1B4J8Psr+5gIjlgDwnU
ekanIZII+WB4WZxn3mMoWPByH7VHf2m9e87Q5KtP2Lijssp8suWl986WB8nuOLcX2qlcbgVPJdNY
qjdyBHkji/O1Pkb4wqoxN1qSoQrDwXou3fzXcfjKU3X1Cx3cYh9QGgMjVIQpKNQZ4Ubs3sHEwZ10
TbR+xwWr5BT4AZ5kgSj2NceB8ByuE1s2eSecpMVmMnuASjTq86g+Y9eNvmcRKXKCtQFX70C6h3s/
DHcH8LbczwbbdkEm7q+LYShU/RG5SwhFzpv2ZZVY7mo0Ly4GJoZslgqE/p/zpQPUsOaUdztet2Rn
mtMkF8ldwhulr3Os7qO662dVV0+iyUD/OKyLKw+QjcVnCBD52Bp//C6Aw5TezN76hTWh16QOvbA/
JPro6YB1v9Co/Mt5ndE9e4G8HNBwj0FC/wP9lwNLLh6vybmPzLgW3rARZ1o1YZbjXFwA9Xs/JAei
qBqhQB8OPfNpuzlY5UcLRQkhEZFNnMsp7hXN2gezN+kBkxX+uRHsRNLNAgCikrShSEyOEkCSiFfB
enCep/yxndVaVyADH8/w9GaH+aDkI2ET223hPpYuRHfa2iZTUDUlkF9Tn4l8QAqzCUJuazccXH94
2SGK0LxS1L+T1aB026eYTJzUTd/i2NDov3O/2u+GADgzsygLBHXEAuCWLITgnfVujc1sg99ya9lG
5VdmcJPqxkt2Tqe+dZ6K6TAmlVrPX7FsxWExKmjk/v8hFT4Hdmr65s/SNEMZeML2bCdpa+VJHuI+
uYyuoMz59utuKhKulFKy/DzHlf8N4ig8mVN7EjI/JW7JJ46go3LLTFNl3V3oU8RpkEIG4xZyHPE6
x+K4wYxqH5ShzYPdV+kL+OOcaJy+dFgDCDH9bZ9oOntjhPwTSVM9lh/i78/WftLyNPbyuKjn6jz9
7inopUr10Dzi1SnG5UE83w8z+snXMShlNILIIc8oyFn2HFOM91VghS40D7WK1B+/iCz2GzR1y/vo
8nz9hkL2jvc6m8mDcWCT1BmggdUd7nkyWdvpUUb+D54nS2kYGEpwgQh2Xq7Yf6pCtua97+7Bj2qp
D75mJZAPBbwTuZgmMr5Gdemb/R0/oaLqZxyx2eL6ORhRItkbBd5drUpQGkNTtSJRm+CUD5sYyxFh
FOnBM1AxU9Pf5lSY8w9JsUIp1RfR5Of2dZ/pz5TWRxNR4dOiS6uSWEoaf0Fl0ZKxvQWK7Ul55ZFA
yhfhHh18+dxDQNBol9NQrmvliC8cKzP5Q92ca8pLL0WljTI+lY0tAJ0YIlGjZIrKYQBNN+lzgYD0
1+iePMDuPZKj1eHW/LhJS14t3K7zJXvvbTMUtqYitorQZ9IjIyIR50eySCoegI45i1yzRk8PTE1Z
X4IVcl79szi/33ecHLQk4A2+IkiGULYgEEEWJu73iC5w9/Jv2wIdTbN5y+TBLgnorZDiR69BYovr
hG7s5b5iCUXOiKaOqmnsbGCCCXyEmsDsVw36VLVZQPlCYd26tZt230ibkI+Xp2TTgXw4WmAJXk6+
wJnzaBWx/B3iOL1wimGflIu3RVRZv3ifcUWYQrRNrTLeFFDnv5D7zEHwMyFIIJeHP5j2dfmX4cWY
cgMnWaK4UdZWw0MW6FPPVm2Ufene5lNiaSKNAaE8Ni/V2Sj0v+/fJv9JZeobFik0bD+2T1t7qPF9
Pu1ed8/UjkRNAISKVc/jI0M//DmhzpRchpp05NlMe9w/zCLuM6R0Dbmi3et0G14z+G0ULunmzPKU
AXiJfa4A2P11x/LFhp8RqA/AlqRuY56QJ0fLnA9RcVd5cbLZ5ICRoCEWxt7fDBgUGgeKydkF7wc4
xYBEaPkpQfSCzAC1vmm3jxi6mh2H3T8obSG0SerhelM/17siwLBicxGxUOpxR/JnDWIcSdkShsn7
y4qDzPhRurzbyreuNROByc+wLckqoBZXVrbCqxkPOPNatks8Yvmr+eIxtNs57AhqjI6/mNyZrEkF
h66aEy+y4SlOWCZttMVsE+c4IJzXemJOzhiVrBzGhqZWDCVzG1kc2bAt/fOOtpY04Al9KKGYeudT
oP8IIxtXQXdRHKZGu6X2MOP2D9qCUNPYnZrfPcT0fDfYQqORBiO0Kz7ffxcodc+A7TzccrDGZo5J
EZ2Y+jBZGIJmyLKzfxJR7/glrU/QsOlgMGRIaZEFLe/k3zg+GntdZ1uJw0EQHq0hUrgOj6tmuP5O
zQy55yPYgJbfFqvDtWmGGkzzVQIV0CLI7dOcQht3yCBtGnDs8+AFcBFYbhi89sqG5AfExWHfAJIy
AQjzBr5grS8QpoGROi7ciilutcETlM5TMLuABSgYAw8Dz4Ps0XnUKv20RrHO547zzMA49cpIBs+W
wnYI3nsSj5Ml0FyTQpgCTLR6uaD1iytSc0s0LzgaijyXaAvm2hd6+EPvv12Zq+pSpA3WJe3yrTDB
ngvQlXVe1d0dthp3wPHPOYAMMXjVDeiApMcOvFqLGjfzHMKr0243xCV+4G2tH7WhdzwfC/5DWlmx
oxConMISsEtqSmH2GQLdhtEpE/8eTTnPXPRRekvD4Vtb855Hj38PIOZTTq6otq3VYF2San+/UXO8
QeUcibdunG09M6q0SbcH+CzhVW7gujKC+l6FK07DCZhpyaecer6EC9lk3rzJ04hgHHMR9uppK4B8
tVmFZCdMbcNjHoVvn2KpTwUWE0DnxmnmqbmTNxsJYyvaC8ulUabFOzSlhzKyCgVzjtgvpDqh/mrT
jFgPUYHy0oJEZPPKSK4r6IaXcNmFfOphRygDo/bESO9287ILrc4aB9VGyvdCV5MREITR3rEw9AF/
5yJCjS4z4S9ACQRtn1jOLm+VoIK7dUm51h4nn1K7fD9AB47HGGKpbXXzTU1odxfytZ8cGaKqOaHK
YCRsxScfF4Xqkb7WUZ6z5ivMBGH3bRmqJ8phFCiXGFmZvUY1c+7uW9li8cPHgf3rJBG+YrAmoUuX
F+FPIW2ZtttPJrqKZJspk8MHC+Z7xhXxponVMy7+FxoPMfmrfVg9kAs9+aCXrqPND4jxj+eK0Mc7
ZoBTov8Z77AHHXNbrz6VBH85FHzOSGOGB7RQXiDlgEEkL9rwYEZoqVAZ+6t5hLG3vPf8InowV7nP
4fJBs0eJpmLHVMU2jlVkFOnFl1MmfXi66eA2pseiIVjFN9wRzscnaa0aBD4LLUcx+ABJXROb9Z7X
FELQGR+ELladlAgn5ZVoXMqd4RqOGMyQU98YftQp4sfnLQgrf27gkrwCfDLP133bgnux3EL7NyF3
2thmgpTmwJFLu4n6k2UgHykDytHW6j8nllIHC3VtFrXyWCddWkI6JqI5zGtWivgvgTYmi+/U5qTz
rdu3K8QCi2vavwGY8KBmU3xi+TjS4/eKjslxA/BAA6SSZuVYhf/n3ZN+/TgjIH4UZNrI6eNHFKPB
L+moDVnpaGu9FWDJm5cY4yeeTU34akSWcQWyf0zOSEj1frjohLxZJj9+1Ls3W7JuG0kRBf3bknTu
HQEykSNXqDu/WAF159lRenLI4meVb8MDHwi7TTnxM0dwEmXURijJhFMEFO7QOi75YnN2wKf/+7Fe
EyZhRZ4Ls2rJT9eQTtEMWsExtOJAODFEGL/W+6BHa5xx3rB071fQfZTcXpwecVHtrmuQVB3129Eo
3gYYeqWqLf2IgsAnSSYnNBWWjZwjcon6HX0STj0BKvoOArKNuIkDN37328nFk5rIIGuFNauZ6q07
aZiNbPUor7bHYZaIeCstzBdBgNMYqkydRmuU5mLcszvRk9IAgggfoUyYl7p7sbhkBbQM2GhxuIeP
RGkjE4QSyNCdhKAxcsKqsvsr3LLP/4G3inHhDd6cLUngTBdAWhTdzC0fEDR2YW3zWr6jtjEclq/7
wlq375z7CHSYDuT3ITIX142xGMQG012vXw0ZhadJLu+iWoSltov7oF6Jkl/4YIG+FcrXD/HD9NIB
s2Tv+8yGknKBXf1+2RFFaHXYCfPJwJ8M0N3A7DtLzG0ycmk+9T1bboeQYJeirR/aax14H2F2AcKx
ATFZJpZ9cRkiFs4yfjJeWcSFtNXRuJSwE6wiIw2CWmtvBBUjizEy+QQDNs7fKTx2u98lRwGZaVNm
wrTvIxhk87oIDc/UCal31xczqfG2i+Sz4TgnKe5jWwpmx6mW3eAqc4/kOMRRWwNIuUTmDk3GyE7B
0MdCf5c8pQzkTFBHnahi0VWrpacwXFbVeTlsVblNTki3o3JGkT1CE7sYdfPcK68kExNETIS5bs4i
VZhWTAuNlRHudYzNojLM2NRqmieADHzXYLTkaNHQzf/aj3Qt/ReLVsn5esBiaPQLmsQ1zEPFQXye
W31D96eJEAjDpYbKtItUvYA6ywFzHE530voDIk2gLw5fm82u21HbDnw4jg3pXNLgoaIoiOfnqli8
2+4IAFeMdcathY0h6vS9GFDayHwEEevX4EWWbaaYf60vEMrkGt8W0I3eCMIGVIkI4bY54/sAKO9u
/50Egc6+yyBG8HN33tRhQkAqHKfpFrzKzLZJCBY+J25pJEqq3ONKEdCCJTKkz14eKzVYHQ2qqFSU
rtg941yS6TG716q4urE84n4QVwkjHTzjl2/JtAoKYFuI84FoPWT54oXPhHn6LPB7IJ/Bgu11aRA/
aT5V4NPc6N7+a9LOe2dToGw7XFG+lNtGkKmxaD+674TkEKjsqhtFnnx+sp/x35PoiWPaMZLxkDXC
zBCS4XePyQY2c1BlcDwlfSFSVMeaVsrmI1fZEy1gtaa8yA2IaVq74VveKyoYhPSE3qNPXiJWjOz8
Ii8aq8F44uZ694B218dD+FKgvRsV1zhsTt8tzl9mgbqivD5WHzX1W2IsNNMqdp4uU1iMoyRGSEVs
h7stDV9xrO40mCuuRAikMXVz4XvOBIuBzKKZ5OkypZbhSIp7WqgZunTMTT+0hobzbBzfjC9wPiMq
poWgGbnfq3AMco2caGZ/9rJYpnrQDH8cHVF2vIBe0EDHM9KU54qCgxhg2R0Y3dfsdt3Hycca0hDc
/+EMVKkmuzD5hd+M1GCBUYhPr3V2+w+wsYy96CsXeTkcu5KYF++M0+k5VLnh9OKp64yYqJ68j5ft
tjsBx+0QHSINVsHXHhWItqYWJTXhUcD5Z77XHS+HGyHfeAb7m31CgVYzE2508DLrd1J2yJZ96bKk
hZZR6GGP+F0tcdaGI3wInE8eS+QwOHS95W7XvtHLfLHEMV6cGFENC+FfO5ZqKpCnBRrqfzJa0yw+
SW2AR0PV7nAL6NA3FL7miScnGf4tpATtylVRsHEluCaWbIm8PfuMWWJW/A/qDeAvYZx/CRPJDQIo
EoZNLXLWMUj4XhvdtbLWBziaYvXyMsn/zi9tmZwkUuGWtKE986DsgS2cXqfYvppuk62mRKcVD5ze
VER39+SkTvUUeEyZoUQn8BoVRlLsaV9QqdGihY+F2c5oEo5BnBySjp7qFo6PMIDof69+ajBPwnAX
vuxTg/ue5oB7imO6Wyuf/BPp8byk2fEAqKnAviVLi63pz0+6+FLiUlYAa0gQvFPW23d7lIrrR9P3
xfFBZma/7JeU1c03aNZ4lm4pGFVEMSzckEGAc5TdLj5oLI0pu0qLKOLUWTanqzsCUjDAyqXNsuFk
ItkVUN/aV8usq6CNtYvTiEhuI7o6Qu3rGkKLQnjHKiGxfVpyeBmjK2hq2yCAt+v0f+pWj5cHXqfU
NC/ipcHe+hr+7pPh5MlSgazp+5B653TckQV2+qeCJZPn4RCWqUTF7lZ3MVb9qlVweapAHCodpYgj
KInIa+5NaygqUsm6mEMs1BJtOTOUMMxl6TJOhHnuuaCWs9uxnEIc+I4Wy2JFt898OKFNgpIc7F20
chB4dnvFEuppF+D1HpMgy6drZ01biG1s0+VNqmwwrd5xBRA5vkD+S+ApUSskOx+HOjXiTNp6TcbD
1QsDWhkcv4To4i2vGIhDOaP2doyjydOKRjQGVIyE4Tj5mfIStPPcQPQD8InlPsTbvgOKxkme6YG3
mOlPKlOKRV1k5Zy7HrvXK7pEGbmU3bmSm1DTIm1I56f0wZgyQo3LD/pNCKF3BOtqXkRgURt5monl
OXVwEuhEKVXoHNwunrFnV5qYQl/fA4jz9WiZHPAnmwNatBti6OsT/Bg9AIzZWQio/wMWEdu7aWRb
LqgeG9Z34kTOUxhvnnM43VzicMIP87xvas1tHIN5GeJXAXlpnJSpLuWd+yU9RQP92tamvQe8wyWk
tOgoNlqDNe+Zi0uV5a1J/Q6D3YxYCgOhU355REDKzZuphe1z7CqPUWU727vLRo6RICBfHmQS4jxF
JMkNjr2gXEB5czIHUlgDztTh8d9vrBoqqM7f6DFEHlFDNQVjY8AUY9CSaGDJVY+/NqTZcSo1lmG0
YtcTCECwO0zpM7zWF9GMM6OOn83JTsmgkG4yhyuH+i2d9HsvoEMnK7KUnjbNZqYnEHuKEXaU/3I/
ug9UAMkVcdcOiwIoCkE2gWyLJ9X47kRkJp2QZd36j785KaNgCaHbeaJ/F7V7qwY3sL5SPWx4TYzq
fyFNz3d2gvqpjbUYkP8mtJgt1YaNUmJFd7gHnmWr2y5JUGPXWlPk5z0QQlylE5Y/hfFb0AMk1mlK
2oWARKf05Te6UyIs1EwHOToh2ef8jzRIK753vG67iz+pQJHivwenuavjMYgT2yr7GRpoQvi4VVI0
zFP7No7sfu9VoUjktLurB8vfyhGattZssDeHDRjOuOBG/4FnCTr0kC2al2Ihg6PeXILAEcgzuIND
Cy/oK1AavTuZvCq0l7dpnYAGX/sDxAaRxh1p51aEPE8IWXbuoHYmT/rRzeQ/UeTIKrqTkUuzg3Zr
vdVx3TQmKrSsS+SiDU9qXLwBQUdCV+SLQc0OFccFr014QHfc9RyOgd7Q1Kp8VMPEO+qKN7v6KeG/
X1oitoFSMLMNgihxNORQpKdS8zSBErY2OGAMIYWcPa0cIJaZAPwdXAKOFxE1O8GUrHLQO7KAdzgR
nvPD+MQwDRIgLO4HCpYH+6EFkaRu8EW2KZQ+1O7dsYQ7h6S6PU7x6BoLJxeddJ3ATY8h3rBfPQyg
PvtxgwPdJCCKaED2sDkh/Tty4eUgeJxZfgFoutIje+hU26qthgCAkfxLw5kHUFE7tBwNgN9JDjBu
+l61i8b9NgXCRaCLhKsM2Yw45R6c2Vr08E1/HLzIDGnEBFxY2F0gdxQYlH4sK/QGPa1IW0UObuWr
Zau7Gln0lWWEF08gz73WMuRnbsnLp80/DiNGNuVDencDrnyBAlpi2FfRKON0doBy+6S1MzptJzN+
ONwY4qUkr3pMwYqKyByhWRKr0ZM1+bMYSqn4cuCahcokoW0SUsIKHA2QYPLnboHF6fH8PPeyH6Pi
PZWl6XJFhN2m7vHgAIPE3lZn1td3qMP67xG1W/G26GtUCSH+t7z35StqWICkdcTg2W6ZIyCEH8rm
EtdRifbtDBEHwoDWDN1WLCIB0FGcpRZiDW0Sm/rKnlUVhjZH74lXnPCFEaMPTPzgZvDCiaL1aO3X
qcyZlkadlR8WjrSNjSB7urKd9RKYbNlxQih9tfq8AuWEZEuVXnL3UW9d5fBVO/QlVeQuonanrWai
Uo3dlBnf2B0RHmpwjcgYN1OiPfrBPbUDvTGC2e0MgUVwcmMtrAEQo563dW1gEC9EJxVx/C8LYr42
vsQN4mWwf9D8/GXtbIDnOo8KhVWWcNDdlvbAX3clW9D8Vlxl5t3zX3rK/qQe1Wg8D7kQ3N180Plw
9U8vNXF5/5SilPCZYIdgH3I4PW4G30jnfLTamGFuUTrF6JMXGNopBRTPT/e/1D46lTG8Gi3tdEvv
jRdS73wTyKW8SbbtMp+EMLVW/EiVLsWBvWDJHKyFoG+xBACljTw0UF0hh2GUZCGlr90LZHAdH05Y
Ol/EprgJxbNLZBu1ZcbGvYBaZ8LMiMjNDl7hRbPHbpT9EVZbCpTKUmFthjOmhH3bWsedYL5vbiRK
rV9O3LShMD0S/4Neu8nhLq/geAYChL3g0p4/BPufq435LPjHGau9LlQJmU6c507pjrcMLurT/wGR
AbYi9y6v+Q9hXCdYtz9CP0narhV6gQtQdhzjzji/OPAt34GSTsI4GLFp5Na8X86JKr2IVNrZnyMN
fah2nDGVw+0oBemlzRjklC6RxYom4gc7UbaHoMpgNdfvksDCy6MLHQpnNce5kKtfBgXlS1P59LAM
+zuXUR/vTeRVupK3hMj7uUPbswNZKH08cMTzQqoPPS1PumYU+ygIHQL9qGXodiFa42FXeHQUyYJY
1xiFWpvedMHIWWB+RYrYc6KHf5b3NScMFZnavjctgug7FlXsOjeU6QaKKynUr/QWSDMZ4E+78wvM
MzQqmqXUHqHG+d1MDBPJJQNnX62g/NQhH/DFDW5F2eH/4L4TxhhsaqjBFNH36ivVDGLJcGk/U707
5/kc8wdOE6Lc48GlVOz2qylFJCOV5BTaMqPxK6VXHxanpb9CuRvpTW8KF+OBAD36uRdWNfq7YUZG
Jys72QOJb0bykX/jHBxqxd9Tt7vFMHi8hWrT2FAXu3alyWvSqKyu+FAAT30SV8oxViMaEHTZd8Au
TEKUhvUDvKlddJ6xehHqSftAj0j8v2qtzpQwGxl2ERJLTU/9liSnot4ctEN7sSGzLMPWAnMZtwFj
SJ/zWoGfYqfkc72T3bQbyRiBictBOu0Lz4sESrpiMSHp6nSmosnSFjwZYwX155jViJv8qd/jrs3O
KAxTosQGpQ1wAvWWXvNm1wmw/iBemiY4i6NcB6pFQUp+EPUWY/vyAlosYRgT5z4F+CqoGAhW0Hh3
YhEaUh84p8zjbhvB1q1X6cRT0MyG8mKlD2ynLoMYRkQXSuH4AABXrHT2lzXVkDlx39hBCqnqy9os
qA7w4Fnpl16DtXqhqqC5UdI00M7W9/dkPZlJfv/T6hlec/ttfGLQlofLEJ+zseI8mcCKpYonXkNT
on/4AJ3SDLgjbI6VEEI2zVEBCb4EC79W8YBFLYrtxzdxcR4Cww0+6oB9YKYpWtpK020rPhBy0435
jAJ78c5jQdoLLkwF+5E8+JHuX8F/ShM8eXIPTTUCuTI2Jc5sYWa49F+tAMtd8fBTX0MpDJdGFeaf
DycYBjL/fiKTnpdvAKSzm/NAO63G5Hp2DViJ1w1KPxadGS5+vOvYUGoKN9kaKHLHSErwNH5XsJXo
sM+jIqLBOhl9osrn3sifvds7JtwcTiQNJ5UbA6qJHQiwVU8OiA6p8I2pSva/38xQjaKXwQmUHwZc
v6t6Wfu30NYe7Yk8vI5FQMxSL4bP9tGyWE59dqUZzLyerIxDwB2/WYkd5TBOmyLqyLvltrel5g8q
0EEcWZyYuUjeG5/s9PbwEG3D0GDmuaZ+fidhwhHYkgvHXq1zKXXM4s3cpUzbYZWJcBy9zvgOeZP8
O0f2XnDULI8H3IfHEZNJwY8RN1mDNGSZRav9+vHzY0LAb7r5geQYuKvyjfkm4S2UNXft0MzUo4Uo
G+ioJL/cpasQFjt0zzBoN/WuQVW9hz/ZS1OmHTmOCMlrNmCnv+issM+xyfc034Rzkal2mtofsiFy
q2qkRSpuJIteP6i0YgLiq4mH5TO6wEhcYPU/IyNYrlkLCuHRb3aHi5ko1LQ4wT2JMqMBbRw9DGbX
ukQaH6xWlVF7qVJGFf3m7v7QE0GhM2KIW8MOug5EsiehEeNZUL4IK8xVP8eiorU7ypEv3m/SfnBn
FoKP+q6Hj8Wa1yjDDIdOBWCSMCULgtSxkos1tEr3d++WjkTzXhDna/MtzQrOg5JEuEZRUgyXzBZN
7/s9DoSWEJWqx79phwLEXu199BsN+7I3ocKub92L9Hjql610HJaFtVv8sE2fQzxkPSAla3tz3Lm5
q/1O4AQls6w1ySFRsnCjg5SlVi0WtLYUr3nDgQ1SqhRTplCiGeoT4+W4f7yrrIYQAjjCf13zqlmg
fBvvpw2Mu90cJ3l5odG9U/tlwzRYP7ZZ3rPYykd7K0RnWi2I9bU7EPXPp00Q62YS72NHN/bN8otp
KT+HnZwIQNsn00/lkSKpdbkZENmmxAlzujpqJrOnaNVeMs9irmZxXgVN6WPTao/e3aEmXsmPfFD/
q6sjOHuifTj6DyR8aLKOthS+NQKeAnAFXRVAdHZU8CdacEzZbuZau4/DD9FVmVBYRIsfIn4cpDmp
7MO3A1uSxa2s9UMDgOqrrQ9ohyXTH5j3w55zrzFejJLMKCdejzZMQHK/LETsyB7WsSfKhS1X7TZa
i2q99NMw6znLykIternme3HlP/pG8mckGbSNr1Pj7XvyIn2UOufgUt5GOaHY64K3tH8ve4eM2TKf
7NycEfMsI/7d7d5+amY/Ll8kHRUxJ1ERZN3HhX1pwCgALB2UJsPcgJhuIMiNbUrZx+A0I3tHuX/W
6qLOnLRJhy3hdQtSMGQYiG0HFbpcLpiJY1uXUvun0mNEjfXb4/7z29PDs1k3AqM9QKF8m3tV9rIQ
GpZhKzVOphH1OJzmd3AKUpqwkUPI0dWrq8+8HHpyu08jtAsncUJGYTBpHHDXXkUX87vaVt8dOuWw
eZzjEw/0abX7TiwUh4wo0EIAtZg+rIQAok3aahcj4EXocEEPkda+whBaOtfU8PHQ9XkCT8cSPwFh
q/yv3jerO7o8Lv2e3WgsC5d1Y13HRwQCmqXdyCV4PwYwKaZwYdzWe076BvRuYYZbCsJb2wDDcNZG
drG4Dp9lrF2TM099V8BK3fnCGLRTxV5+1T+t51X/4Cw86i9u8kyj01ZGWis+Of/G781snUnQ2lJn
FcrAJnqIsvWy7/Vr2sZgQgreMjsboSOafyT1tUOudmUpDfQXWHXVQsVaFgvZg8sdn7sAbj2e6u11
YS5jpWq/oVOR3gQKC3YNghVFP34cSu+WEZsagRhNv1YJwew+f2KFoO1htiYldmCSeixhAU/X00u3
mQHYFjiImDG0kHh19DOhwfyDPbdoe+dBJV4g/zRkEPpUGGMRKndow8olhFgyLZmmUsioiFjHSTYr
QrSXtzsuHx2H83kSLYiCicjXMwJGsrxDjYHso/kaHMMaEc0k9Cl4nd2ff1tho9z888emc0VSobN0
oyXXwD72AMcDcJyZtrfvQ0CEeCci/mSB6MiZ9p9ZvAxEYQZIpvbtSQo3Y4EdGoYeZm5z7R7We2kK
cTiA2Fgs87Qhc+URkSfvQeh575CWW/JQoL/jGotlu6BvEBQXykqq04Vk/DmtJggHHRNdQ3Jh+ON7
Lak5HFj1h9nB0oaTm27LwaqrFzTe/zv+/gmx34OHH5cExMCxqoPvmYjK4ZP1bnzj8xr1bhVASPRD
xmy/FCnAgmWDx/9f7N2qT8LvTnBegdlwJvwstpmI/1Ov4vpevSEGuQb/Gz4rUBk3rGpu9eIoKceP
J+NcTMWO75YuU2HEMXGi7hp39+uQp99qvNCR1A8bkYdD78HuzQXhOiYThcP6CnJv5/xeHvE01cnU
hjaoLeTGETQ0B87UWLaEY7vgz8vDWNwQq8MKQaLtXEorJUrPnv7t2oRSFTMdqc0iXG6nxn7/MfJH
HcLZumVBMv/IQVziWSKh/6u/Lv8eiVwr/GTFU+RiBcnexqq0qAo+mlIak+4SgzkXdcNFihjRDBwA
kdtbxcZsqVzvHOj/8BGpIqb7naSLMtLik1Zf5lXfQWBPjqOcL7aNk6rJIQbH3sdWQ7lJ3/zRKE8n
90nvc+WMd8gLGww10FNv+21T6xdtQZ16hitiXphnakl2BiHSgqtgpRS1tcRu//ja2zT4VW4YVWnB
0sHfY9cUT/LhxFYhaHpfU6PZ9Y0Y4JAYSOVnIVGi3/v7cNmuF7dcaDul5+eewYSzxNVR8ttJDMj8
B1WRByxiT6CmLu18cpjabMRy+AOs6spOBJ28qHqC5vfsyFHrasRLnk8Xl/chuYg0MNDWZYkWXrpH
bynDd2QIMCrWLbSFrBTrWdbbdWtGsj7tfp46viDY1gbsAJFa6pWfBe9fo2EQbpytrLdgtTl2R5Yf
sANouO/jln9FBiekeb1gpTyZF+VBNY8SZn8yIEwYLFzkqs0l/NsbsXlZ1BS2b9RjqQGPvm1zx5Ys
YA6LM5G2GqsyVGHX57oHV+tIafWQIaDYIwuyeom4wNPm7Cs5StQTXNmKgcaHH/8ssZtBr5uXWTve
eFXeNzGSGl6rriS1h/ZIjUTngYvFG1JVKbjmNfl6UYT4znLxYa8pNKjef1P0uFOH1slPN4tHyz5/
P8bfs0tuYCeAs3QS6NlCglN3YkXRO43maI0PqHi45+HEEYlyQoFwss7rE1zKO6uZoWS5SoOLLVo3
63TPvlw398BQZaBfMotnJH+fMrMWJskm2z3FNr5OHoTivibmUcWuXcDYfbEY45TXO2I4+HHbCM18
6+/Puv4G/SITDgxuEbQfkpJmM3uo5lQ9yQWcuD1e+08EY7hZGGH6qLYacz4dMPhJeW+CJeZGgsra
gQtv6+DV/JIly6zByese7RMJ+vI8B28FhRGzC6CTELRCyFk0Kvt5khbsoRndOVV1ZZBXjzGYtSOW
sjUqh+hR8q9ujhAPpUj8W5XKBdvRncxMNcJpVd+5go/OUIv7CheFNGI4WhVgJMwz+RvLU5GJSQ4w
a9zSTyVGQdecr6pN34QwJzDq/gGiRqNhqbYvz2/gNrSBrW3z5MddoUc8KyyspwCRyTROQpa10b8E
bV3mNVJpNVaLYTui3audQfRqJo4h57pJsPWyorSiNZNPdn0DwZJ1S2F3TzLdUzHqwyKiKrHLYTr4
dpubaNtw/m4FUkc80wTv16gArh+zMTKGbBHWCm9wneNCWm/OYulsAM+J312df/tMJ2ikzI4MbdUy
bM/GE0FBzwwMJUqOhLq5uLO6jkfA9+1XKWIDKjvOwH8/y0+o+GXklQ5O4lSAcrtSi54dWjUXSvlj
K8m+LGasW32qtWd1lWgLyGGKzzU9GOylb2X24zffh9XhvoxrniUDS8BL+GLRCAXamY6T8JGsf2QO
fj5Ef/3PiITBtRl5Ii6NGMVLgWVQJG5ezT1Pm831bXpAlzz/QEeUQQ58fFWqIgjhOMUXiF4wc/Vv
dOMNSVZJ8cRmdkInpfxPiEB/G0yM7IA+isvWsSA00UDtHQOx6r3S8N41VVvO/+ULDbknU7SXiJgN
DuiNn/qm0MeSEQL9Avd2jko3clcDRnCyuZ2HXZ4E3+NZCpepMNnfb74CvAMXOgI/pjNCjhrYCPeD
ludBIxtLV5Ket8e34N85AxkncK/loZROuQ+TxR6ByWx6Zg8aGnAWUqzypR/ZoB6yHDzHOQCz/sz1
AzcgOR4biTVqT9nL7FLW2hC+REEIMNnDEnccYM9OzGj/mYeDzfeMLg7BoREyj9WBmjLgmbHsg5sW
DBNnrYJUKuVeqqVZJ0djOoBjKUgi2I+oE43h1fJOrBa6WIwz9A9ntNpo6AYFZGaip+rZBkceiCat
pkjKRTLwTyC1PS3vxDIQDiKbc37V9GW5jL9K8QIwd/f90uS/MPZDujbg4Va3At/8rP1uHlfYu2k3
K1eb4CiRlTyIf5wMibEzxG4wK/f+ozXaydzsAeOFjVCiOII0VZARNqhnJEFjyMCgy7dAD+M5A/Ca
B+51Y394ss+Ij+pUkXQWEr9rCTuCeJf19mHqmH76DpIIR4GLWsqPmHZGD3Ir4MMIhVE4ErnFdhx9
N0g9F87NJ0Wx0k2gvSBO/NOGum2Fb7rCh2e9JMGWlw6IiAuYrf8yMY8AsABZsidcE1bsVUYVAMel
FztqQdrsfkliBclqZPJm61ltJt76uqwfStcS1tDkzgsIPHPksMyPJWKIEAPgvO5uwSBB+f66nxRh
HAM0eIFtX/4xxE05XLcXjrWJKrqkL2EI7BBVDbufE8hn4SmnOj+tsa4n6L23ErBhfJn5Lk+xYjHQ
ToCkF4hIfM80OVSuUMnu/4KEEUBFndo8u+rX7RRHtY1yzDLllIL7dI8pbBZfZ2cuV2B+Hibtsrpe
kQ4gqMGKzJEknfXTGePkrhlDpstmErjc9afcQY6gaEV7nxqJMmaX3aRr1PBwtMdi3ilrhgvtwmbl
kVsIKrDx/WQbJlGDO6cOJCRQ3e2PAJNxLPTdzO42Xp4EypRA6q/sN9/yLJP7rrNF/4wT3oqSVYfW
bw1bS26KB6BpkOCiulMVbyiC6E+ovM2UAKI2bOAhzuRsTkB369UrwOD98CSsPPdx4VlEFEb9eJBs
V2kyfxLB50wsVVcVeYezZ2+Zc6dBOEXlTMsCrhS/VucU2q4Ry2GmO+x8WzW2bmYlYZcY0DEKm/df
VqlqlOKVC4y6pUtkEHqX6UoMKjryRFAYuHiOuTG6i5p46JjYPExt8fAzgd8sJ0uAf6jSeg16KzWO
Qizpu1zv6GFDndDKSPTcSCNz+Xvttxw79ZlMdMMrgqbqt563wJi9rSoBSy0Ae/F0Y/N3praCv4cP
EgwAwVD0REyjP7krU8oUBFvIugdcnvTTsspvd7Bk/eykvQI1A/Ve93fMMLWmqLcwdxUTgggGR2/G
bC9vGruK5KVWQCth6sdoKwNOB8tsZn6WXASRHaDKRyojbHD7pgY7opaxePbgtBWkPfUfT/kX4EcW
JfXD1PgRhFeZF+9TRarFWYqdsU9sHGUrQ8M8ga8kttN7C1p7PVgtdusBYMgGh0plWrcZJjWoKAOG
NAnQvsKlVpxm9LsZ0yi5qTwKtqYKSDEItsMZI2hCogI0OocRkYyZKcsh40qUXOCEee6hJBMIJQfm
Oqw9xrj/Y9wWIW8Z+qz1vE1weCmIhfvSP86KYby12gXhRMthqgxsDLk89H/ccTMC8++aUwYQKN8R
pFxHJRoDsSWN4l88n1MZpg86z4hXUMvaVVu7FbqKV9xenlxjfbJnfyBiaEOhXeFMntRgj8XgEF6c
zxbUhCb081RIn9RyIQRHFdlhgH9RVDp21X4ISGelAeDPsId5pbFRQfkWhbkrGq0kQSvm4fq853RM
ko1mTAoXrPtGTGFbG4DOSXCGWfv4kufhhiLrdl5XQDQBKV77TYqgkyu+wukTG6ezOdcan+bH++X3
Su1mbCCloY//N5ogT8cP3zMBx5LsgPjSNp0le5zj5pyzgPbAkNZefCXOXTfMk7WQB8j5Y+FodMxC
mKA9BM1UoKmwng3TwG41Kt7Lp7C3XmmtsmBrFIju4x9LOTNfZbag9XCz85Lh6e+ETbJSkjOvxaIZ
VzNdZbUYXyxbXoTncDMexYYIy+AbzHHi2XbKlhUdB2KxaBI3emUi7YJFSQh1WPBYQIR2oDke103a
uueWFHJRg8dFB+XKA+uikkjj0uLE0WakwblGtc+M5rbETFzgMDkBvLSyxA129iKDrH9CKerLHirz
ApV6bnbJtShos8oiEn7Zyx9rM9NgBWVVJHNdk/unZTnLQeefHOXfg7yo5+Ss7fj86TIj55y/mhbE
YeySfNeg9nVewTAPaZBOXRQejUBQwpN89ihj30TwPBDtACsJA/yy4hS+uDHQEWF2uXebEha9XsdX
Ggjupy4gaSzb4YXX1NJLDg0mwc5Ijsi0SJ2CsET4c5nvZQNA1fm6i6dy9YM63+Dp/k5NTXIdx6zy
MHaDGCfNC+SmKH3I93PY4Zkv4J1emfQi4TGRDtFhBTOK8FUdiUQDSq2wujpwS7iBKzgG0MS08ZUk
aIe6H51FqVaT/9IYXPY5SMAtO/7jiVvU6BX8YmzVWs+3I1PC88k5etuqKV6amEO/x44ec4/g9awL
g/2Q4LK97cZpJj0Lu9B6//1uRmNaBpOi+gTEvvKyUi9rZ9hidlkdJyFfyQM1Wa9ffhk3GkX1jvcf
30I2fQKEZDN45Une1MwBHD4/6y4iap9mfjEBUaYT41YFll1vMNc6fMJax/BNhX5mgBZtDC4SIGe4
SYbxuBevXz5AGHSOijs7QDukntNpygw7wPKh4GIAU6apg672ZXUxqMMwY4gp0uCkQ2B6e+BidQFL
wzQlX+NmmNU9joeRs/U0OjZFmWKmjFGsyJXi5Fb5Lk6rKjibV6/iyXQ/696gYCsuZWKdoXDDSGca
qQ/o7gZyF+D/N108bJ9RvZm3my5/8lLymrhrQ7CWRKB2wUfEXNaflYl6mUs8tWSt178GYNkbczuO
ji7EWlg+27bu446pWMvG9LjHloMUTeWw+6ejj51n4WZepShQgYYjFQCTSx5d1ksvNSlOnbr4iYH9
RkPNQxzQUWsyNRjChv8GK++yAKIRpoTXKbM3yDmmFkuWcT+qlw8yiLxHQZJGkeFQDWwZdD0tMvhp
X3AAOHmSZuRtNU0+jEOJ8tROEpN3rXSopmGBwldzyHqvuLpvs2cC5HUZlFBJw6Vpoa5yfiOGDWL1
FD9q4Xv2imbGw9EfGc9FtAOso5MUx/7EF/fiOc+GS8mhRqadVtIRuBVzPjEwaqGlC2JQpNxTDs15
mZZ/DKMrpDgRHEphMM1e2zx6oqrdpIvoNZwiGONMr1AR5XGBHIzOgjt15w7/TTtDy2FrWhmUzg39
wzznUaH/w3ZjTxSuYk2NXiSdoBdTOb4Ddm2/gMhLIlp3CztXzSb6a7eVqA5XDHG6I8mnzZBe/VAs
0sQhVa1TqaDT/9QcdV9BmD/kcrr9CGgaqel3HVnNJCit/8Vcw15enqQvBZhTGQOYb9eoVkDl+7+N
4c60Au5uUMAN8IzZ5AaEWtEuE0xm6Nbcg0RQYf0Y5vtkyV/HWukwhPC7FDwci7zdwIfZskYS2Uu9
hTKJIoAvhgu/6OdVNtC1rS8kR6jf102rPLfm2suBReYYYh7ylCxCeBDjbx4m76TpZMXEpJ7HrHqc
+Jiqzz0AVVUlUNJ3Ysde68Sk16SeyIljA2sZisChbx3lbbe4CzxS9JeiTgIkWxzJ7hPnel5zEDqn
7t4lcs7grEy/7/FwegamAkBLlyBvBW1zesMoxsK+wi1PpD7HvtSmTW+iqd1z5/1h9ApcVtiuXkEc
aPEmYySqyKKBfB2bcduEhNzHjNkO5HJG0OM8TVl55hIavZNMd+kDTcZNEwaC9jE/DdJmQl2JC7H4
c2wTIWeYti6EKAn7+MX/Aki9+Wu92STGGOtaPs5I6Ph1ceYi+LWHdVVdTRpsm4oMwgeoztpVX7/V
btkau4BVUqTePYc7pCkvHHhakwZOQcGdXPwM2AJ/irRxK1HaHNCk24Akm4BOU+ehrIn0vT6Zw9vx
qGiry4Jn7Xz3O6QV1zJmG5FqXhzseOPs7667yMZtw56oW82lJwTd6QIQpmfS3OzyS6OFEzWrJMyI
nMB3bfmoz5pZlxJi4H/79vdiloOqTqxHE1UEg0WrJ11izfA80cBfnMRq/iD+e9mRG4QjtoXCZ/8S
BWTCbThtwTxzKtKuflw1KyKW5ilrH3ccpHLWJnMHkL42bqqxneDik6uYlxg8JSnBc/HtBSzQtM5f
zLrYCZALUVC1FVyBeiPia5+A/DaSi1dvU+6TIoDOoCT/I19POC6fcHA35VMJIVU+0aFpyVXXLf8h
SVg9N1dlaHRnsKvBp4TaSYcHco5q3QwcAXZp1SBmUMYsfmLq5t6k1I6PHz8jOSFXnq2kyr106zfe
hU0calprCcsULcCnWURp0h8lvBB9ghsBjHmikHslut7tDUTrgzosbnAEyo5ZKy9FY6r/oNF76h8K
7QYOuXANnL6atjqeX5DmYEaLFhTMEYrDGjU0BmQzFNljPoOQMiJnT+ka6CV2OwjMslpNl9YoA9uj
oyLyk9RitxWJFoSFDF+OV4cov/utO8LzMwGheFCTOPYeDyRcLklh6Gqr7TP3q4DH9iyXxawOEBCO
AE8d584gyZV+YHocaAMYbjN6pFkpkK9E5kTdRPDlFT5Htkgv3VeF0hWOGksWSKQybOtduKoI19LO
KxmViKWUpqMqNbajOAu+0h/ufojHkEfqRSvZf9ehhBcUPs7xwYdHL7DdCzKHZbaZOrk8J8zXw4nq
ig3lxd3I4vJMPI6Q+Wiv2IebMlTtZ16x6E5ClL8t5cwobthgNccYgIAQLLWKZPx0WplbErc59WGS
+1DFW7D55Co7F6Sj6jf9OdfLP34Zjw7hRV45eixiSkdbsb5pIJdOoo2DiD5727otF5A6+pF/SBZN
NV5vph04zZ2E+QjaTI7rx2CynDhzJQqtJy4MLxB8MbHA9glDsSJL/qCDYYntN0D1SNu9mkn+Qpkm
nal8ZdFzSGZ5aSdwZfRNSvoVYIi1ra+S6zqLTN+31Fsl/UZnwq5u0onIWMBwuHgjA5lRB3IJDDZQ
HJaSMPz4aDt//oTLBMTRqiSPwATCQBfROJrAx/MHLvkizJxIzIdiziOEQ9nEHguIjqPhdD+eDRvH
SMGhgkp47jg0Va+Y5Y5mFXOyp+giiy6yGE7qBY1BaX5IvRaXsQC0HNALsBYBBEEzHzvTsWU/WkJF
uVCim3ZZuRwFCfiNHU9SfdNLD8MldgRuMeQnYYRlKh8bnbw9azI0esuH3aPXRzAX9KAg67kNXuSK
TkFF3lqd4F8aDnH/5/SJjW8TrKHIKKGQDK4ohNCBHtZCRZqYh6BO+CdKPPAs0ZbzPAuwbi2bkjSV
DeCe2MbwDWYHzFHjR+0v2yeR6zHtTERoKlJiJ56DNuKv3WAUjTpVECPSFNBwuGFnYLOGC62R4CQx
jbp0KpiAvsBJcPBsbZnfLSGFnUJZynx//PVcRqIG7G00PbY9k6yd+5yj7BLalYDaOL5AW9wBscZx
qelxNJkUpDs0I2mpxPlu++uj5BsMeOY7aYcJowJmENqhsgx3iToblHkMnyNxeFmizeTgf9VkeRsz
hjlY1vyjMNRnRbaasXXtKB1/X4C4CNCGZKnKHT/DPJdCXHsIPzu4dsVzOKn+7v3DvzBwBnCuwlYt
VeRGx6dV17GPTf8Bcp5EexTvccKtx9zOuxjMLmWuoZqwNPvkV21hvbFCwd9WtNLqbEpmHU4s4GAM
IQX+TeRD5zX7teFRtxd0kN0BbXMYeP32FXxV4Gy5U89ac2BPGtIwyCbn4HXveUPQdbqVJ/qQ4uh/
sPFd6YWLzXpc2mVkX4lvF+X//Yjx6ZkHRtMxndyC5kE8ORJC9ONiupXgRSN103yjsGbzjRwLwY31
YYO45mwNzeT0zZUobaRm82HlskIjpjlFRUDVFN/KCmtbTxOv0OXTZl4yIPg+NA3KeasvnnsXpTc3
pubrC0RoZmJgOMrJnHzFt38QkLpKcRhiYVw/5QB5mzBCmf86H81O6+niTBfjeeG90LR3LSiQyQ+V
UlnSxKGUZTFo69tWPI0Cl7YWRfqlBk/W2/AQr4CGAlv6nFjKVSBxHASEFJHkioXd+Jd2BpOi7WoJ
H9OwRdF156tWRsvxA42NgpKVGfkBtsGV0Yw2GOxha2pH1Jy01RPiCsUqDo/88DxWsNhH12nKTzbY
I6rdiJ9hrUxj03bDjUAxa0S4Ix75asl/5wIMFEnK/urYKuXmtfwgFvcuw86Zx0YZ563JU9fZIxNK
25I+QAmUxqudRVcJxNw5/ZZnzL3OHr3KlUN2me0TBFdl9jle1QJyUulKrz5Cb+GK6mw2jfnL1kvn
89/ZS3LNh4syjnMNmhZ/wBOitRefRzWk9AlE+lBZCi+MCRcRLmwyJJ6viYGPn35P3u/ZDBnDdUkl
otZ0xubK8GLRRUfVYAFkvNyEard4aDzl1UEGGY36wmjsmwYppvuYkOZMP69Unz4mRpWgIp8RVzTt
VhiLPw/1v1adbVo08Ulv6P8yPimKQebOjEQ1+JclHO8afZFiTJkbMuNlRsLY1cCLcDL3Rlm1eJI9
tbKjhJ3B2SqPlQQC8DsZxcipATHQs6KYmFgN9mz1HaRK1b+f07oAJkhvXyYObtrGInKXtOClbXS3
oW6gXqyVR6sfVI4WeS/7AzTzp07x49QWsShSspfP1CR1l4FGuDGaTSSMdndeGtEQtfG4QZxbu5wl
d1tFNs3Oj92MEoW4fv4eZZhVD/7qTOqRpM/3uc8jD8jRRn5fQ50tk89nHElUfDga79hmvn2ccHbu
Vk8PGpUIW9K2yCgKMAQXtpbybpkzbbzEesfNh020udi/nqeB3g7E5dTh2bS/ymG0J2Y+3+a2epm0
0AIV474XRoFOEfFbiyrSPm5tjCIoXyK2yNPpduNcjJumJ84xpNF8guayQRwR+XadxpPJeggmqVZH
2GrV6QogJ73LzH14vV0FHA3IcBa4EIa67+RYB0n2yljT5G5qSTLEuIxxtGDQ70eVZnsqHFvAD3t6
Tpu8Vxe7S2YcW0U08lV0EXIybkO3BXIbILf3acJRwFX+fxc0bYeauxN2eWbu2KjxvRKpcEhlIIY/
Jp74namXHF1kZlEDgVWz79h2RJD5DQY1B9kCMFPLLFBrMHEi+Pa4wDaPN806vpuGp2lpRFO2phhu
OjVbwRuUdPXO6h8tsj7bxWMCpD5j9Jq0Odmah8PR/02Ij3ICLODdOM0ACa//ine1oW0Gv3zaruhn
6YFX7Q57f/jaD0uv+SVUZ7xV1AMnxwwoKdV6FRAPnFIS6yvFwOfk5IJsd0zOK7KjHuCewdn/X/Vh
WYSAYE1cYj1YZs+JJAjCo1nP9bMeh1YYbbOe2/JcPH8xtOB+nI4Hd+uMAn7xUQ5ae4cpkhdtDwN2
wzfJjnKKHDtzhGHwT2nEBlZyCcVvVVBF5B9woIL9gczPmzI8UK3wFQi+08QFS+i2AFd4KdaEyfPo
lEQtp32N8tbrp6H8TrPTWIe5pJPdM/UPX+eCSVYYWK54XVHXXnmGZdFydAaQ3B29jP9SVp7A6d9g
K3wXYZ6dBMfMimzyNVS68qGLk/Iefw+Tw96vWtEvKfO9Ia9m+zFWL21C+Y3v9ES7UESTz4P/q77d
bkChxy1uXoDq++hKF6C3E8hB3j7s5p7NP9PKRHDwpHRAI3BvFXy3DXDJ+I132FGp9TdrPzo9IVgg
AMe0uSbqfZ+cwq3DqfHcFPKdM821GRjkz20JAww4aVXFyOkC69tIzW4COcHm+A+S8GZMRCWPIoQO
5UHctYWxQCtMHymSi84sv1iJmOz3NtvzdrTjPpn+WzGyXDVrn3Yxz76WM96U0E2m9dysPUJtVC8z
y8UXyumRTDRs8zl3To9WnOklo7fA+Rm7JPOHh9adb4CXr1HNvNZIoSf3LT/joDXesQ4mxgbNgZMc
EPLgv8H8q9xeLaIHZ8JW4zfq7VxpHYTfOJ1cE/95urxfX/ezcB8RSBuf/TUOlTq1LItzsTC1lT5k
v/NWJ76qwBdAOt0/YQWfNu8Yd8dXaemLsdI+7cNORdV6mVRjFPN09ZnsU1mE2BwkjjIa7vwRqq1i
VqDmljC2Jb8AIPikd2P/rt00SVOd2kZ0/gv/K8C/XuLDHU6tMCf3/fYvbX26pas1L3NjIJahaWzz
SPTwKkGp+NulS3MjrMyA+ESB/odDJ5gZ5zJK4TvI6zEwNq40tg2zywaIPe7TQbwzziAR1QL/ozlt
4vHQDoobuz+6sdQlE4GflaV+Yn1HAEt+9jNw3EJTRTIc20uYrKuEwwWjQaM8Buo+gKC9fEkhIvUe
cPt7rY8ZzEjbbe918zpBsIYE8kvGnbs35uequC+pT53wssxsOlzURm2SaA8Rg222pDqu/ck/ewrt
KX2iJVZg4//+871I7fIzf2RdtG5zJhQKiRFwTrD93P++3q4SCPCNjsIVUpnSm6nT10H4DrYNQNH4
ivXDjzEZ5hTg2+CkxgImd+PiYpp7GWUJDrUpA8X81BIDiMU5Ct0cHt7MCCLTouTRauT/Cu516Flz
sTuA/xAmbJDO7/TwG3kl/NVwV3ZAyQ4SFcJUWIRSNtx+EX+rP7PYU3w8M2cUTxaUswuvHI5iTNs6
sJ4ls2A8avbE4njCaUS4XGwHkKwTSXT3Yda+e71oR8g2fXIEU6EJxcQNq+exgbGLE8ctiLQJ7Ggo
cVyseKL/NZyI+wcmhkm7lcTF46RfuKtnC+/Uo+Iq/mAZllTgVD/bGcHT2Cfk8QgRfZztos+TZmdv
OT+S+vUgXVbNUNDcMk/iH/YB05+EDNcCw5gXx9xWgtdnDinbDCZP3blrNowYyN+dgBId9Nj7AAqu
QR+n5DBi8O9OPiGaaZ6K0PZyifPC9kLILreXjzXmHA2uX5Prkxie38ji3QVAqTE3F0O0NCfHbnqJ
2be2gU4b1JkdM5smkRnlffUgb2Kmu+pmC8Ebc+sRyzXV8swC+WJ0mDenkEh9F6iVQLD1IexJxxrj
XecDtBaBEdjNjKd2g8fWFAhHrBLwgY8/Vs9y9qkdmpUSHpIDkonJWD6tO39UlrDZ2RpSajMy0dSI
vD+5tY0EjsCLLc23cpJzXh9bG7A2dfpjT5jlp0v1VCxxXEWFuXwQ4f7KlokvBFnDbe8cqOUXdf+g
FTYsN+M51jzTJK8IedDsjafftOQi4+gfulxaN+GmHXMj4avoMOAq3Tfa4XJaXnECD6/5+foSWW/f
XG04az4h9gAvB9yzIT/117dFpY/g6GIEvjfQGggOpWneVG9gdLZO5tCMOP4c5AiQeNIPnasvuI4j
AKpWCV7sAnCSA8b1kezomrOzUpgSf0vYx+HLGjeux9de+rrT5Fad/QJchaQ6kvX5hp9o1eArnCh3
6Ur3zNSNrP9R0hGcRP+OYpr1HGjGG1cq1VuUiyMFasoXS/weD+nKGNHy0RVhOHVe5YJr2mJ1qQPw
XuVJt8x39aKs7PGagcdLAfuE7HE2zSX5vx+84gsZnTcBuIYVQ9UnmKd6ufCyTeoEBcduL/DX1ic5
Y5P3QHvIzngJDKJD1z5fV5GNAZ93GlmqZ9+CdnZ+cuqsnJsmjJ1uLkefE0ZkBSqljBXJlP3/MNqu
0xr0JlW7fXRw1gRpwfUrSqEo9rRpjWELaLdZGj8XEWkOytFpSg1oZdcJUb9tcFI+5rTsZMTw/oKQ
1QZb6mQ6JS7lRrcTZ7Ikay9TgZ0zLVX6Pt7eM0wKr4YOmhUmGAul6PZlWtaaQrxynwzbqUB8L2NK
40Ym9CKUUgEMeHNo5FP/bbKvbjOoiVgnYW6Tf8UD+KX6OxfNs1qQLTummhbtTtx3DavRx7JWZMQj
sd1nUe1hJ5x0qbwEZguH5HVsYzluhjqIJHKc9c8BbJdiPBTFdNDqYtF4dP2OPsXtjxf/2p/4AgbO
1iuN2mmz5NaienkX0Z5DNCqd0p6ZlvNkAvitRo/J8AfkjNq1uq4nEya7GBfgwv25GZWAWv5DPp4Y
VtXu6HUh29gOLNsMDjkjslNmDS0jJURz9M1gxWH/umL8RqD4w6TfogZ1ghWvcBAT0aWez4yFAzIR
uWRkbXBIVBaI9lEc6JJTd0NK9b6ELDhiEIkNnUl4cQ623zlqLg4qpInV5qBQpiolzDQRhF9lw/ON
VtWd6ZDrCqQGlOHhvuaiBKpm5HGsFMGw7j0Om4J98Dg2wzbsKNg4QYkyCt/9eZf03La+c9hgFasf
QVdleaGC/Qef0ACtlOvBARjwF6Sh6mWZNc+8wuPaBOiRYwINVRNb54wMrKsPYtDwhYWiG1VSAEYp
WenRMmZOx90uQRHVkKk6htxsCanins+IH3iHMQfEQ56vDFlE1uIGp23term92Oxv4AeySS5fMWkD
aSJYDSMqFofnrLRM0ME24VfhgebUVMFkU3/839TwJAWLCeqCSEfI4lgVsjL8foy/UPQfnoFVlo8K
S1SkKJSVlhYh683Max47VhNJlQasYxEd2nvih8LkeQIAe9KsF1QhwR3p9Lw64lBHS6pwfYm8nTMU
CcUCVlFyvdixLPkv6MrLnCHCTFuyE3+LgGysGXSDi/hnbv6/WHmgX0xs+evLUc9PcmZ3muP5PhC2
daJ0mKB6nCn+x7ePT6FtmoZvzeXSm0sEqVWoPtQweau901nUXwd/PeLKa9Harm2HtknbFe6Dy3gC
CGeppJ03fLUvjZ9qF0Zp76efKTJkx5XCcmgdBtPTD2dpVg9zeRCG5MO2ag5f/WghkMScBTChvxKd
uEa611Sf2zZ26QCKqPNIW5gTVYTFzs6dAJbIYeVJsKiIth+UzBBfw+E0vL36oGVOdbtluUTgYp7V
ZtMm17f0c7y3BfAPbD8RQTszlS+AVUX1UwOjEBmeZC19SnFye6HMkmAKpaEQNzVlN7WsamhY+aCO
UaoBCeWUb0Cm2OjAUzMuX2pAC3tI1zYhXR7Pmnq/Pt3CwYetke+1KSBRj7+7CbLVma145UkhekS0
lj6ZMbdY7wz+Z3uLgahvvCB0T8Puaq0STtsUoN8aIwrWg6TCdL+6uD9IET3D75me4PKCxq1hQDN9
IyDW/8ReJ2vJnJga9V1+36fZvZbX1gxKRv20c2jjivE6Sgzq3qVOS2lKpi5XcFdyOS2i1+/oj7H8
hu99VlOHjIrdrroNVJXf/V5lQWWuHN8+hHGAZkJa8rMqEyQpEd6C2mOhBCdacu/7r9kwrgTgojn/
pVTyBdEUntI33/qO/MW0FJ/v7nyNcpUlQOnGPxVXj94Grox/bvLfpLlMzAfthtamJ0oDKdxZEt0r
NeoeobXi7WBG+yHqGCinORQKL9bVvsju4Jf18AcRu2jMkAY1ND3LY4Z7SMIQwsDAYeyeD+YNk9LH
nE24xJfTEXWXfa005TNGupdvxEeYdNHXpW1eI+iET3t8PnxUm3/7PKwdfa19yNqXE1Vwaqnb5+cU
Er4CPwtba/Rzb4oeMVL3DxHl4F80vLqmr1PHcaiJ9c6CqZqpxPk06cGCXiewKPW++7ut0JI2rw9C
mekpwxMBR9EpXfUgyv5GzFkgYfX2I01EnthDYokzZTXyBUbZwLEHaa/cCULoBsa2Mg2IuGJbEXf+
fxFGD95Qr7c7qPM53koAoCXLiu8r8O3AUxnkB1UFKzB3jgeNDZ0MuXZnAMCnEnCOSmEQRHnvOED6
HfZPwPsyPJlWg+EnqfO4QD2NpiveygHOT+aNd8GmJ8DwLci9gNWXHCxyHopN1ah4SxnA4kXan8mx
d1PukxBrVMygpy1nTm/v7i8PTdyNNfVEmeWoy/969fWEDtd0KVQgkRvGyYJcwCPltJr5cHKGeigO
cFUKvqb5MOQLHTrIzFj1WY9j/Bm5GUXFpaYBzu6QHA4+UwQqEMS0S3Ik70OmA4aVjrNJ/Y4zg3/h
Tm9oWwyxJSpTfe33ZZu5/2UOdDe2BCiW4Jw9bLzssKmVOrsVhLnYPFXDu7KHeYbqXkl42TUNB8tV
4wizy/h6VPU+z+uH6M6JTf5zuU03E/itkWQSClbJc7GRwefuKZpQ2cfIB4qgh30t4ItKP54TFRDE
HB3Y+ly2nJvLTQLXATyb1MigLQesc2sm+XkfQVzw+XuEGpATsnHJKlRQAVkrr2AFdUq7sUolxmO/
V3ocmKTkTvWcfbqBlAE2P4JT7sNkFhDasrji2Jc/3dk4EglHUiC55Pye/2sD/SoR4F/X4Bz5/k6E
1o41TBs2pVF9p4Kf3+GGCrdQOD6WMsoeFHj4BFikfEfggFHHLmTOVMn6PslqejWjGyTzEF37Zmgf
y9V2sVNAoCRSU8iajDcRAZ1w3WjiuVh+5fRgGeTp89zJ+LoQrWsUmN6fo8rizYeTQ9pp7hIK0SIM
43HVR+MmulJYpte7GmeUKl+rn8XEDfCgV/TQGcSANWqPXxCmBBmWq0ocKhcQ6goS2rwdVXR//Pdz
qqxYniv5AHW13UsYhNjZYms2zgVihDy5rVTagTXoekGhFT5bqb69D0vDb9IDjCIVo9nM1M4qoIUG
WCCCew0q/Gl6pFwx1d3aD7Zy4N+PptLulhqV5qaAHPCcqa+ufigkybyR9wRYP/lIpTva9BJJroZa
Nw5bqU74lVsdhazaZhoYrZf7sNJJXRUvATzkbuFWd2r+S9PU8otKN4ZaPFIVVjULQXaCTg97zEL8
uYcOAIh1L7NLvMWUM9aQHUcCqgkdkHccTKMtlY2MqaZahMUiyvatJuG6oiZGUS/s3URBTmDGc85/
5PkoG99P5/HVme3MlM1WJ9etfFybjKvQh2hQzlHEyei5MmwJSyiU5V0EPSNqgjCD2GARyV90l0LI
tWOEB+bvZUMODREdkngUI4lVE4JVuwOQs2T6CFsR8VzpVVHZzEP9Y/fpnQIN0pNW3FERx1Pj/huM
AtmhkZoCtFWdA19E63XNCNMQ17DP0wmZu26n51YrY34vBFTSsutL1em+0o9AqLBqsIK6fPYtnyVl
KusAeB1wI0lCkYtTY8JvSLbxvQtvkxtzib7qKeBh+pfPi4spnFA+hCi+fxuPlvKfRipJVFoHsm94
Ojbrzd0CmMKYrkQIZ8GCnAYr/8j6LAOLA9UkfHpWy+29k1sqyH5yfgx/p+bi2kIjfaHCK2f0onfM
97RZiLndwlVyN7kBWNKDeX3JazOzaZMxG5K+DhQzWvrKofTXjQjvd6MlsvxaUaWYKvccIKZX6GRb
82ydyWw2wX9ufOLvQmb90BwA5fObd6K/ncRTE2N7ogQNesQsMuxJ02+GlB0AydY3Mm6dN6rJIbQW
xGIPYjxxHu83OTh5RLUcdo0IyZ0AeOauGD1uw9owygmwEWfpw9aSiNB3Ulg6N4lmgp6u1r/OgJ3E
f78Z9tpY6QeHwlQlIsT/F2ZFdzfbWww5MgF8RgpCw8otbPC3vCYELCu5v/8kVk69xUXx9unFFcS2
cV+wBiYQS8MuaPaLljRTjC/+rnb2HVOVUyyev5bjKAvFjtXKWgImMsGxXOjxrmvjbERpsLqQQnzM
6PEeEhVlPKCZm8bPhHJWNnv9BETyP1h4eYvWUkIelMFOKaPG8IPqv5dLv5YS9pWjyvyhRN8PqylT
oDhSoYraGDNluYxa9tw/cJCfEv26T+EbhqEu33nd75XH+LTSYewAq46OVpUGzq9eB+UmPxOcMO1a
vpaEBZ61PrZ+yI8HaY/zKkHc5nhviPMPg9sX6G1GfhrGLPtBSGbAWwHVOdd9klJlomrBhdtSh5hI
SL/kadc+mLeKIZ15iU7f3aTlC3+YpuUg37ULFjmpm3m/+ed8TkKcmJr081uqMljbAP/xNgRgYJa5
59BMuayRmJoNSy+BwUiAVUdLWKRpuK3G9B6jRFRyqMELGdJ0XIzQS4huOmwVex7F4ypcFcU97Wpb
bfkadzAudWU7RuQeQ7NA6fIj0WVKQAjDVhXGJliB3MKF/QkFhSpl8vuGmPqobdXdLsWoiwtjoTrN
7MuO98wTipzfJVlEdXwtSl4Wig2TXHGj2NebdwAG5gpWWPfvG9VsQKu+2yzbmv+0ydU1yCyA0r7M
nCqAyaIEm2oBHLISHmTTd4vGjSVWcqBnVboIH/15PtPBw13B6q16sGoM+qibjwUoScYyOi4XMfQa
FpjJTAQeeFJ15IvLS9umX+hopxIfheGTy83nl2KXt5wMhjqWxHeSw0VOwGFVlEHJ5TehMd3dA4F+
tGzW9/KB47cc1fJkc/2IL0FFG9UEZUMYr9H8u/OoAgq5BdPRAVKbzrNRbzVEP4P3zvPqghdT/1j3
/XrUL4H5yf3KZ+wH6NeUelySP+2GIFeItYAE/j2q7FMoMWjrMSyAeZYlcEilNEqZ2ubhz+Tr0uIj
BtIKtLSZezjtc3/4MFRisBYS/aG2l+7+LX6pWxkyW9v5a+hALqwDImY/+QmMVynFrX5DexvnRExm
VvGeDu8u5E+XfHcYBrbcRWmGM8cvYlH+p9XCEmjsrUzqVa0kVCTBzBPZ1ZaoA0KDxgwaJDeEHS4C
95x4Q56nlhcBCkRp70sYXtRu4MoN/GZVygzRTzGiHTAKK5vvL+WK/0rceWKj6kMZVHzn+Hppo7wJ
FXz5WabTiTUAwUEqztB8fuha36UzlG1VsxzZlr7UZrEn0XKmlPgOw7RVh0nAD0dSb5QpK5WZBzHO
HVFaYWSXNTMoZ0/yj6Jbd9S1qkjBEu7XKmHLmSDpOY4RdQtH9HzTFK+B3RpWp6hzEatTAfoLdvzh
DQPOqOZNrwITP2y63V3kHR57SSofGg9sr8nhv3Orh4xaMfgZmS6/aywwA+9quNqd6TNFlLfTSyO5
zgvftEWRo2sgldVsEPGrkfPm6qLgv/B7lzBNWpPPNFmsBM8VcRuNVZulZDsMBoio/mV+YX+5oe8A
Eqa9fAt6QhhqMRPznIqZJRuREiwKAuGJtUNPBvlLj5s+366dKXlqBJvv9jEFrspOKYaxgzest6BY
mTtVhG5GpU7GT52cSvnr9ZnTNX8meEsVq6qkHP9/YJ/tX0Xi3GE1q719Qtj+DjjGDmqdhMX1GhIl
V9G/r4bybfQ6pGkclBVc1egszL0ivjFDABwrw5iD3swz6hWcjiZfUPPV27NUXOkj3RHQgjfdTWYK
SYo9kwdR5UuEwWxi4L1YAXzQOE8dp0kVA/N+JY0GITjrrCL/HGb7SRQQhU6Bpgk4cPXE6lCq46Y0
z8v0Noq2tS/lKqt/G5SYNxU+Bm0cip26hCz9fOHn0P4h0B5dEHkhz0j0qoJPLRs27bq6TvGz/Z4j
45yQkYBOWY0bHBt19wpY8pJ06oLRd8K1hd+FjDfVlsLyvYH+jNeDG973UJiMrdrV4v4xHwH3rc4K
QK0dAeSm8ub4c9AtUGgj0EJuoON2Ms0q018BShDwZMcpT4ZVe3urjzEc4lwAUF9UWllEFHOCDzzS
61WaBQfynI2H0HivXUcdMrafd/FJSDmTDPFVfjjxoTc974X54O/b5nG6W32vgWCF9xwoqQQKZfrU
d82aklvrB/hl0n+inOSr6pTbV5U8nEV2bgjDUMkewDRDO5EtdvAW6W8sqv1NpUS+85FJY/SO+rgv
SvOBFwgwCU7CQaBwiLRBE0swVoGZz/aZoQqNYQFuPM7DAG09uHvS+QBzR1MaZ7MZF312RJXrZwj5
ThyIeffZTFX/frD8USRc/IFkw3wRt4rE5KtreyMSbI4r3xz+xaEOpcCFMOoXzC5Eu1XDffZVN/4I
W2x+AEbR72niWUANcBz+ncEZeLvPIRejUYfILrmoUvnUx+mKiPNPoP/+uOaLFhpPAdcGSxrywAct
cMXEtZut5zdJo1cRhVHL723/e65TP8aj66uFg6Y9FlTyoEJ6O0TSkLd0Aw48vERmbgH9jONYhH3M
Da2nNyOHqV9oH5Mir5tdsnWqcdtMcIKX31rRvt3RvcCduoOdxYsFasxXv9gx7AJfmeQF5H4Bri+w
iB/cx9xmgf0MIXfEDp4ArWKbxuYqy82u8YJvDgVZJ1qrfL5gCrKvSDaQwkDIvCoG+l35IYZMYiJX
aEtL3Ah3WNfDnHEfEHUELI4Nl0SlSUva4ul/NCWo+VvHatLy1T9jRlEGOmahBqYSSc6iXLAt7Ewv
J+E5lrVmPm/FYiyrBFAWzz7GZjBsZBNtSMu/Z7on448xXwyF+te6Kj+5pvt2F99gcyzJH2i9Rxp/
vTM6cWgL+vrwdfpxf8idirk/2Dd+CS+shNQHbqrjpgVDelSkdCtACyVIiswwXWA6hv6bpatkdY4s
bS+KvHbmSp/ycJWllvOFLcWId8/7Bh1K7R+8T5U5+r4Q1QcHkjHLfU4twPWjwBNyTv+SOsvoEUzV
I54Pue6xG6pLE+OUZZ39bA5BgiwpdJWmOKckIvse89HVePw8zx2YRXDchyYpikzsjhBoDYS1Ck5D
oyAf63gAXeiBzsfX65l6D9AjWntheeIfKrhYGsC0+KEtGtR0f96I5pOR7eMetpNfiPYkx2W3hUQD
LLp/7e8yC7rBNKKsJBlqEeM6uAoZZ0iw2XhWUwdcHuluO6xeIvQHzR7tCGmmWhr08hOuCxW9sOaZ
CtLLVpKOT5OnShHnyJxArcQAAhKdvBNnvyt8eAWFF4sDlkFH0eBYtvj9l8mublm9Lt1XE1c9eBx4
8UfJ7A9diOZSmP1VCX5sVeidxOgqIouhGgQRFb7n6TkB9ZDwKlShjmiZbkxOF0Q1x3p9w81SccbB
lEUqj8bSbekLVyploE1zBeU1AvAEDpVHC5aAbMB2Mg8Y8HVXEfPFqGnv3zoyg8VPRzDYglT6cQia
L1RB8JvzDiLWOqZBQjrxgmISiNqPyerL8uCoGu4AXwco+qRnbvnQGbu/Kuj6c5oJTWGPsJYmT2a/
yzO5TwS5sh6EAJukTRp8qHLGpfWGQpf8YYQMS6Xi/hCrle/GgLjBRav1RpzsiY1cOR8hw7SWq1SO
I5PH2p2qrNKhJtTo2Q+p3z0AdWS6ozg4eMAQWBxnTfZ+6U5Wp+WYV3mp2N5AKhfMffaRYOlIV30E
fk2/6tWcQ/xChEwQFlnAyHYKFxd8zOQCYGvmI033fbuUa0Hx5RkByaLJkU0WlDMOwUfxd+sAX3i3
ee9kSK1BP+QbhtFJPHPYsuv20p8tqFIEK1kq6hBsqDoUS1BVvYWiEDdbS67AvXxAj9swwHnfUUvf
SBq9ZTV0Tw8zuqoShlLB1cBUDHhsNEf2/h0UjGmK3wkYypdh4kFrPDXaM0K5KnoOqcFPqnBq8fJ/
BoDzk0786XKppOjDDkUfhAueRtjtoePOoe4fLYQ7HL4hF+wHXDj8eSqZhhjvvhdDGJcld9sH0KKR
CfugNfu86XJH0qAxkHwAvOPnCJMLZNbUO7ierKM+eSzqdqfWtXFAxcntfmrpYzInEthLsNZutIyC
Ad/kV37Q8C/1Yq6Gj1tfWEvdYnhy5+nzTSqJdD9tAMWf94ZScSWVQwBSpsPTikIkQj9Q3OUbKjCR
M1PNIrKV4uLiSfLen7+enoZvqO8UpGDkd/26UX8VR/ucpE5cuqgBcdKqEMRNGpydV5YasDQXqV4R
dmGiwQvk7c5tV7IdnmyJPxun4iAzG3xSXWqZnAq8txvM5KwTwiPr9YBxZEXSP2+6Z6qbKpM4OJZJ
uJydE9Fo5/heEwh0goyl6hVo6wc1u55WFTXjOAF5oDnvgZjh6PRGOmZEchtAKqd2nepki+rujdWk
CUEg2C3mo8M/aZG0Hg2FLyxu5HZtPMFkIpW88UHEAnxEI7AnsN5UYGSnWRfLsKEfYUwCMU7K+oV3
6ujtpmmCBjG5E/WP2EiufBXhAhO3CE+rNo/XDDcS+MXWe8JbIzMtGOjrRHB9utI7/00H0eI1yGYu
OlejbS8n650B/LHr6niefzcCOWjyOAr9HNaQiBSytEu+ggQobt6qdZBC7CrMc4dLeIXvz6fsqbiR
0UsJup3+qVFzJ4h1ojz3OWNJosOITjDu99D0EolcxhYh/cnIXN+1meNLr4vAO5er4hxzDY6Qr7Uq
BfKzXIri17FM7WXZoPgVvL42OTfVewNCy5CJmV1V7jqCLKzSi/3qB7Cigbqk/h9Y3MxJOMDgcDEm
tafKtum7M2vZB/OD8KbxrQxWCE/7MMn/W2kYXlFfXvUMWLqI90zL5RclRDQ33yS+ug3KQ3QrVgYu
immIJWMLKHnkqV5iJRgdnAMiJXokh2CkicOnmMJ/ZXmsyppXf4izbHRG/uLzABj89/a3nwmGjwRF
GaWtAkcNvMx19tUyhaTZl9nknEmUQKyxNIcWSBaZ1/EgA6cqSDj93UvpzBMzFYeGe76R5qr90pdS
FNxAQtsYTPeW/u3RmzBGE5FJcNsW1nnULKJXYQzqIAITgxnkU4DaZKWle9Lm/N+3z/tQ7yCDnWFM
0w+XJ8QBYSy/dfSg1FJQzre6Z987KXjKJin+r69J123+zs/IjN9/Ut9D0Ro2LKRMpjNGVDq6q//r
VAZK/3XgtjpVkLzVf21nZFN8Kc8Hh8Rg8xnkkdWpL3mdp3P7LElv0J2Gmin69/Peup3PTjp5Q/0M
YhuE0X1qdcKQqPzffDnUhlpOIhli0wuHuLIL+MbVZIB3gRYFRTzdZ5xcVsT7IUE/XirWXX4kGX6P
JbTKMrZZuP4XrkJigkcMHP5cC+96/nmV8+9xB7PVmI/bcUalu483DDCEJBxh8GnEMQFX3IpByEje
4VJTia1qolUIbtbEfwBeDr99tPKbkHme2Ek4n7GHhA1SKAgW/EPnEHLVwWYAAu9F3VvDkmLW0B/D
smOqcEYhO63JWCD5r9+ufTeDMYjtzIFybSmMDjvS2d/hFNzoGUvKdwebWsoNnpE6xXKJC2kvVeO6
BcmmIxIgRsQjKOOBhiZetEPBl8oBfLO1pJq3kiiWEwMtDCKmWPRaSybv2iieNEbWKS7QFDdwfJwk
/1TnlMU13US25iZcwL/8/baq95YBPz1HOEeWGHq+MWt2vCKczGBTE4bKi8TP2bt1aJeLc6LAfshR
S3D/DiVpg62S7bAmg1bz3PQA9xD0T9kBhGFsfQ8A6AgmMJ02QXajHsmeCsDTSkLFl6rBNFqrjTLM
Zxq+76FqjhTCslZ6gxbZK9CRzJOnE5jDcCZ015kE/B3Zwe0rlkDnVo2tdwJKdz8imwTyHZyhPb1k
IQIvyZaH9uc8uXm6w83XluJMfnyoKcf51zi1CW5GfszePVdrKiYwvL00gZtlrxMFNMjzrFldGFF0
qCmmeNrSlND6iK4NNkpsCLISkYt8PBW7kcq/LdDV4jMYnvmuKWlV7MgwMV3G4fdDsl7eZ++wUGnq
doRIa5XP4S0FiD0sJ0kj+4h/UYAzTP1jsBt5iUokGrzquxND+YdxRkKsUfGA1+BtH/R9I2G81cNb
oYZlCTBHxwfsyU6M/ANzGkJLVKVwWI9yMQOuzdH6+7L/I63+66eogcNvPR5KlVzTuOAuJ3uU6LCe
m7ciJ1gRMl7ZWT9xE+Zr6ZWOL6tihmOMBa9h+DuX7jCfVbVKFYgQvNyRFIWCNauhe+pFjMxIyejC
HkDOy9/F3smbub5O2IzTeOQ8/scajVmLXoJ7LGcaIRulxJTEyYl4gWBs8fswyYS46rKzr2uxb72d
nW9The29nrJUidIQ5BM1doVqhylNsKFFo/dPNrU0hJjB6MxgKMy7opjBg0706AfdbN0CMoQOt8Ey
t5c0cxjYPZJpJvOPP6AzOowqotqh1uweWoPlGk/T0gXzKkm4ed1dX559Qtf0SGlDt/xcibRNkT5N
sIN5WGL26uTVBpOghBzGwSv5zP5Mj4td9lL10Pdzh09ZH3BvCgnZcm0EMt57vtwcYfpb/93OMV5y
IpxoR0mKNzDCN5jW83Xk9ZCvGHIluUBlcAHe3SY1sgivcsnbdgNc7F3CccSv61y5vX2hJEM/fLM3
uUUaEV9m3iH4dc+5KoAwqIAubHwWxMkEoC0Gbysc4rU2Xh0qM57mrUZx77cBe0JNsL88ATlHp9Ls
FxuQWkqqSE0Y87e9nJwCVVQbfqA3gNu/b8ixEQOvnN1akz+oz6br45ZGkkMs7fSEooRZleRw+sXi
nK8axPsxhFzdfCGnaSGmJx/+TsW15R67EDPgHuTI6Q1nF3ZcLqivYqp4m2Y6FAj87FUwzZiI5+a6
R/Bn4tayfy5vyExsz37fM+f98T3+gH9V1l01ulMpHKZgs5mLYE7uVsfai6/CgL7r8EUsjWF3tqia
h99LFm1q/0oenJ06+vOBks64v1nKzZVkGz6CoOOLaXGhW0AdHUNX4bGeQHbB5Wv16spXaRmsXI71
buCnNlpCH81lVoQT8ZVTUihBnV2sJnkIAAfK5mcLd1fQJyMQkKQQ/0FKobEYjuBP74UG4JtKIBki
nNC2zZsJWKp6y1CSW2eGKUZYxyqklenKxYiUjOysVMihEQdjlcFZqimFtfMk74ShJSEewG3lpAzP
FMIAXd2kCTPklowJ0OHeJL6zQaoDwFQDnsE9pBtQDQ0c/fkVEHyaznCoG05R2GkymfvhmlElMX0x
z7OJwvoZZaUo/CW7nwsvHtbl2TtapAtBLHK38y6Gk+dKtyWk304trX9NOZz/hYESnL1L+lG7iGld
RJdgH4fdvUVEONFGKh27WHLQxieIvF3Op1Joz956D1XO5XgbePyKVrQ2vrpnkyW/5NKy5VfC7zwd
j5TjwkVXmReHEy/dcNefPteoJgaJIY4/IRCod5nBIYFusJzOxGKMm68fhG8xskDLRk6qXpQm3P5c
DH22DsV5zvMG3sAIBCT8NwleNca+cYlptCzPTKUPFatn3WpaptVYtmG1Ny6ucDK7fy45IvEYXxoV
4bA3rm17xyf/Y31TNcK/GgmFHn9uyysDz+Y61COk/PKPOTW7gvuJjBkGfvu3k/HpkdmgqQhzCoNf
WLKMWnQ945WibydX17esEt5n6kHttadMXTDDpGcMTSILrcVfZzPgmHzYy6UJF456MctowwskUBYe
c81n8dgdjoG+8d4UaFbK8PBYGd/2jJGFbasLGjdkKDib3ACSrgZT5hh0olnHxSL2GPLVuEZzoaiL
NZF/l2Vumx76iidwxVVGoUbAXnCx/O27A+oKqeWZJjwTrpvYYuEpX42Ce+UxeRKzUP6d8I8A+zm8
if9MVbE8LwSY0a1zxOGj1Jxeuu90ezJQgphONM8qQzTfmRHhmUDUdhwWgYS2cSnJHTUnOllx+L7r
Hg119MTtp+ZnrWMjAEk9SFeTvH2rEWjPcVxMqT0gvl4L5sa1d0t39cpWETit8IEJLLb4hur8OkoX
uh6KF4cl9f1FWqRZm5ljhjoK2KAU1XRdYXZ+v9JGr2LB98imIEfpLuAvnlICQUS6SflUoGRtBCK8
jEgoRb8zLh5q8rTxL/DPCRMf52KONG5iTvQ//gItl5mNFjp+kBaJkuYWCx/p/q1jtdyE/zvrSoLP
PW8pW6wc1Oj0aWZL2Mr2UJQXWzrSDXYYXj67uCdpRKcL/wtz50SqC4VRcvvKxNILw6p3KGPyo8O1
LrFt13v102olY62maZZuBoR1nysKZ987c2X2XOhLeSjQnO242XWM++KFSapYvQF7mApW5A5EEmek
cQcQXvC3JCFnc1TGgE+lu5ZS7VuqZ3Oab1QcxxvKITfLtrpC48BtymiIfXM6nzahzRriL17Gck5h
F/VWqfZwNnjcA0qFKfmmzNpHetRWZ93aNksar63fYx1FZy6nQfSFzXnv21SYjGL2Zf2N9EAiByU9
s7rm0elQj0A6lYcTl6X/5pAf1yolMHKx/Y5YaK6XfU35OpEWtfVauqqc6ORwbStGKVLo9S1Mv90l
uPWFZgKc9CeFHi1750f7jFVVEC/B4nWwDMYmTv6hHPpHXO9TyuvEYEaCo+Grl0BTSNEKueYPV+t+
pbM4gh+c0NZ8CFKAPIDyF5lj6xb+N+ogVzypeHwbaDyxGrWdx7pyFtSxv/bSp+IOw1c7q0hcTxI2
4TYLTrZuMmNvBbj2m07Foof8Nvf9e/lICWpbHzSu0qCGgYtqJ1/SEhx6zagmAfEb4xAHaXmqiKNE
2ai1EWC1zUVzMnlCKIkf4xTn8swRSW4jZMm/zFxY1zuH5Dig0j9F2ZxCuLkNQu3AQ8tT/GWpgJzU
Pq7t2O9Dmp+KHBZ6S/cgncqIOS32gcx+5VaVYabCQY8XNR6eI99R1S/2I0SxWZLvCIsMkCYxtuvl
JLDWBoYoVz5Yc31jVIFuOEfCQKUKJ/B7i14EIjLVeGItnniW3CF0qEdYsr3hChNPpzo9sKp+rLn9
Bv4rXzzuXqFjwSlcAL1t8/3S3TCbiIzz/MIlY3Y+Ykq5pxsTw7VZbb3iS/Kr9RzGnwzz70rO0S5p
HtDRR1YbNtdj3Q2gfYqlvbHMVxDYsJwfPZoPQfg2X7ppxD2KpU6Gs2+j3+L0Zhnet/oq9TIPpqjz
xyWp1B0Bk/4qMznckBJyBQOxavCGsxEUuvQ1WstQwK+sZV//t2BPE69zx6wGchWmOzsctc4M68Cz
m5Kp0q9vyhDSNAHSB70R66nLXPj+98FFAGyLTptpfiJoD4b9Bw0xBiofTRS4R3L4sf3HSwWXgXVs
TKTuiwG42xRmCWQHP2+B16QQwLOGx+92x/uFtnCzQwEIqYyxWg502A2epOePaq+cfoOFBHRrFmwp
zBLpw+JEQFimJjr2ZoeFf6w/t2f5t7UoKrWU6V/SDzeMkBTBzNyEZ9Ls5jl9lYhOeVZMMejStXTH
oD1Q5Y1mP6IHz5fQPjjGCwwq+T8nxwzmtVXqoAJ4HiQe+B+7Tvrj4vf8BF735tViap4ahOFsW/0F
ylndtKmh9e0e7TmUi0yb45+AAG/3f1+5jvl9SxmkPX1WXuOu9wmwdQq4OI1/X8IJ12+ljNLDtDyI
a7atxYBhg5KyBwjHicuAAoIwteCQnmAs9anuKrLZZi26EN5DBz95EtrCMfl/RzvJNl36YOOkzMCv
LRRBVWknKkvy0asRCtAj4W6VHOGoBfLN733laL3HzMXfKIcmXB2H5fNMww6bWTWRSXh5NviyZVBj
vXEnUgQdbW96InmvvAKa8PltO1rX3FQXG4f6bKYm6LJP8nOosIBLTIOwZCCsuMDub/bIxmARGXqw
DvRY4tQrE1sb7uceWx7JLGcqq0jyGb5BDb6x48ktpX263gBUTwJLr5aUE7shhCnTpSUR8Zc/qq72
H6JD0NJjqNBvsnnt2n7Tjg9kfn6G842Ux/lVXQm/3XWWQklxTHh/dukHBHM06+DcEsHNTR8hBEn4
6iD5ko9OteY8F+B1+qOj42JNInrhaf909tBPz9Ja0AsA6DdaRcBFgYntlvvfIiZn2oewri44LCEh
tthlgtjPjd8C+9qdJHUwuvE4/H995vyP6ByTh1jKoYwlaogLyRcGxWhTIAKoyCbiwk8UbSG7/I3M
qAqfyKUI4qxzopS8VmW7KIOv1+H6Od3e/etCj8jOLTuGoDDXbtQS8s9bFOsNTO0QADniiZ7q7Hix
hVn4y5OvXqEuPtgQQDXA3R4Ko5E1pj2nsOEyN8/kDfKX49VeZCmbmWgHdzKazAA8+pL0n7wY8yGO
EvqjrW/uB7818gSsd3FfuVPZQDmMyVolo6bUUyYE7y82nF5CXqDWdXv8ijgKQ3wHbB27tYkFzj79
qRLQRLGlr4gDZZwbjZznOWbJ6HBjoDgT2ewB+RdjzKg5zf+Xg73kACJu4yGpv/SqYJb/IwOg4ldy
EfVi/gyGIbwNAHK8monzoPcN/gNYx/cYqKGrbvIutkSwxUP6tkMbz6X9AFGhfvNREQMd0jTRwrwW
VfFVNsh3MciQcFfmRKvR6bgK6r3ltvKb+VlPrdscBrfmhoy9yeIVXLsJLYilof05MJ7GxwHG6d56
0/LdBY3TFQS6EwkVY7+/F6ZuMcJyNR+ophWzk0tPKpYaPTdtRD+ZU20fwuxu8xApMYmxFP/OM4zG
2fah1mc97Fg9oWNTe96a1Eo+t5DFYlTSnPUilyVC3KFteyhRQ1eZTA1uREB53+CCZrGcDSsV/CJv
A3lwgSXiycUAP5ACe/9tZm40hVFe+dyPcpyZBfh6QBtcrlSKVX3MmdeL3MtCqbRSQxA+4UZCq1rA
vbGtk/ZL1UQsLuZDpEIUKwZZzqDQNbe6x8yH2hSe1QTv2+ooLMyN0vuZjw9ZKwuf39x8HvyjpoQa
3V5Q4MM/DYlqTUbBsDMh4MBmMTAkEBeTB/AqV7+/e5UkMmYxUG7zQkgV0zkCv2TiZmexM0UHu1yD
4wLUlm6u4RSQk7ZL0YOQozvNy663vi61ZPw2m2tOCpKHviARlStnyTPqDEWCYfMwGerJSYa3aae5
k0JpSzwCtfjU5g8hau7FO1+7YjMgOAGZWztakJOrZgKaBUOaP1NV9HA3uN8EDpdF2tVbUimu6Xlq
g1TgRbFTW7STGs5MtzvS8lyoI1WpY9mN19OVIF/4NEb8vD2V73HWb4IC4vl+N/XNaaTocfJHN+zf
+2YXIzlNxPAcZFtgN3WmCF/rT9pMfmtXzv0TVmPHKpxG/kGy6S2y9cHIKY33wmNMBielqVOIzzRy
+AFRzNb4sjE4+4C6ZeeErHWBuhb/a5XnpzCRwdJ8V1b8fWR9FHRdaIQFi20OJVzuSGo1s3+KIsLf
JwDjVSXk/LYdISmpnCinkthsXW7lekxld0jScl4y3YXb31AlBIypQwlExZXVoOjzDRKacfouqFFT
wiu9wSYYe1lpSQLvXzUWDlhbOCPqjksT2lHjtv7qICNIgQj7IbH5PWy/OWYDyaodmdbjfPP4Qbr+
E1kOts0y1J32TUo4kO1YQP4sJ4gsBe9wals6E46QvxnFJ1euBXUqjm/B+EtV8eCA+s7KrV0EYd1e
DhqprcoGDj/YGN3pROPDE35tZFvqnPzXEmaaH3YEt+zcwdwnNfRfYKBPxjwl9PKLm9gvBcO9Mhx7
OAYIHXJuCX87wrVYS3cQZL6elC/3+FHygAW1tuYapT3NzkLcRNx1sRAOgLyNEdbXcwJy8UnjeaMI
cTZAMj8Jnxm9RVVLBX1IbF0up3P0lxhbEorPxUmi0RPRqztQqqKwMnDCz8DdIp/XNr03vfBiqtZo
JphXqTn2T6iSLL9TDDsiS6OuxmwiCtlC87J0+cR4hgg6FVPilfnxxS6tng+M8j4axSZz4gCb0vff
RTK0CyFjwLlbozwnnTRWL0cr2bqXQacMVPO5EqT9qSDixr+U8EG9cyGxBSbzI2WT9vI3q4g1UtCR
u439G67yPqgG7nWLLO7wVN4x6NtvZakXu6KBfkAX7VnHQCMhm7n7Yv59t00Up2bshlJ7BpXFo45c
fT1vCAQKdvfnB9RTgHfaP7T4WFpyBgeB4y+9BjQqJbF108IuX1KSUleIdkc6jaNQmvmJwy/sO0Wa
AXIpDrh9DeaREOlqqPbsB0yhUiePNZQwvw0p9W8QNE8N3OsGfbPf2LRlLc/f+XpZWPXypdEAk2Xb
/p3LrBo24j5We+olHyHB2R6SwKj6ewjKYz8znGBOZ8rvLQRNnVvYXTYkMLothIa8zebg9fVS+81p
MDpgyjH/v3wdFvqwz3NUKfzdMEOckOybSBDaNiIZiaTLnRO0ePFX/OQgKHNDIZD1dArq1+yreQrj
xHbYQ8YrjUDXZiwuM28pLtBwHTY/zXGvznTNrJBPxDwFHaTdXeKCN4xG8lpOWT4BnoF8o+9C+1yL
tu+HgW5tYrTFdSI1b+0M+FYTH9RD2a8xKgSz+JX5o1sr8qwyfbuNUVTpjftolzs9DQ0AxAHUwKqH
wNxKJYmrgLztmK+njQ+rGLlDzcwgbH+IANgJRp91xNFoIlwsa0cuJyME6N1/3ZcZpglLKw6VWUhq
v3+Ik/N6gwTh044PPk7h2aee/ndxmLhAn26/yk0wglCY6b2AJDukkhHt2+0Z5PffvU7qsouBetEh
qWlQdiPfMpmj7jaSC1ae01+hD/0Q4jjxBRLXX2nZgEWTRFbgWq5uMwTgOqWmV+t6iKKbowYpVBPU
mPH7fDrs2bmUDm/R1rT7ROd9PNJZZf5tGpvCss/s4hUFexToBw8wfRcc9UcMGQs00f3TeSrenqin
sescnO827TX0DQchSuYfyJDQFAZ/3kV7PARMBdjhlKqTDiGwrTiJt71KEZqrhn+7gRIq72Z2Mr7S
CJRFlKmtFEgYEIh0GfAvStrsY3R63ib9khr/rUQuF0xPvDa5D5/dVjlKYdIokMRX9CM+eHrgOlDE
YnsLh1UVRRjNms/O7uwfZldpNC/OPpp5VsGf/oAgTlbRDnOaXfCNrW8ZLb2wsK3uXIVkaeXZaQ3q
NaGTFUjohd1W4oE07QV6hIMDSZ6RdYHGqzqkc7R7WwUN1YRVVvYl0paS1sjDLeCV4Pq0xfpoS/X8
d1gcQ3U7XAeKQRRec6IggpcP9d47AoQgyw3g9AT/0C1zVZ4yUc+ljNbOHF8Jjt+RWliNUczrbixD
eyXx8SM9/TNK2FASVJkZQu3x5H/0r6YcfQ2Qby8EK8G5LFJlLGPGZOStyWfY1hN88y4ZzCH4l4bc
vSCveySxoyYIpimGnro1zZd7wCCt8VxPKf6LDUF3i7tR3CSKrRgjerxbJq8/QSLPvBnDxw+KubLK
TB4OHlYxZiIkagarGNKak7EFTZZfw3w2FN/Cg+Zu6RTWvP3GounpwiEWEQm8pOTmSgfREH2AZ7+Y
wPoWb5cXVTlLQEde+t8DIC9aWt9XCUPYoMGAA6Wa7FRJkX9fMLueQQyTXHSMNUz4huCExuamf0rR
ItdhcsaapJqQiN9kU2Hkcr3ir8Qhow7g0CkARVcSNR5Agq8Fhh97yxZS80B1i175tpIi5HlSbQIc
hBva0gmL2g9BONVnDZTtjxLwW1mc/kRIlJY2EvFeb0MIO24zUXtDTILYmz3uqoMfG0llEz1WCLTv
yFJ59miLBD+PGkRIJfA34kb2bgFospo4qn4z4Apqfedy5H1Mpfd4HrSYSpLm57BVfE8h6COy35cH
wwiR54sas6pPUtG9wK9YDzaV9mQgTp23fml+qpgBEdm6JsEGcvPxeSYozVwANNoi4sx/Sz6Apx0B
6IASpa6woaq3p3kLG4jJa3qEGBC0f3NIGHNbhfNRfhbJ1hd61Nf2mikoWEzgnrpaoB3pkBaLNlGF
eWu5L9nqN7VtxSk/Vy6i+/+E3tC+b2NrhEaZ18MU6Iq4jEJ8GbpxAN3IhDGP3zZYN39ExX93TiOK
sSIEiETd1SLjTSl+3Zq19cfMrTwGIjx5MHIuoyc6h77qA59QbxrqY96SDQvM7x2BabJkWXKFqKp9
jS3iXNJt8Ux25pmlrRZx+ISvXm4zmQHWaza9Xbftja94KXdK7DEv7WEOE+RUg3t/JPNFJECdOE6l
2ZoLDMW++Tmt/+MYTt52ZDRaVPezZC9rHdYJjCg1B2HkobYyylRwFFbicLzgkrkD/o7cwMuU/snz
nHOnSVNk/mp3yj89ua739wz9ELtAigu4J2ZJDyg/22/RcoRNs587U7YGwqvm+h0PnclnUYyvsVMe
qvNQBT/I+4NZ8xVOmXpQxSvOtJCf6mUam/MjRrlKZ+D5rDDFhXoQXrlj0KKLuI9KnazYXa6QU7Da
PC6ueBCeDHvt1ZhtHnPX0bdRzpBUJT3wcuCl/aL02p39BdUL6ZZ041grt75fjCRu6drLc2fKu0bv
PgBHrs+lRd6oZhBSgSifvT00V+zUvgSDkvIT5bkQfSoV68hNe2Wvmpv1jtYEpbkdLBD+LpFnE8f0
ME8O7KZ8vT9V99xgj6sXWUr8d3Eq64xinS4PV/fPjYy1HZds+huNXnd5g9ht48X3S8glPPr4/jw+
1XvVonGvTnmPjeIXS2yo/NMhEfI+vpY+DSARfvnZzlm4pIcO00xGDKmy/lM7g/Iq71/ygldt7amv
Q/Z+diC9iCEHhLvfYTTvG8iBu0+n6MddJ+KDntXeAbMTRCXnjt96bp9YkLHq5a4unWXKPQHsftgj
9E8Aaqnydy2SSXthESm+DAYwj9Ih/IFdOkDxeY8Ncg1dLwFdQzxjdIFXawqHD12Vsk/ayt9rI8Bt
i+uXZG+OsDZrwTncuZhfkzmsCAI6zwK0jWiabynOM+FbsXVimteBdD+NfbcJvINHCxVQtGSgk3+e
HTjbRHiMJ9Lfimf47i6xwL2EwfM0ovQmspNeCKV7A7dJEz4GdetTH0K9ZZElSFwiuEx01jXSJarS
jGzMn8xHT/YcpRghGWcv4a7OMUzxWC3KpJRrOtwA6TVCBBUX3PwaVySgXam7S3Z5UqJfVreW8y2l
pQsj+SfWF7HgkMknqGvFxfjUgzx8m/TYjCuhl5V+Ah52rg0VoT0ZIDubdk+8wMopagdLLGAkObZO
WPAYVuu/izFzP7P1h/qJpTTbFdPrb47pY7gWlzIn8L0FuNEEBbC7ri2hlC48uSq3xWwiUk18LkBa
4IiBSnK3v96f40ap5Ti055JFoZ662mVEUQkGtyODFk4wR+rF/NF8d4+8APslHJenQXPjCm6IJHWx
PkPg00dPM0XeAdeeIlreeJu5PbtNqk8Fh88BW9g3fMXoHRrnhF8rfMGxT8n/Q6uwHLGRbdkN0thw
yL5Q9VVjw5ApJJDVeC/sTfSz5aScs1TYmBj4VPLO+8gxLvZXzumPeLWuZwuuQEqN0ZWRzTbM86iI
AJa7Ll7uaFhSolAnYU9Agv5xI/Js4/MESZcdcw4WI5YJjUyXOoOr5wOmXz4Sfk2q9uiVR2XgwDNS
PRIFUEaw4T9wN2nIOmPmyJhKqIDNCOPLl2yAsMXyaeelFBsbBGDc0lWNWEPI1I6HmiWT8V6N62Nk
XzO3Yuj6ZjgECncD6vLy+5JnD1pvQKztMMHWZANjg8yN24Yl3GvYb9yhWcoUNURZtASbFU5YWLJO
+ITozY9vNZP9t8Dk0TCShF+4WJn0fW1hfc6HMXeEldFoIwBQJprox/HQCDSbdN4xCzxXR2YcJ1mj
CSp0N3XHiWXrA+dHSojvhCTl71nXwoQNcoGuHb7pC/RXhBweTli0Kq+LMBUaXRj125yOLQIhszrB
hBbZ6b10AMdFEEEqebfN5cdgNkqmZIb0hQbeKHZUJ/FYJSkolXw6vMotyjiEwiaELtgo9SYR/TVY
bG9U2iJCor9Q9sJGojso4GtUJ7AvEYcaJoAoZ09fN8R7nYmpGjBhkO0VKppZ+maC++uOXqJoEIQz
GZg1n7f9aumC/u5zproskhHOQyeBZSV6lP2AUHfWVix0ET3V+DW0LnDQfcTczSxeGZB0iQZUe7ci
t44erd88jV0L5RFPY1NBm5ToLNRgCPkY6C6Nh5rMsuGcRH7HPL3BnF6u3BQ+fA4gh2P0kD95ae5K
3o35SZYxMFDomsopdz4eiervUp2NNskijNnogmw+aL9g3Jx62llxnPntIghDL8D+a3zSkaX+XCF3
1yrRvtjv3r6/zG3tB4ptGk3Vz8ZZogVqtB4Q0/FEeC26AwutqLsoMh3dCMKscQq6sByIH7mZJbYR
9en12n5HXBaji4x+xWAf31tp/7Dc0k44rzhXYifcJVwr4Wh8x4owATodqSRceJKgn8MTp6FoMi21
hU8OgMS71m2IZKb/pFi4C9h33PNhBG68HxasoqR0M6jPX70ADqNykzAi6L1ctE2REmzexiydg07V
/VwbxXtpcgQuUwUzWIpyomg5CMZu0mFDqMysadG1GAmlKvNldvwUj3MRmOW69GZZWIJVwlB8uZ31
Gxd1k1ml4BNMQoIK3wtcNJYGkHYvkPe8BDvU/m5okkn+aArrS/T0RQQxG4PrHXwlNVNUPvQiueBv
wYXwU145X/cINY29rvzN1XVQk5u1eP3WpPVoyCNfiNnTKrRAjEu3BbhfVG4j+4/QrX61qZ2cKOp2
fyCBC6Ak8+C/b2Ayujxg8x3nHGLFPuedeP/bUQ94wmSaO2C2KMbgzG/eWdhSiDo8iMj4SGlauYC2
Utf1vsAN2hxwYvnyo1vAYz10ugAEA31k+isvvJ+YiZB4oMDMrudXsWym6u0AQoi7N3YCqziDJIjC
m7YqaCSkMDkkYAh+nYx0jEZX4J/341XJhY5fD1l3dHnyiK9uPCouKMbw6xWOWVMCM0i6N2l1XN3h
TcDX2ztE/j8Ye+A2EdMtGiwhEuEUyvuaEK5MXv6tNLv/wx0NZK062BH5d1KAzt67Xg+gMuu9zx/Q
0BrfLMV4ciPqMtLeSPWED+rpqQKZK1damNSER1PXFlwtTLOt5pSI7SKqovXpIqzq8qO2kZowOXEI
XZj0gAJ4LXsk/lM/Ji/dSvwOlRN55544zJ2oeJ0XENLzBmxeUrNqTnO2mimJAd5JPih4aTypbIYt
9B9brd0BXyx5xTEsQhCNK8yIWIZ+cR8Il+NeVfIOdqzUs36/Oo4ZeZ8kVVGZ1qV2Y5fv9y1xG2li
tGue4Y0x9d4oLOe8W8uoqYKT+llL5DXUN04eEi0zCkLDM4LWFG5jKLfQGCyN0UhAkVslUmfmlpcd
dt5QtmrwyTT+4wc8zk2cOMWGhMhu08ui/B1Cx8agaSSDr1VDq6dYNSvYrDxThvT8n2gSm0Lhu0n5
ollvaoQ8PpakFgOo4556zn33xKQHlwxBIIILQoKauwliz/ccz1k3cK6/qdbe/hxK64T95vJPI77N
qNWxL5pVnw8Xxak7Nzo3WgUUN+3FTdPk7hHkoY/uhXC9jDeCNunQNeEhDFPI60fYR7Yp3ZuSukSW
lAheKgysEPAB39w+IYLXGXDFciZ4gUMhdH0zybKWpfZ6lnlFqP2puj3uwq/SUJ2csgKkk3qMY0zm
Z7FDHYqGbZrjCHlxbbeVNVFfOHfILq2GAWgwhDH+3vOaTfPOsGFpRALADRKRT+f8felRR8ybBayY
a6JUkZW4YqTvZS+ETvupkHirQm9d98prK3MVlw/MxxujMe5VR9FIO1pBtTqDQ6M+AgwP+ao15f28
Vw4L30ExUIllCb0lJN3lf9FVPIBseQOH4JKzm1kWstO/NmOyxm679hkae89nr0QgO9eevID6Mx3k
Jv1ppvTVn1NKLI26RyCfAN/f/EdIjNztbBe+D/QlRqPQ9azfA3kRV6dVxa06fC8DcDZrteRZTG5M
UH78yynIY2WXn0oBEYOrWczPIUGFPmf7thW5hgHTgfFeA1I7QNWzgkUEc5ItuRq2RuTK9yqulFh8
NbvdGj5hegc4QxzdDAj4dSwBbTFirRu8VWrwhvCMPiar9SHvt38Cw1kehLBpTxkX7Jn7GLLmkOdH
EAkv81u0nmgGNhiVkEKQN7wjD97pCUVrRlTse2F2QZn6UFW/FCmfBQaRwfaWafSyMMOCekknYoU5
YFr2I5KB5eBJepw6/WmWmA44delYVi9RIMV4Ajk1tyZNjkzzRboItJWJZQencDpwcremYHKk3Xff
bVwsdXVwBD2hzhKAcOSg11hZ/XqMry8XKeVoZ1d3QXfZZDERwwAVxg1ghvWTuYxWnEsP4sIsPSBW
wqXMNp67fWrBMwMmmvUH/yzVKYGfFy6i/ymbsPFegcP+Gg8rIR/AcEwgbTXdoljkg6UqKw2yJguE
1/nt7jhFBypfS5q+fQMK+AdhbfiEF7zeADTFefwnHm3Wiuo8cqHlwGam7VbdcEa3jFGjGQgSOHeE
pnyu/ya+K40zjM4HeN/adtZzsP4HBayXFpFfj+vRIp03aMhDBmNnbqkv1l42GWJtaATokU/Fmpyx
tMuioaBUxR6ubnlf0GMrcai/eITkODqQ7ODDUtOMvvf9RMejI84OBPzAbfr/6sgjcI8I2leYH795
BRuiBuW4klfnB3rQukZDTh2MI4pndPQg2fq+xTA5nD9N53J1S5hEGr4/b5JZUoGEV842PKaNojKF
koe7F00gFgvom5Z/68fmZQ3ouC8J//lKsgsKYkx0D2cTL0sMIbMOE4yni12mlaabtCX2FugKwEbO
l8JBkPntGwvMSMFkM/Jx8gv5vE4ZJb616w1uUrU1RHXVaEf0Lx2qy5R/YHSPKtgWxs/Lk36Fndpf
oOrNuiIWxquiEuwG1zYQvHS0R4id5hK7SeYlpZ5Cv3FBoFT6leH5bFRHmwbQCbArW2LyS36+sQwf
nmrJnAhFoJuyGfm4qtQ5whySBbPrsORxZOTqOwrSmz6yBoFHlxI3wJUXdHWXpYGyfQKPrqhsG1XF
s/bZBW90hkLH+Zc8R/wrSOJkkaSfcVZrfcKEwuh3K867hMBnLhzUmZMrguWG3j9noo1OOG7iQwUD
xq4EWR10ZEKcMvkI1I1l51G3s72yxbD1A9wBvanPPuVkYucoJbuwipBDS4YXqv7jmHxWHRU1/9y1
0XtiKzfvIXmgpu+ntwGfblg4kHaRAs/xxxlQjlCYVHG0MDmy+8/XXZVSAnHUkbQ4xfHNh1jzMizY
hr+WdZCAnDpEdkDxZG1O0RmYNymlJ1nLg8z1IY+njruIyDZk86H/lBqIiRIZGf3ZLCowdcULpsl3
PtCdVE+dXRPtEgHQSs7ztUd+WvWknRyoX/EBv8C+JHXT+QZUD/ZphR2r/gpQYfZeZ78b0wD7QOTW
Mx9cpczxwj23DtIqrst0f6zFSYddl1TkP/48UjK3afHMvY/7/Qy4QLAmW5Iv9H/MrPC6JvwnX460
vx6LIj4cFja9rh8EVu6Qs5ZUxoKPvGuPV8Y2AT57vYv95j5MQJ+vZQtWFmwRO5bDXxjvsBOftBWy
80epchZQbLo0uqJVLW6PK2L19Y2etYsQloCvGoDKJiM3K88GxPFpfPJspIfwcT6ZbdgszZPB5/tO
nvAIXSRoiHbDjKa0m8+Y/0vj8LbiU9MZr7RlVC4MSd1fH683k2iAv76+2pdJAR2G0b96PoIQ7SqX
JiyTDDJm9jYX2MN8k6cGWJVAkjss2mlkU11iaQmwfThnIQrsfOeRI0jR0cLdpJxWYxyphwVSyXL2
OH9JNvS2o/G1D4d9kUuBc3aRBw0yF1RHUxrD4I+pDeqXjSSv29/Jp+8PorXAWv8cgNptPerQ6in9
YDRhiRTDWbs72oRBwl6j5l6AJPxfcaXyP2FMnfJ02+0lvWQt8wPLkgApBe1BSnXiKKTCFif1Tp28
3DEwkWKB1r7tlvkhLKw5qsAusRWYN6g7vJxTMlGYftBS8Q9qZdNiUCJZkMPpPil3YT4BuI38vimb
G3WpbldJyleXQhpW2gJVIAHvQ5YuIYq+zSK/AIUFXaQ0xwAblZ/sQm2D3oXQa0wEc212EHWO8SEw
WznG9J9llDwps7NCzdKLNw+CbRFW+HmARu1BjGAgK5UKk6kqSdUdgRm1LUfsysVM02Rs5+dkzHph
l7MeL8nxHZ9V84EEtLPy96+e7mwGPF/vJ9VqqklPblOuoIsdafYjw4t4dxx50vwA9HhY2OGLMgZH
O1AYYK5r7HoXA5HiP4PXwH8PglZYZXY70wzDjL14nDsre9zppbeS8HGPm1Ny+gMajNK7AFAwGhYo
PZmfCIus3NDhbqLDXAzFALidd1gnUUfjDSVINeM3o8brtwyOTuqJETFzc0SJNPDrylxT9+4AvKOv
CM7fagwxkGj80yl7XF0O9a2a0GQIDFwqEIUXR48yT17q75hu4z1HLe2YVdaaor76bQE9xlL9d4nQ
jhwSCEq6ItUH/9MCO7mLLnMg+0RNQVbJQb8g/e6/+6AjVBp8OcsUKGAWzCNPikrKl61GcVP7tZQ3
ARq1xtWwM3Gms+QYqCMRGMmQK52GK76ZNjYTVNKLPDVie9F02lDf+I+mIfRerryT/+1QZulL43ij
1QfGrqIoKKkoIW5wPupvTjw+QGOZOYFsqrNtQo6RVigNx3X9sVIfAUgeAKSAqq/Tk1bWOYzLicK6
Z9xRUTwUz/pOfjqDptXn8FZ/yzku1w3pMG5HmZwDKwnHeFgCT9TrH/kY0stcbiS5PStPgAAC+yUd
8JLV9+tNmvVb9tiorvCN1xtNdr4anZtKfKKjphXgqxrbYDMES+8lNGm7pLZVrdjLEp9d/cYQEAi7
NeYyKrJfmyh3O3CQBDMIc5U7ADJPZE8C0hj6pyu5NrpsV1INY3WFTsQ6vkpqycMMfp+GDjYNkHst
LNcKc9zbfhYYoEpmw1Dg0PD6BvvkQKM5fXbTWWXXqmXwutKNzTS/ECxh7oe/Cs2ScYsJgvWRiWrT
M+sAdJYpT3/+LVO/6pmrhP1gfurLq7hDdaJnNIXWAvH4MQCOy5mE3ug5X9Y9IQy3t5mDlvQBuiFS
CvBlF7O9Pqmn4KgIRkTI93SSLUCdHB4+18T8ElL7D/2w0HyUkMm+UKaYKJW+7/YhUlqRFpgBDRV9
aHn1lLMfwuc8udCeGrLOJtfx6K9BUa4bRtGdKONqy89LfcQxwWGgFJ/Nqdlio3oPYg/yzez+h5fH
1DLrHWplswnE8TZziyMnn275BTaRGexg0FZBVWcR6yOEQWbuzU2hcG7PgVZFA7VkzlW5Ms1t5t/u
HEdqxIjAIaW9g69HzX+4vtd/EPJLaqKGKgXnO4YmwHOI+qKTT/rE+2AiGcWH1ZrzIpP/6G5qULC+
mP2SPfgxp0jsDjaS5T/Kz7H4MTHNlq0aDe2bv0ljnebj8WEFe2N4OXL0x2eYUpXBaJRIGrIOCeZT
xpx5AlzjsrqwvRY8eNCNyjlA+Kq8LHKYb9JFpo5A5VrwUdaCNTM7BKEVyqg+qDdRFPJrdbGl6Y4T
ybJQ0tQ+5QBcP7nK0Y1zJDumAijPtEUNyndSBZYKLDUhzfwwBfj/D0qJwHhTku/TiQIKT8oEqdAK
sjSNt9Np0fDf8nFMTFSsc+0whlDN0pTjqY0I3Ki1N8Qxm5RIhEY5ZkT+zfWbl94hBTlk0Hw7vQSa
bpJff8n1RR+igUZa5NA5Dr0atSLAUt6id7iuWLF8o8Yf6BAiRXXgv/GOtBV7TqPveGsDYdjYvnvK
9+Nhdkb3ZrAWh6DP/5RxiALn7mL824/ekaptZ0UXC0TgFUFst5vbGhduCe4GP8iQM2ufscP+r5yu
ehOUsGk/d/hwnm4P0FTUmBYgXi6y16x8bv7saj7z05PD/PZBwOlVQf7TTVf0ZumxL9Dww7+iPm5e
pINldf3mD5bj3JddE1+qo5Zu08pfBDxeWuQ0PR34uAs88zaFoCDEZfLJb2KLesByYThk3zBbCE1T
1msDr5/cL9HsD6DwjjXH+tRFyx9NvsIegj/ahMQgkf681h15lUKWysqlb+nLPTfClklD1uDtwEA1
fOiw7W8eiSOdrFt+PQcIsD4jDoQaVRrkel/Del7sAo5rP4bed59V4tCPD7L/jsstuSy2QexyoECa
vUwjhs4+LmIgBJKoptxSo/3uSVcymgOWCvwDwTXYmpV63gNeHskHHEH/hBuNg81l2L6HWuXIBI0B
HCZSCt4fA7yu93kBcaVD22GDTG8BW8aAV5w8U7lyabihgaEPO6iW3WICcoTPI/5KpGn6IwvMoy1e
O5XO1UTtPcVrCy/xPzTa4U+Y82gQpLz+mMqaP+kD1ECvySFLjiNwdQOK6Po5SC6yJogoxUvrLCaT
tFP/i3pkkHDvXO8uquCq37JyT3ZxCBXms3ik1oJI/CwZhYGwt0CmsR4GGW3BjctKAaDZ9SoBOflg
877oFrQ5WrnR6SuZ5SAymZP5aq49OjknUmNGzi2q4KrrCoE+EbuwL03kUcyEeaEcOJmB47rXMBnM
IMpRijiBew9st3uhhf26dSDhVTiIbu1PAnLRSfLTOAxSDLGJjir7AtwCre23Tu/kvc//s3sQfmlJ
QOBYuG1pdqxmwpUMHN96USAbEIfNUbJRpKAYj1Nh1nxD06QDjhfW9pLc9kz3yR7+wI3x/6TiabB4
B1+Q+lSRg37Bmq6ndNi5WEE3VG7eKtA7rhET77Cc00HIbaGj5pwmJ2VedYQWDqNjHo1HiNXBXYLT
JVS1DAnNOnFwTNHTdP9Pj0ZADFmQT9vOJEzSQ5YfmMhjsXgDy+2YX4FY81VOThuWppa2o2kD/GEU
2MLTOY9re/hL+WJeIx9Ma26+bkFp+OI6if1OxDFSmn097jMdiK8x8455OGRpAMgcjbQ4WFlvDJpa
z2nN9txYRAJS17khXSHuFBaT/iWOijOs5DCf829lzbttHQxwOOA4ZnDSxQQRdk7NDf3y9cEtKv3c
w1cFEI/n1GMVhsIzUZ35xq8UlBSDiqXNcergSUOXrC3oMQShSYqFnF7psaWU3efjr9pH0GefSG45
HrO0rnw2KhQF8LzTCre3jomxUMWx1zBdaMB46Um45zTPbCt/AjkjdhpTaIMCG8061z+VGDsn3FVw
bMNLnhLyYGWEqI89leZdOADOOz4bRRBHz7pO5WXwu/CDfUZPw7bxwoveLpQaHgVCD9uTCHRx47wP
2B3ycLYLYuLfRBL8xPUkLiDdD8Z6Z/oSIIxR6gBhGb7d8h/NnDHe+zHWQFeYOYxsb3VbOv0zML2M
nlwCRFWH23sPJeC2tcfRwwOobADHgzQyUjyBnpaIcHDqE3vX6ahMk46l7s8ZMJcLlG8rCNFOyk+Y
ritcZ5GAPzCmoQ34trlbiFa5H4Mhlm9l6ckx61HjipUulblyKf+NyQRRLEUCRkxUm3h24Pd+TRJV
pFYkJ2kfrW2/LXb5hMGy/tkgRvjqKbHI6kGNHMRp+LnMs22XIhrC3PLGdI5OIw/khNk1cfxjjsy0
2hWQaIh9t+8PdNIpvbpTxZBJRiwT0MyHD21mS8Wf40irCAWw1U9xRX+7Ljggiocn7ibQk8jXZQOJ
lwv35X1jSyLeygkfPodKYshSBc0cGWCfxslPbdt2q3/3pB476R9u4/ByT1esrHnaqzxf2cZNfE/s
1hYsDKEIaJwSdnQbWRQUYqiixrolyygKGZzvvQAf7D4Xg4ngimQFBaLTtOlJXWUjWC8/OmZnWFJn
U6zq0VfSYXTf3c3Wx3Ec4jWpzLPqBhzhF3sW+T/0uZQcd91lK/lU3URYcAnG1FXu3mpbpoFP2Hk+
GIC2zxIH4yh/UdApQytSFfOnRBed1vhDt+pFcRtp8og4f9clNcI2YJMczGl9CI5VxLc+aTjNt52j
2cqyO8IMByI7vh83BM6dt1dSbDVH4ObxOe20CpKihwECFjyMNbpAG8lGhbIuIRTfKSQ+jgDOQmUJ
fM9jAqbo0M2JfW2CH/q7pg2//9jLaDpJJ/UuOLEDOzYIAxKTpWwHqHHPlqDBBVBP2Ew+HbxGC4ff
x7H6Wn/Ic697xZfXX1Fw1pNjFbgLA2MD73RgyqA5PKOxZbQNc/pmDVbZmrS+beDEHQK9eJfrPttY
Lexx/kzxbXSou/0iZfjwwpOm/gMSTqsCll69mirDPcdsam+sl9/BpvQpE4joIe3tVLnvDOYQIR06
vZ+JyT3I5GrGL+7KG5v3oFLar9QuzT4JDQFQMFxu9TjL2adXkGng7x0JkAX9W9iwG4ymYBnrbww+
vU74jKgJxdVny7CLu0KJ6EsTK2JKTE1XKu5hzpQUcbUZE50sO+wvCLmtheALlO//6iGRlldnRet0
N62Fa3IaK4fXQwUw16eVujNBVplmSUrP9tt2n0fXfmf/YlxnzgQjWY1+myLmmlUlw61Lufhe4QoY
ekNwKa9uyU3sclpwm0dfLB7doGgk4aKtR0mUkYGnMTSVc288k6a+6ZAMOe/0ZjDKWkqVdF54/ARe
RQPXNuJXhEoZyElW4AVw0Rhqsm51USb5uuvgtH7Kkpg/pw19Tweu0roDnaCyPzj0PHgBhhKDJDBw
S9gKYwzIBG5eNiNfOiUIbZ7sdp6kADW8DaCeSBEqawkF5yNbRqX/bMlYd1hn2XTCkaJSYeHVsJ8O
0NvKtx1okM9XKR4dAoJdMYNdubTcY1CfVuRdy/Mw1pwDEjhzTI9D5INl9FyJAAN3/r+IZhwLbN+M
3AeNdZUn1244Tm1B3jWpBdXa1oOePunRda70Vwr/h0seg5tfmqW0mynZP8Chu/V0DsxZnEvcqeLC
naJ8h+Z83Y39sDeqkXQwgSkv5gxZFx1vbEybye78zCPX4T3rLAf5Bw6Mg29maCgziS1tFroGYdPu
A5/p3DtMaAY/Wwr0qN6oIqWpbrOcsi6OeWNeH2zgZkUpy5jGsikRyJlOMdvBx8jvMbdH/Agjc1Ki
HcYguJgorFyftYwegIEq8sN7IvuASLtStyuTUWCE9MkN2uhBlpNZrF2itB+7L8Ca6FarTyEsGR2/
5MF721Ul/1pLCGKC/PMY/4/g6reauamDkAbJME6kb6bEtzfz+JgVrlhDbtweIx0dDFO7G86lZKck
8g1RdNzNphHTUPTiJNwNWO7N8gy75jd5dcRHsvO8o7XEznYzQmghNUg2DCbSYBCUuD0g36R9vI5E
5R2wN8VnAn0yx/pcOTpc6Pr+TTncH5rYOwssHqbqeC7e0FjauEMCw+ovJzU0Sa5U5BlY4nzMQCZF
6MlHuk+/QfoeIMagExxr+hqz9MIXOqepzIq6vkNd439pbjFUcPKKIpuTyCpfvTFOH8hD5MF/DF6v
eVaHQ3aMbTSaYmfTnSqvMesSODkxXD1yd4ceBmHhCPfYUt8oZNL0MQxajL67yGaVZOYIpwW7/Eey
48pqFJnpYzIyeAoIUaHg6ZmMbb+/dAr5LOJzUao6DJGgKupBfZWeEFnUk89FX61DO9wsMhYrQGBY
zx4vp+nSltUzQQh8rhkkOKlbb9ndX67ilM/kgwXGMlh3E4AD3B8od4tTWv2WhI07vY21ygmvIV/H
RK2Mx46UnxoLSWZ6z9h14ngyD3iSeRTLGbaT9SPuCDtQ1ufzjjqxBflIYXGkTUICPbGWbCxsmM12
XHpHHzWoYvYcdkqf/42KI3upShoV/58IZPRfaWU4C+FYfcoShZmKuRotc83UHs9lWCLhJyeVSzR7
WaqmRfXX01I9sx0PeKr1UBvZsOxGF1NmPkQ5ks6jvUtaTrPYVMUVeFtUTdQV29ex7xjTLY5SauTX
RMMN1B3pj0Xthd/KI/QivP3TmysXuhOK3ofudg7oRyALwdcEL5xMZetaagbqixmozY79UpM7SzYF
X7imteYxu2IbiqMKtUlha6fyy1rjU91P63KvIc4s/eqsjLJzu1dyfaDBRZNUB7fpzfqe4i3Lz/Q0
e7hXTiylwhuXvA+oHRZybie5wca3/YNJkbrBRkUfKBwSJb5/MFwbKm3YZgqv8VmeXu7qCCvtMFSA
8TVNs/UMSNrQuAU0cJVJhvx2bdxJTD2eRbsjE2VKL+yyNiQARNbRc77+cxotqEZDEG9wAojlzfPj
/G5ZSkLq/ZQUggpB7kWskjUInVx6SRLThhdIHAYgQiseD9+7EOEz9blLeBGn89c1Ae55GAqRrDKN
N+vDcleAeD4M/JoCoezIYV4T0v3igVgvqnstgBIgZeMxFJCrYbESlJRrovpb7EPhE51Z155vmYkc
a7S56+qiHoAbv74X5doMR+9Ad7ADa/s23GoUKTZMZcnsCNuefG/Jz8YX5L6XBvZ+hiQn/I9SiySs
S1IHMOf7SnKAkxSrtRjxBSEQM9/2xqVf24Wldy0EpdI/ZsLCE5V4/RNgqZvvx//5C9UkDc97w8D8
jUQTlK1/ssNsitzCLyh0XZrY6oN1hfAVYwx+pBYDAHCqFWWIvshaB1Lc6XahcY5p7gYjMgWQfoi6
QPrd61+D0JOVlZYInR99i7OpjCN+Bu/tcy3gV2xeFTLuTTcoFiNsACNNDto4YjGoNFtaAZeA7O+C
4SsLkwzSf+KcwMQIMsO7fDB3qgjfho/D+6db0jdi/ZzvfrEP8w0D0i1IwPMAxPoNeZDHj+YWK3tb
wpbKN7uo3kqVhpkJFFqnsWfjDdms4LLdhw7TfSH549oFff4a222iTrOLrO87OtFcod+6jkhQMcJK
X1/NlMLKH/o3PCfD+GmVVJe2xFnBQwns9UuyIYxCTud+ZgxOLG4b4G+Pjywn57KY6yoNELbNnnqD
52px0wmIMMO0pPlCigr9iUlJrIZHM2ggug+Ea779Y6iXJltmSXvpEsoN3fFcvjnS6HhH/iYHsXbd
1wNku1uUNMxQeu4nUje7VcrOpEMYvLol303Aqr1EJzOTCKHiB8fquOlZQ1OjtoEkpPFuGgDs1ecG
OFbgGHJEz1v/DLstTSxDBL2yIBHMGjtBSR5WG5exME/3oibtdgOVBH/ohqvGqR90eL22XfYKmsXD
XW0F8ORLSRZl79JelgXSepZjrp6WT3+SlovgRjjhtT/d4tFgA0wQ/TT/Na/zSJjqgKnHRxw8VYbw
qcNJYvUj0+YyynsKdyZoClcE74Q4OP545xPIaQya6heSHABRycdxE0ACfkDFfmsiGW0Xw2SozZXX
1vusOlpAffL9OBNCvMIbTMlQB3knQzxCk6zdlUPJB4V4BV6BKpm+Ee6KJ2+Mbh78BmSjIZbPduwk
pV2R9qLibnGSYjXmreE+H7N8aIW/cKaULwZxgdy+v3vLVthKJgkvKVfqa/q33H3PyQnSVkkLG2Yq
rohNJ1qmJey259JbPWR57J/VAaLYI29oLGFGsiTC1dkftcPI8gCIaRzuTBfm22GKNgEZvGfbSr/d
9lmFM39pYQTJ4b5XuAdoY0Z5QliPgu+XZvbTvzYh+/jidL7RX499cnQWCMDzIe+eUUHMH5HdYj0X
ylor+r5d/1TbztI9iYhC0hB+6g8pDxKzYamKLznxt78sryp3GuDa4JC/F8/BVQeH9YS0aK1ikzPA
dsyiRgZ3MrGLinx5MFjD2hyiFPJsbc3ejczpkVm6mvX/WKrjajiCVmfYlSn3dydyM9xpuIOy43hf
yvDD29gfWmwV5rPKNl29fGdDAJrsiOKNL4kh3WH8o+ohu4DUsOk8KfmDj46xYPSApHBjIDDw90Eh
1R8J65qFFPZyJLUt1dsBfbuwjKALGK0JJ9AnZSJHCIsCwERO6hkBZh5ObsQq2trk6d07WSktBgT8
AMWbEEm++DBeofsd/24LFeBabwdEAmefKIrdVgypY0CIwf0qRzQymS3GWWMjkYqIOslq2D3IcK74
by+QfW1TqIPJXiL65btSriLGD3B4K9S5MDJgHmnIiNG9+vwV4q8cLt35OQjgk9DVO6dF1wx9T57h
PzLcKlREA/I9HmeSbJFXqqqzwNdbI73MYAjX/SSt5zL84KLufLK5WxA5k/R1IlcrsfDxyZLE9UyM
RJW20u+N3Mi/1rP0/fJ4GbZrgthKjTaB1286v9fudXJcl7DsuzhHdLR+Yqz5zfO3vrbu3AdegFwT
Ij5bcwQuZVpmjRQiIMB4OoBufdnQG5b2zGOv7HW4SG+f3MCyLUU9Mwrq8y3nKVZlwy38QqpKz4jH
m9aqMFIj+zDesOf2bJI/NIuC6JhjfwDuEEQI3yJKgpBkHjhHCDmn0y1hSW0Lj0wYob8CykwUr5g5
MRK4d1oQgv7XVYV/FWtts0BYujBCBzgoVjJc+Mj+VfF4O1VRm4lVYPqOvOmHHa4fQvmPm+6aGkxg
l4j+T3bYmpzB7IIOcHkLLV5YUm4Z7j/XwfPyVY8XkGH+Bxn6dRI+ha5u4IhRwUinaIVf1gn9JfZf
xYaXSYwOx4YTr1c25WiwpvpyuW5J9D/g9iP2fLE3E9h2KiHJdAzxYnQDt5KAgrGQnjtlmJDArUN7
J+MJ0nJxvMDsojPjx+58Y8/i2N+Rz4VeKAuqzzuQB8qtWQbRsfFhF4rJOFW5AiumrKOirCdXqXgJ
N2P0nnmMs3/fPG34bhcwWRvtjqXyrqJ5ge/4TgiThjWccwQfzxVwSTi/vFtvfE+jUUwglY6CLPS7
4ZKCS//RjecN/ZWk0S2lZMUlrcoXojYAD0h6W0L8O3HHi2CQQV0aDZancdzYKJrN9YtyvHV4p8OU
uPOly368KAQ/QeWroj6Zd9f0WEsPzYvKMyXcUZOq6++fMo9b6TP78+5xsxPwaaB/aPpGeSWhQzCL
N3Lx7ca9pPOAkNzY2zJX/QcSbFO1OjJxGqtHNiYEQJe4OrcX61IA/9VHrt4U3SqX2D4trAHteoTM
+fGLDBvYDatqRp0buKYciYpTQtMRvW8zpv50hz72uFINzbMFiBHLgG2GlCC+y//d0CdJ3Po3B2lj
ss3CbzJyyOcuFKXMsEtuhDD1BFLP7ddIJnbxdb00OSA7MCOR7mis1y0eNTd4Azl1JusnlIkdGVHf
X0LTQN1mVC7oG/vVWSBY7wzqqSyoOh1a/7lD1QTIfRvQSQz+cZAL1iFdZjZ4i5N3T5P0OtkAegtK
UkI9aiWU2VmCn6ZMzc8F4Nu79QIuZ4/tW7DM18H4ib/nPpX2vdlOiryPDtk2mS121JJyVVVpDIR+
5BEolmQ1wp5kGHn4+2xsykXTCpw8kWb9QZCXZLfPmPEtsu2Rf2S40SQz67NRlP3q45LXUgUv846c
nDLV8yZlDC0TCnfmF/m9bNqifjTRUHnQd6eh3QSXvLbfgR0h90DgF8Jo/sbTIYhJJawJnM/Sm6oW
RktZ1sAqfimlWx+tY9fruXNK0ZpH37hehevAFu9hQ6ed9ZpNVhhjrJqWo5TCV1/L6y82fe+lE/3f
+yrn8vBNOqJBHN9xdam6+qyiQHA1fLZ46r9UPNfOXKl9drA2cl4vao6L4J7S+IDiVIu8hq+a0dJ+
njhewPKgSWc63Hs3mFPgrnqa6eg+WrzWw7vqHMua1mNa+dkVzRwVMq2++egocBIvEzsU8HgHaa5r
c/JvfdIn27AHCPvNqw/hAx6IsMMq1Eb3nEYZ7c0oDJrOdzE+nNL1YML2bdg+42DIHbu7hLhVVJx4
jVnodAL+0GVQazm1S18UOsH262Xs1RkqSLcHkxAsim8P1m3ySxZaXHpPNoufSD2ql6Uhs/viIqjJ
tWTNbTT8ZwodF3n+Be1kuegWdw3oJyRnxnuZSeiI8QZdcgStl0kMkTgBbA/8jqyYwmtfyrpvSwMv
dNHej9x5qCeaRdN+1HMzoThScFHAQeDOGUw0MBQh/AjvYHwM6VGXhAzl1iLW9RH8sqEB58TDNf5i
1P+gMpL4QidObRP/nV9pfs94zsyt9l70qAKPdOBy8EFRyVWx9VTsuZNL1jwxRseoxFQN5L0FeCPT
usBvmTHWiQT7SaIe01ESCXpYDUlsTnHa1dp7N9rqVDh1iWqC33XstsIKjMZEmaMrETsI7EyoPaDz
TX+PtwJKTYAtSS08UYAIxygmRvlIFOzUNfDCHGA2olho8svqjWfrMALWl2C6yxNLJ/SvMGxu6AME
iJ3UVa0fv/YbefdA8GDeUveUPaGEwcmg7vpHoaQAsRg611Sc4GQA+mrSnIdflp1Jci7cE58P62yL
1+xb1UOE/JMy9sWd4ax/nxpNjNpgXPsE/yzntBSdNcwjfYI6MkJv01iaoOlMECKmcsAJ7TyY0tGM
8gJ6GLJV6J/36cbUArNCMsnjue7FOtpakMdPWfQfQj2Ag/RH2OWzSNG5SYImcwZDfuErvWw/B+YP
iiOiPzBdgZLEtOXtUlPGlQk0F9fFgE7SzCVSsmUYtfWLDygsJHtLhZ9hDWG8M+lCWwp4LYd1HyuF
OeRYQuKowa7dYHM1p45OKsuozNZVGgLGg9fy2Dy2meKEWPlhM2L7KcHzfQRieZu0KGscRhCLudiC
WnRlJughDtT6B7qomdgicSicoZJw3wPLNW7Sal0mcl+Z+QQeCpr6JQtFej9TaUAIKTWGOiYe2y8k
M2XWMRCZdjEuaONDNn8S0yF8v3aB++K4j6kiT5btmAMiZ1BJ21oG1s8HguD3lDZkzMEEhwCTN28I
btwS37IMn1zf5aNFVdC4E8RKtFGryDFtMMAaRWWaLXdctMqTZchYEyILp+IKUsyEftQngRYicl8q
Kp+nfEaEfIsKvoK/rjvNV+iUpa/1QwLl8QBwdfrWFV3WHeDAOQalk6fHAhwXAbTXia9l2+VQU383
aiX6iKqmZyEbrCePE1AjUrfXSTbxBxrGDIJjb7VljoePoXtU3DitlL1BKn2+6uNxz0BzGyR5hdlp
F4i1sIRgTiiIeGfSjSSDyCSugZ4vUsOQhqH8jWh2hRqndDS2HuV9kEm1V4i11pkqnEDvBAONbTV1
/KgF+llvA22Lh9Kar0q4vSofwfexWbiozaSDP2TiABHxzTsiyeG11R6RzaKZTtOPZOfNiPhaasLg
vI5elLhXC/y3kHxEqBXy+dlsg1DXo9Td4lUWGUif60boYX0u7CQjunVXgyrsw1iDDXXurJEoZ9As
gXAopYFlFTidxDQOAwDSyag2k2qkR7mvt78XlC1DcIQH2kalNFAA+ys1bB9BqtAylPZXi9i91I+2
2eh7y7tZG0mUF3geoM2+G/D9LTWdHejPg8hu4KtvLyF+MnBCRF8NsHKeUlAb+/l9ALVeq691WEM9
udKPk2eHzB0Mo0w/ES/HaU2CBe99XLue/BO5y8n8GEnuVgp6A1k2yEEjkYUETtIsfc3l9mg6kQs6
qMcXqjUmK7svaYqx69M06smM4eX98USLgcqq0D1SY1iOTrnrX+OoGFj65EtGhTXGxrq0PgbXkxaS
gwB+l4kh1jR9Gnci4vR3mfXL4CbVmcJRg2yVAamwIntIbs7fFgBR9FDCWiwaDKK1Ymd95tUcWd1u
kJNNt7Mr5M3JadbzhnlkwwvG8eigt4qSW8Y/4yXoksMuOvVsaZucGzqfsqiMhY5pTEEfDuGG9KGE
MNkz2DtWDPvvMS47qK1tqrQQ1giwA79WH4xIm0X20k15vh+g1ZJ8k/XPmkM8kCadIxhpYGRB/Mtu
HMO69zPDzFrJzSxTQvkGrqb3YE61P0bZAVi7vNRyNoBFVlA4tZl5sy1neFMXwxDpipUDywsk5PZf
4R4m/ha1YWFkOid8vFgVAaK+TJb8nZdzFCdM6cd+fjEVhs+HvFBm5dQfoINdPYSjkYkIqwQWLeNc
Jwj7gxeutOt9vKLMvS0JbIka7gBQg6x/TYjtbIFm8m+kSQb5NTiyTN8floAWcWP+4bJJdA8X5TuZ
ZbqafIMmUJ/4bbJ6spY5ofRR5KhPtrZNn4BVFBBz4zL2dgizLgG0cTuEFStnMKx5Va3C+huULqhf
Vc7zVFxu32KCrdFG2ezdRdWWgp2e3xlwK3+bx1OPmgE1iBsr+dSiACagk8aaTKPxhwqZDoSjGdRe
GkBeMpgbsAXS2lMmQ2fFji2slmWhdXZhXMwiSuafx+Y/2zgpvN9tBH4ulKNBUwvqaiYGsvk80MCI
evdXG3hiZ0A79KjaYub4LMmoL9CFNLWKjwPYv7xPdg+TUc8Kc5jkEEwSm/fPv+DUT+PsrW+92E9Z
lM7ulEm1RA4XjhmzWax6pVvQAUqcJkBJ3sRCHg0eYag33rAU/oFEgBu29u04duxVkVotEU9IYNLy
X8xJsqqR/s5B5CpY9cARAZErOoPAGqeFMH0QC7MceUW+bgk917vM0VdA9SOsnmnWA/2Opbm6Btia
N46uYXIMaI4gMtVxTA4vVVCAjdD576ADTVFAR+1WkqZGtfkwdwCZQtOY9elT81UXQCTBgIY3wert
PpdKuXCkik1aoN3f8cil7anPWF0n19QVtTnWj8MNZ90fHLFCdEjhvplU+YrVO4xrDCeACM8BrKQ5
K0Qr8MRG6Caw9+BldrwAYdYc620wJ7c+HBP5rz6fMIdDMAjC9agT7gN/gHIPZgCMPMMAOaOuLp/D
p9tG6d85HJQofwA2yXAPTjFX5x57SVoM9SJn73D42V70PIktXo4jv3594vZz30VOzmDHt8qK43YX
y6X02fNwChrosFcx28/cCNsELzRSsUFaVlApxpDzgTlZsQqXRopKrBPLFyZq4orx5Nf/lla2PeMJ
DFpmcIZNfhe+mFVEAwmKAYxREoQTRoszjUQOwlo+f+0fKAvPKZ1crKPCXJj0+XVZ2CsuaLvdUFko
DZp/DouPNcTo0aooP+uU6B7IB+GBCAc1bAlHEaQD5BbSwphqzk/SBceVWlNod8h4RVB54qgjGCBU
Yy5aQLMHIQ12Q4EoNgujRDET4OiJk84SpwjCNDT84xWhdd0am6OhIhzyacm/Zlk0OvtCg6aqK45d
ey8+nSu9MWFM1EMGDvHVN5pBR7Oc4Cqg7qrTQWkU/QswwUX4+u/u9xKW44nC07xQivbTMO1GBByk
F4ZadeG5F2JlyVdRi18S4Mj76qYegBE+cuvppkWCfNOSTH/LbD3DLx8IGlOldVr4yTqgmNdH/jRj
WlWOpH+FtL7Zi8zhhvTNozCj/dVMVxuK7EBzuDQ5NPGryP6sadQVwwMMeKntx89c5KRzqazcvPRD
FzuD86Wo2ijTuc5zIJWOS6GzcZ/Z58pdswT/jboGzZ9IIKni26HDeonTaUeEmGQAAxrJB72dt5MN
TiQcSe5RcoqwnlsH1+RhgWpBZoiVc7qBQZXCG9ymIa1cD3+s+I8p1yWmJiTrEWYUyYQCGsL3EgIm
SyMH+VFSVWxsWD9pDy+Hum3FN6yZra+Lc1nb/bZOe1aksA4+W3mHmswPktO5dCN3ElNe/Q7/naVs
/mfUqlMIqqj0EiC5/WMcXLjlC5/J+b8NJn+UOODh4IBEDQu6AZt1vXECJIwMeRwJVbCFobGgOeQN
kOoqd4Xigp/ICijzwF83S2+v3xKahToyyrZdpIU154gUmq2zMUSqTZaHleHKDbVVD038VeZ0LLU6
G/0kEL2ULE+jiYzX02flZ8PCWHQarLRxXsjjy0F3assbmx2MMjqUoOVRu26dQxsGC0iyZUAkXdJb
Y+YAUGgrtKbMpfpknfjtI/GJklcU3I6s6MuFO8ZA3yE0MfPkP475dff1GAA3SKTkVxVjSPYdl2qy
fQmp6FUNyfJklrs0IbSpo/IGMH8s/0G121xdfjMCDmSMVUcE+yUSnovcT0NPGVi9h2Tme0mlA7K4
ILfWOekpSIMCWBK0slTPBmJpKbiC26Yr2B3iURsGIe8K8ceVDJsGMk74syUvxukUL6ervOIBZupl
YnjnT1kMISRYZFwXVhKRaVEEes48cW2oNY4+v6kXCJJ5RjMrigPLxY0fNkKdKJribnoqXDDG/cst
HX9Gh3dRYwqm+ruzq/wwLPIHPvFKsRBG1r782sP1rpBj+yy0qwXe2WsuchsBc4IUCLEaFSfblXEJ
CTrEHRcEKf3qZmbQH4rTFvuNj/yc5NS+5gLCcSrrrwRnpU+a1zMbe0WvcHESz5zPA4PHovb+Ey4v
gxFMvXDYPUcRYoHBR5OlC9V1bLTa66ybrMkoC5ckeTKRj1BykdWIkaajgbP/EMiqsS9WIfvcg68/
J0j+NZMJRS8/76wQl/SGFXRvxyopeInJLTcIR+6BdJSCCZTP5bR/jYi0N3zWrHioZJua9LfGa0Zy
tPNJtFobkmOi7WLGGhUSwNpaakHK/ARMaJxUvdlAPuki/t25bKzJEVnGmmylBuH3p92kiIqsGeeg
dbJDVlb6rMkZtMybIVvD/Tm9jIbFmyIKAITQiB/mUFhHPByqg3/xeiqTaY4fD0PCC+FwgT9WQ/xW
0KzUrdqacfgyRScn65WDSbZYSJ6nq13yf7461g3X3KcP8jy2TtlXACVsw51IWd7OJaNKWgPYZBQL
xIl6KhActZXbg1Jkgy73DFfBESbR27Sh6YUastzCGuHav+UDYsJKXXMc2TMuubRPFmbB0smUWZjt
IVDqe0hZgHCz3qpOiQ3N+y1dd2IvvyStshSnrV6w7zPenSqcVyIANLeTjanIaQFTv0rAtYXNCyqm
QRaziC9q+5+E0jjUThYP6fJEoWqU5Y43kHwgucoO5/7NxpDwTAjXtBXF8VVERFZ6s6UIfgqWfznK
AjDLSdOJ8c3Nr9ngzZyQyvHq41N6/2x+N6msaFyVxG4sKIkor/IoI7HKSfg/gGFSIre+gcwtu4wJ
nQqZjmwP+8A0lT8KygX3lJneQoQP8/v1HAuaPCEvijpd50na7i2DpFFtql0TU/zuax5/lAnfukXr
WkXt9l94qz8azhnLRQ+t98MQbGj2P9T/hQ4byN259Cz+JLUmzo0U2TYgyAaDfl7wV9ardFEh8dDu
AAIYrCIC8mbcN4PyvYQKV0cb90IEoy2LCIKCrDi2X+sI4FnirQp5nwRU1OSJIEdbT+5cOv2lc+6/
W9/xrZEy0YStjedWPLDXxofG7UEkRDloesyLPAj2m6h6Wb9iXUDM9jcinBl1SGKcAeChzmhpkncQ
kCkh9Ae31RylHpl8czHKuwyX1l8UC0+52La41e74vETqtQMcpiBPo33Ks20DsO/N9gpGR8yp3xkz
Zpsd39WSIhr3a76B4FEC2lO0nmhSVSxjtXtuKHqvCam0ykykqL6jl784rDC9xD4A6sd6Yy4+KZzY
ZwzJ31Rc9dG9MhoEGTIPfUncRhZUZJ5k37tmrEyijWHOFDA1GvJT0qViW++K9wP49XDZNdQKFzNB
hGBwVdgFPYN0pyZMTajaIk3npd43jI2Te7h7+Y82ff2tclw56S5LyV+WB6GRLWPkLQEko/rPHEid
Wg16ci4d2/8L5E0aRvXu76VSNl0YmjlKZDZcn+SVJQ5ofZ0fWKy9i6V3A1nXDOUmo6QcflMYQUTz
z8GPbfFCJydQor+efjRw5r3rhZlJMHMUMmpFELqH4/VhvaySxBOD7OAboKNvGtz7KMnR0qJ48pj4
gYPVU43RCCFQqxAOaqlgCQ2zu8x9yKzAmUjIHefJNGgzVaUv6xkW1KCBkppd2ng8/ol6PyVqbvX2
G5WKERvw34TRdIeWK10Rm9yAqnSbgtpLNH5JsnJIIg56AMFMiFabjKmr0d4mMVY07/6YwTAirQL6
nOPaVxYu2izyixrYeo/7KY9DTe/XUBsV2o4NcpHb5/fi6T0KG833Xcj5V3WsHvikG/SbMq8mM/xQ
kza50NjiLj+RePQOrETRPXxTynQQ34qBIpMovbFHgaoJGIP1Hj79wM6gpDIrOUv/2dC7dTaN5CSb
DMlAHzGPCP0WpP/5eIi11YmH46TqXNZdp/VKjNpd4WPQxjIWxKT95JkS/g0HQpDE1mF01/Wd9EoF
HNKb3rb3USLJzC4F+kiLTI5232ZaEG+3NHeFh/3T2WZYtHoZSb5tXiS6+SqGz69uNawdnRh9SbAw
s9RkhTkpT3t6Y+68FfULGHCp+Pr3D1lFcDMXmRAYwh8qF+7aqhlNgfZfl00MpJNsiN1e5k0L+reX
EzYOfpJc+iA/6YCzUf2rulz90gAxXizP54ROOU4Tt0SoEV2qjKtPGzGBWmm/6J3ORanCEMT7jMb2
V09dW9kVLKT4pLpvMsfPCHz3egeLK89W921tyrhEHxvJgUNrsz7YFubZdrwOo9tdZjO+0SWJcPkH
3LbYSZiOocx8R0B6zKajGwiNPooAhGy3BbBJh9Y/TntkeoATzS+gf75EUoaXDroO6PQeq/Rm11hX
7KWOjKEQo4QyeiQUN0dsYVpiygWFamWzg7sHTdxFmQFxmMWtDXGluJYUP7Akc/DhAnklL6pvIHbv
W+MmI1ryUDAeOMp0jV3jgMYS40pT+VIE7q5uGr8vXBIi1TAM3NjzIBmpTUrYOd/EhXrNa2QHO3Q3
htGB6R1KcG3GbwEf1c+vP1Vrr3yYaFXQyaMPAGMYleAeTZbV0U1NHamNp4XU6/gu3MKCU+6JCXyj
uDo1yjUstHmLKVcHQG/1oIDAlAzMOZvVttSW3aTaGiTY8PgggGWdZEvkaUWs2DF7spyFYmRkXcRJ
kzXVTbjXEOuMSdR86OvRgwZsS+NiMbJhd/Wno0cCrXZfSaN66Hv3iSkNbI/6enmRrNOQm7f5QiQv
5MmOjrbuPgxWD7guIjBZNn9/6Fbp6P6XYLwUPpB/fHvB61SG8HqaQ0wra73UtoREr17tKsoC4O1h
W88sfXctob+vejH/rqRE7LzPz8uZYG2CdxCyVouwbJrtXbI1Faq66BswbHs5IjITtzeng3vZwIo3
g5TTN9Pk3QtX3mGbMXKmBRg6AKmRys9vZI/pZvY2FlehxjB4azf6Sm7133B/86AUycUulL3fZ9KB
3ARL6EqmwdVVuSrzwcByE00peAD9kiBH5XLc6kYzjCMZNloagKQNcNYSfHvDNvy2bHIu2hCKB74I
WDXC9sEtO0izjijqxdhtIvXPH/MjyHbyjrjenXlEgFHQ+fULiDeih/dZ4dbKtGau4B1XHiVNlOGX
N1/6ILW9N0KPjfod5M5WRXw7iEsduE/vWuWrjCFnFG8eiEGSXl/Kq5Ku1L3R3Q5uOpsT395rZfZL
L7tVGL2/r6GckWkXKUvy/v98smatOtyTcRCelfJyaYuh9mjbSZlEzY+h6jAonDuIyzOOsQkhc14M
xaDcIQFjNsR6kzJ7PBuEhJpbbzBaE0U06WLfnoGLOEZIf31XbB3sx9KAN1KgnPkc3t+WXOvuYIyo
MAyHvAKedVW+iEKisuASQAYztXDMlFQffGnCYAr9G77OxK3R7wZzgcwT221u5bZ6sAefXM7jV7An
sc4kWIACg7Lsp3qjNN7PzsIBiKq0pKdjRcJafnZqePJUUcNRH5sPkgqN0OuOZfAMrqNtGBSYTSQ9
qDarRYz2+/keBq2WTb9CZ240+OlC+jrlmtGIw/MBcNVmh38Cgbyegw6thhSkthpbG7AHw/TEre0o
ws4cPr1HNmVNEx8kPmJjbS1LPGZMIEfoAZAs+H140sb0WgVDA7Uo0Ybky5+S3kDYGDuvRUJflBZq
GM0O9d1mZa21uTOVqJYe1e+9wAaApKxOkapH0ZqCaRGlpFL+2a50fJsBN4RNd4w2noYAYd1qnhTa
qXVHi5WHcKowGcewRvB/23XK1CuOCbVOIe2Gmcnx8IBE6DDLtWCGYiRTWXyFG1m8uDQZ0jaGdQ2j
dGRJFt1v9n3iwTwjDzv/Tmv6blrNIj/Fnc2aU/P78799eGA7wIuhkTq2XaalzLFkmQAGUTkKwhyB
BzirvBalWISt4RtuH3GhTjwuNf6Ni2xa2GagoxCmYpt6hOabuXH85+UsP20xCcNDxY3OkiyeSSxn
KdpSXiScGaAauY15oFsSsDy1S0vlEA370R+bKClYp+jsrCP6qb8idDW5N2oaeUxo+5GDEMJoZhoZ
zLa4md6mxhmuX4IDZnM3gkX0jSK93wO6Dra6ifs7NH9N3VO8NEwxZYffyo6zlHupa6PN5DC0wUsI
52kHZDHJvVIRuTdIgo1mVqmZ7LqDA8yzgMocV6TLj9o42kraJy92ob8n3HXvjkgULa+U03wiNGyH
WVduhZDrtjmwDfwX7xm1j0cyj2xr+y8fFLDvqnlg0O+0ox+JnduUsl2sPbWaSnXma8PAMXdx/2+i
u5etlppzXXnhvgmaOaslR3+V2+dv6VSotNeQdkA/z90KpZhcWks0uWC48TZRYFKBuNWDrZ1/n0Gx
dVW3q4tudUlYr7EI434Jib34F3x/X/kfC+w4A1++jk2H2+l99nPgI46sUyqk1xZzXhruhP5qFF88
nRPngucK6bc9WEgAK/QI1oyIb/MR8dwZc41/EYONnfRxF+xnI/OZ1JWdtQ0hR5Xh4kSdH58WhuAZ
D+Bdf6KtrlEVMMf7LxEpAEplHgBZ3nU+QHEJ9iS0R7LBWepnZCn4Lu36BkPibuerX+6FW2KyN+7T
cdQa+XtPHrH4kE/8o6F6oCaiLGi4nhVAOw1qJT3dMVQouALcKW6g8iG4rKd+UJollzmYmmRCmaec
QSb71y9W1zdOX0Enpk2PppB+rgQ9vk9gZ7kZJplTFfPyOozmrFfUJCAUGYYT5cPf5ACseAzrCZBZ
pobmBwYCYq+cudvAzSPsmVyTmEhPFKKPt3nEvGfS43bWleX2P8meI58POS8N/IG+e15DJ1pLs0Tl
Wu2PHapsg7DkC+HjDCvaeAS71DkmvC4Y/no4QzZ0m2xAVerXiCsoK1vTe4JF/j9AB0NW0IzjyhMY
tNT6lMr8f+BKSBILwiDe3miveRB6zUl1EPhRPWqjfWcr3crN8OBAR9u1T9ls9EGz101cayYTcQw8
QAx0wrA9uvcUo8XbSRHUWmZoVRzKIOIT+RCJnAM1kLaioH5joHjfPJYy/9M7/zNXdxSVVDnMg3UO
HWNYYCEjBQUmY/jgTH2RjHO44S7ZZO4b+kOwE2yLeNtYNrnRK06c6A1RPBED4NA7qjf2PyDnj9o1
4wNgh2EUEmR603N48V2FMxZyK4PJn8E6/LikgVB0f8ByiEO+bdiJlXrLXNqk2twuOCgsKs9CdpQf
3TPV6Ktgu2XhpxTHelHjN98uZjmRO+0/CSY7Y6JBJ69zJW9lXSyDpwBxA+8E8c9L7H1F7jHlfhAB
5urOtCLTXdYngFjj+yVwp2OgEWBp99K6q5GHd5hMGIeuxFpVfL9DRvnIe6tTmnJzv8iTNo/roq3P
Hf84N37fj60JgWjk9AFCvP5BrrgojRt+SmKTbCq0y9zbsVGKBrjs2bziFG7CGSSiW5GUyEme/shL
eaYoRbxXAOWcJtQs7KWHbVLwBAesWMRMzKmdKfo+/lwiM3trtzIahyM+sRO8TNGJbU2if8XHKXnn
wrzSvpI8NUeImKjDYJ4dw59LMX3m2WAuVVfRR2NexnZGn7X5uLMBtnyaECO5YxAyl06RtFyJkyRi
3acPagWT/RVanLmdzYomW+R5D24QIduePGcnOhTlYu8bVjwo65RQnyzrpiNY2AQ+2q6gCNlB31dA
Bsf0U2mOEmc/RhaLvQYtT2xhDWjLVcgSd5M/FjpnxieLfn56Y7AlFSkqVufeDCdZr8lLHtuIFj1N
IegRT49zh79o8H1XSdMOLvm2xthbLPdWZc1gQmvA5XI/ox+rS75fcV7wCSQ8WhtDhB0T/mTen45i
PgHGemueXmWm85f6SUTiaY12nF49phxtlBcH/Km/FPdSmNzPCqNq0Ojlfg7WYp44BkNmVZFhTA8M
mG0AjME4W5/HOE4kdIT58rSGREAsrKtPArHR2LBdEmtBMF+utziESsmShAdC+ROZcp7oDqUSmPQP
Jfi8EMR6Gxecrfsi/vGFm/0qxzuwtEl7JzTb3BAOy6EqM0YoiiHUY1XDW4nDnFacqdu2O/C5SOiE
EgqFfx8e8bEqzuiFergY9CJlPiMN9KfdsD+mb3K5lXixHFE1ZXazuD/Vogl/4B7fSdlvq4Zfj2/z
SLjIa6vyOteDrCPaPwRxKLk3j29vxiAmlUJAI+wfQegG2F8/Q8O2j/ha0VJhpCIw3lFzYuZhIRiv
31wjtuqozamwSpyh3HbHeXpFsValxX0pRK50feMUBtMcoZyZWBXvCS5GlYC8Xa+1C9t4ZULvv7jQ
zilIm3Hu7pJzSDu22O9vDWcli8gHF3XBqauNZ0Y7HePEMKbE1S77/As2YD4+HA1QYLsheFC2SJHv
dHXXys3hjaOtR/Kv4O8U7Nn/PzirALbg/z+58QbPjZRr90G4k1KqqZ8LnkDui7kBWKZNKiEM3CnL
dkFEacNYReTqzWjjk7IzqBrKKdxFLjSqi3Z9juIVMca45hZHBS5/cGNjEkjrFkY/XAByQD9my1oG
xVK7U7SyFQYYspJofG0EK5a4rwyUALfjo4NSmEuCNSwDR3OoptXuyl94Pn0wX6/kBjWkbxZ/0HQv
TJmOQyFjoxek6+8agDqjKpd2JtMYb9tkrdOz3yRgzDKRFGar1KpkLkGBM/dSRKpXi8FON2U2nJ3S
uFCyOnq5qbdkFN3ULouaVxhS/BX9d9VUDpwXqEqzW8gfo26STP63w5nBW32z52ltXZcj6AWQz4NT
I8SEYO8w83AU1fMHCRzc9NsDxH27lrcoyYNXbxE3p4IgyWq3Y6uh1Iugt9Dtn9MI5UjlEUbe9hl1
813wCwuWaE/PZ/REK+cLSIoeLA9aFXzdlKqrHnytPIKp5ynRzGkVDsC6qEdzX7SPTMHwMcadRbkk
c0hA2ImtGqBd0OE/kApdAOUZij38NOzFWB0Udsvd7XeYwr9Dt90wxFCnJRFSR6NLmML6mxFSuDQq
nzAKVXuC9lCq2UiolKfACsbJUOeRf/RVAWMOXTyWshAj6H7+WtAlFGvp170jodh0t9cCvEUsL9JW
CykHtJZIDrjhY3as39heI1uByaWqhtMeVLskOv7Lv10o4/cH8cJ0qKYv7oAslKGMfbbuDKFrj+HI
fzG3Fgpj9U0ZgqtmP2dOZf+pqQ77PHYQ5sid0paty0tTmYxj8KQ/QJN7fTFGKV/U0waBQf9JBKuw
ukYQjHATucDn7l5eZN/PIv9eQt0rTo/sMbUWPh74orPavRe/7S062I/1DDco2BJqAJKb/KOIoicu
0y1cnPO8R0eRO7miYBUPnz8ykp+bz4xgWCH3bnBAFj5DQOsIZVL6e8kErWhpXh3ePkqGmxNQLH6q
9UukfEFY3m8vBpIfg4TpHWhiUTEO6WBP+oYy2W0HokjlYc/34xRe8mG6vJTgdMmW3+MLhnwDodU/
8YzIyDfXa/jBGcF3hucEtqT9jeb8ah0LzfbevTxCHqULeD+7/YjAm9kfBwyLLTFv82I0Aqy+70M3
fRe3SKhICf98/Qyp55xJkDvFtDPz/8sJ+UAcZPHrADBAbEjpd/HniXRvaUNZSskL3li4TDTSqw/m
qVYzuyyCi1/COWsyzOIOC2bQ1mA9k25SshtjYfjAZC3V0EU4M/xTNJmgAHQ+ajELe+cokuqA25gu
KHS4VUniuFliohviwLkqanBngXEhWgtW7qBjxM0U2XgEzmECxYK/foCursNYjeKSleODnIAefkvc
3SDBugnelQERV5U5DZXeN1avJUca5BoNg5x94NlxuXEJfOeMxvJuCwp3YTDYy/+O8JwjoJeW/m5u
7TbjnS2TX9ZQVxNCVQ4sbCbzecz3ngEkvX+2GvZOCwQi6o/8duXwkCOkGfJnSx5qePnx67eQJ5HP
c3RmtHBoQeXcdsdcc0b4CIQSl1U9uu5C3dFMFC7Uu+D9exYA/5Sidm+POX/jOSr7hxrm5kivlutu
NhHVMUBZEk23013cI7A2hdZGPdVtqchnlnfz0t8ITTRLhDWD6Bqo0uUOrnZNcWfdlOYLKUPEu5GB
6/mA5dI0zc7J47UrA1a9lB6KCCajb5tdFNz7pEdxu7xPjjCAsmm1A/lWD4HTitKxnJVT2BtUxu1g
6xwY4mSSvuF0sMGkFsvaSYuD45/nRemvXR7VshCnY0yJbxeSt5bG5sCxhlPHBkuJ038NUGgPdvZA
sGNP1nbdwFKMTGQCk/FG2H/BjppTkOu2YqtkPYnQgKrNjChgVguMQpWOeDZ0C7OW/CgDmF1FD5un
Urai4B9OQeVljdDveHmYGZadE+pdFfRDMSoIkjF/jn99+GIt5TssfkxAkKuCNG+dHsRLMNoXqxAR
wlR5NmwEKbTHKfejTlVXchmEKQalqWeXdirwQkEJ2xrvP5HS6kGdea1eifAebkS9zUE0VTl8ktEo
w/8CBRf7UqY4VGxcSsiMSP/08KwvpG+Nyd1pLdPOUZ9SsSDCgTzsjBq29XOOtkbQHvqDL6jaO6Id
bzKUxgy+PVrlhr3bRYSzBHSvzwKYtTh+khf1o38ZP9Yronp1gCdIABNWQGTIirSpH0fHk3QJjDbS
a7ijwU0Cl5eS2N3mKj50ECXCmH3RGMQwpbjWgq94i3sBpOGehQc4YwCfDxiVbNpJ7Q56AC786CQJ
HjtvyX3kw7OWrlCxvZV8pkZmTL8xkjpmxIFbvsI07ci9YMWTk87+6wk/zR+9L1lcJ7i6lge1+RU2
UW+uFDSgXb/+u/s7uL74/bpZeBj6R86S1Zy71unGMAM4YfTz6srw7ii8yoLeW2pi/iyGuA5faa/Q
YbYA/Qq8fkolxuIa+dempNFmPN0H2jiml5P362PjwbuR6utAUq70lRdyWyWHWY8otSE7iukk5m+K
yI8eNMmtyUS9Wd5CMVfwEir9nVbT0YMCCgUOnR9k49p0PFKzVbqdKXvUlfn+tBHpYqRosIJ4zGKM
VwQGU72a2nMN2NXrf3IFWBCqQyAgnpJbvHmqo+7HSqJneg1DJxEkViOctpd1fwEsOiJwtE+sqFtx
0c+8gsN4TVvt+IZ9nymsIrHkjwuweUBaB1LEoCo6SrQN/QFc8rw/ecxIF2Vh00EV1/9QROTeyzGY
RRaD9WhZDfSzDe7t+eKroyhptow1ESNeX6a/kgH5wZ28gRkzHl0l0ix9oPVnBiNfFvnOo4dWuKmY
ls4XrMFZ9bSRiK9uCSJuwO6G1lQpFhI+LtDtG44gUCcvyy31ZqdePABIB+c4b9E2+ZasDQIWi6Bo
NpjbTG/RrKRqbuDpgmfa/73OOBpYs0/YxyTiJtzQUqb6PQqQKs5UCUrxs82TAftwfcKqksu6CMHX
b2p84UpWsI/yEx5Z5CTHax9nczfezLwwJ2cvAAFuKY1TaOxVBiXBdwdFJsQmMSBe4mCgW/TvYl33
lYR5nHI05L8FA+buUdwkTwRB6UQr6LN4dBkOLud0F+k1FsTs5167fvFBvRSWAIl9WFmiQaKZD4SI
fHniRp6cQtJ//LiUo6GTkcRHyRxEtgdPH0Ses7GlZaJh8qsVO1fj+831YBWG2iHt+V9V0iA5GsRG
DpnD8iRQ3+SNVKeXj5yQpMUg4GQW5WNuncfJfWHEasR/lT64nyfkaIfZPAvLgOhDuLp6diS89CAH
9UBPXZCJcoEpKREI6N0ZqaWWUnW1XbClo7X7NYYtAeohTiaT33OM4W8HJ78vYrHpcnagzMNUiCqy
5LscjJlbehZ9snFz+ka+VLFBK5fnH7Mkez2JkRqf8SXLGIvlTI3L7jMKwYfyo9biAqi6qIx8bCfM
KDNm5W+OqwwJGdfXYQeQfA8E2a+OzGZpA3Ml1PC3HlME1+3tQeZ8TSXcW2R3fmZRvQWlPX+VDCOx
dRnipGvrv4NEDcjvjVD3EswhKvSWF7A9nFgircxfkaMN1nFyj3KfVM2WcsmAUUPZY0BZx1m8dhiT
bn0BZJH2TMC0J8oiGBvHO3KmHLbtvCAYtNNN8jBkhpG5V91SDohHxpE9KmHbDFzLhfx1SeDTnIJD
+CupXFiw7N6LTi4wrA2J2sNR0sg3U8v865YGpe4k1MPmSaswI6TZfHddU5bffU2JyhSMETVq2F+Q
rYBuejQBay9RMwOTzxtoc6epE0k0OLg0RPH3YFBv9b+PTpJ08IzUki0fm2NRyz/3/04LFWHH8gla
S0eiIByKwkCG6Xgd2b4Nhs61MNz9w8Eg7Wf1sNs8sZyy/0JjuZwJ/FO9WopjvK0Z/ykJZXae0MO9
xS5/T7MRckBp8JMqPPfddtlyg+AZZd71KcoFagXJQEuiCz5CF13bwONlBL5TWS9b8TltD2i7+CUK
4n1LCjjm/C6HcPSg0oYv/bErGTvdfQoQr6/dv/QULuVOaq6Ya1Ig/lbi3STFaH9Rc49sPhoTggM+
FFyh/vB5Lgw4qvASPeg2u7qMftsNlKknybgDRKJXtmq6gVai4054Sf8nXbMrv6MtgRYeg3qbiSVB
piSR+rFVMlS1YBgcagkD25yJAKlRdUwMvlp0HV/Wgwc02AXNr376a5UTElU5s+u0K0QGSisq7zsm
ehSZg5r0B9ANGoMKj1PGpQRPrqC/m8tYXlgNszE3uofUxx6nKlM8ngvhLoEgC8q1XSNkiawSuGMd
1FzThM75/wdYiDzpTvbsLVfbt4L/mP67BWdlXZpnuqaDspDwwI461vCwtwVjaIgWHTEGBXd8X+bn
h/Fvsr7H+ZaK2Y0btaW8Bnk+I2O9/StWdLU1q5ZPwHAvwl14iFP3skqun7rhmj1Dm47oCF6wfAf3
aXizLpAcdnDjKo1xxw7wsWZr01iHOih5FKiloXOxcF138e5eBJMr5XRSOMMJ+E4eQFJMhSOKI9++
kaNwuw9WJcTY0bCe3yuPF44meITVmRgldp58TYcupGbNpXgzxQc/iX+ooJJK9yMps/JcQ3ReqnNV
gYh9fRw/MVvhU8iOOAaNcX6lG5avcJwAZLSv6hxft3mtBDvU92BsAncoHO+bFHsXXkVGXc8E1rva
HdAuX2hM2s896YhDWWgB8tgAAC7BuzYTiJ8yHClQQzHXsk3RRikbC+UnjBHK1+OeV7TF2UOI0iox
AtPNWpxPyIWk+yLA+vH+adNPc37utxzycnZHqcx/ItZp4CLQWH4S6thd0piS5hMcmsLZpbz60z1L
xObA1qQsEGkAw49Oz5ODYZRfJNiY087PC6Z2ZAOSdA9nrpVdfiEcOTgSZNUzbodR0PCRtKv0Bx7z
bMYON87Pw/v6LY3TmDEKwwN9nHDQQ48+ox/o7PqmyzPx0T5IKR9Qfhd4+Zf1TpUPOS5WXJhy4voN
sGHGNxVpigr1s9Uiz8b0PO2iAAk2Yqd37y4gacFf9vQYcHHbfoxrLDpWTCF8G35kJtE0c8MPuJGW
MqQcmL+d9+rEUEZ9yXXj9FETCszfA0b4x7nWDC+X5HlQEVeAKAEc6dOMqp3fDr9mjsLSeuIUPC/r
Z9N5f0el/sIj8d4RzXMtTXzACwO9LStgrlpLEMJRL7ew4FimZ9VbgcnjOy6HphyeA0sSQj8neiEf
fFKjnVcVS6MUmXphSPOX2s+4XplngJjL7GCCZ2ZtKGvwrlyYPU5Zuot0O+cx0yPkbdUKqlI7iXR3
IzRdCQi5m3ggXeTZi6pS14QG9ArK3b+fi6adBCpcz6J4lP2Y6rZ1vWRJJYd5/DX2BXeJWax+m7sF
4+PheJt46LM1RABjT5EnYXe3Ez88DDGOgkbvTgzvoNVKB+0+Z84r2HSqNERYToKi8oEDzvKKIbvo
A+r3+t3hs+ETPmUDrGxHmLNJ1hlI0VDTTDfZtRm9IdHCPfv0LR7NDhH1yTw0BM1qSXnS+yz7sYL9
OoUZsvBmk7j0kqXHGrDa/L2cw7LwtkcTISaKs/eEmSHr8NLdNf3Cu4t3YjV6frBFy/JvX1KVdi3Z
6Db1rcCGT07qftOHJdK8W+j58hy3wATG81eTjvX5kEXn4SDpJl/vo5Y70IMRDoNRFyEegISdQ31M
D+8nvQS2jZwD9eJFy7U/yRY2Q+aMpqljiM5GDZXcpUVlfKrIZwZUFlD1+WIAXeFFTe2KpcxLKhl4
8edz0lIj3pj5kRR0N/9dQVBazfw1Pw4mSxzKtyeC55zUUkMlE3nUA357NjIGGfF/HTihkIihICdu
05QdU4P0qZnLC5vB9rZYtbnRkJaiMJwh3gAJ6Q2bGUwCNQV6Vyz791Sq3TJmOwMFOGtIBFv2cep3
w6sRVlJPMIC6sBnRb2CEZ+MzLuVhKy3Av8L58XLjcTebtK4/MdgN+XUXuI0RF7nh9k79KRUSeATh
RcbWvnwdI0lsfHmHCQBr3qzg/29YpnJndmDjascFaXgHZf8reh8lSo7TBODAqmjnxciQoWG0D0GN
9bZZmzJK9JZwnTbZgDYg7XWMATGMIFzQ4s2tkSaJ6ap9q2sgni9/3oM75q8usFSyWzLxWyUcTYsg
f4s0DYkKfSYIAkOkX3uKlXPG0e74dQ2vMIdB1i57xQGEi0DsyWm4F9a8KNoOCz3gtioJXmSUem94
d8jht+lMMO2f5DujrINLMG7dFbL4RL8FOLRojl859y3oKlKchKPFV4PMTZKuqzhHWqRtVpwuAkAf
EZ5gkbUczcQF9NNLXFj0r9tSV5hPzTNSET1TGhSzl0NK4AMo4oMM33xpPVycQSgIONBiIESoLJ8H
iK59blMc+IyigTidtSNtF+KmAUzG5Oo+coNUzzknN3zY27rWlpWDJ6Yy2+HEH6X7o0xDWab0QDqQ
6WLUf/YgI+0EJtpbp3BhgOJXeMgrdVWvRE6eV8KFXNLhg4AMbJZL7V9zGWrHxwN5Y0XT+BQo1J96
g5yYpvM6Wxbp5Pb7TG4tV4g7Wj18qKne5eWOhB5jUbRMf+V3JYjAcw62daf0y6G9RIjKoQ7aH3tz
TwI9rgL/DlZ8e2d07A69sm8miy0BRgXjcU7z5DpKRyky8koiy3MesWbEGFwVeRnj83XVyEa222s5
LlKtTrpj0SwIP04y/NUZMEbneiam8qq9cSDgt1piH6An5lNo9GBv8vHzNKG+j4yAxcpkpmQ5DfTl
4EgfSG7Ka7BPKniBrSQKSLTRhYMF8r52UqA8MEdgiimtJ3fZFqEE1GO/pmBPC3FWL4ty9bZyFjlN
KdFWU9D72hH86ojXQXlMWGKJ+L8uIztW3PhBgxaV8nBk201WGxufM/rkh4A+we7W5Ac0k/PAqAWB
S+FV6Wnuu1v59zhAPwaqLHCOSyrsTOfufitNJewKPR9Nmh0HGC8GipCZm9HXxp8lJlKv4Umlq0Nj
Pg8esxJdVDWgBWuM4TrmdhCXB/zztgjxxeF+3BxQcvUKg16IRzgUX0BeSYowe+DfdS3FZ3Y/3xky
tuy0ETihiyVdvR5hZaNbiciENC0Oc2pHh6xBGpPNPrFUiB3RjZUKdtVRuMdzdYLSdeDIh2Vhwczk
43lb7BCZ41MrZrameUYw748fQTIUTXYwiIweXCvnImDAA8ntXHSlA39TVvQKf9VwEnZiBhi4+wfb
NvsIz+cFZTZ4KML+8YPIXS3jp1JXuHyX84FfSg3ZRkjERW3T1gipXDuMCPJYEdiMuFkpX6xoA5Rq
s+0kYthFj50lwYELum45+MIuT0t9BBEvRlfgviQK/+C6SoyeWSYVcs3Uev4QEJD5gQbF6EVbtCNX
45muGOWvyvmeT4AyqV8wKCla41CXVGiso0GLhAYPoi1f6eye9TVfKC+b9Jbj2fAAFGF5zNBEqxAj
ShWhKsQSEvvlBXg10rmOj1gXBrZIesRMgb6XKLFllrYmVsDVITleO7LQcXy03acthi3tZkB7leIk
z/UmRmnCFLXRheN9iNMHqmK3YybUFNWL48xKiAbK1TAqxFOZJHD8ALz909tcEM6lOHGMvlukudGX
FqmjlHTYFL+CThpJmaJWpA/3h8nCsX1tpWK/CRPg6wIFDQQ5uAGFlPskohXYLvzFx712/oNW3pxl
gAfd67MUvB+sAD/+xoxBajXx0uemd8cwbOszh+ath4zqlGM+8vjmTNU4MjLPEgyUmjm844hHTxxX
LNrjKQU7M+6MjDa+mxoigP84Cn4NGUyVSilg8yajCgoelBJKjYVhl2EFi1/kO5oSMe7fdHtJvBRE
GZ2R1OZR6c4ScSywqBCENHwZ3mtrcljMM0QoE+4TR1Q1+wKpC+u8yW5h2BethHPJhwfWUipoHH8x
SoM8KFFg7xyrZhWc1zKTDaKEgvOid76Dsd1DfewwaPW/+zKGpXTGuTxMVyajimTOEI7CLLIinEr+
iWqEVnPcWCfNnc70DbtYeYGOvQJRc+B/wcdjTCUVgI+NoraoHL1nIT4+TiadoMgBkzrUPWD0fikj
uNxt5y/8CEiFmTvHsYfReGUuAsKeTOlbUw8ql5afIkgiYI6WI1wSPIn6kGTYpUN1QnncvmJy5Bbh
QaroA2F9flF2uB4va7mveKMg55WFVOzxjW3BRBoXsfHIa1eykWwITxVdR3TsRaXQP/7T+Kexo3dY
DHud+ZxNlCb/yw/Ng9L+fi0yEAFS07KyME/+KhtqEl/f5BsO9Y9br9kgvvuQG1r6qvRzxjnTxQCp
khu6jr4IVE2YCTw/kUDwY9T+MuVhNrImvrhpWqKq7dzZqRy+y24NylXnvtjefqTpW8Cn2lb+HHrq
V2IVcmj9R0gKF+wJZHFNTzbGeAK52orZe8uXBzB3AVM2Iqk0JgyZZGi2aZw0LyyHt1s6Vo4yuCzN
AjONTXsYEtvpKL7aFEyLoAv9MIlTREP+XfuknFT37g7fwGtEvZ9PwzAkEhT/tNzSx56dFbDge6QD
I+u+yD/gJ9m+wDfZogvMCvEpgajlcvyY5SYR7lbn7xZB6ZO8sMFDbimoVZSGbNds60dIahqv1qgU
Gm4tlu5UfZ+IzYHGI+LN3MhSu7jbe+VZEU9PDIvlZDrnMNIGGKwhWWF7bIzJ1zY7js2Sya95F6zB
qiQE8lc5EsU1NZ6p+BKkjjLsIBbKzoO4oxDXhXECzOo2DIfKMWu/AVzzf9LE3xk01MlmjLEXFwMi
AdAv8if6RU/z3nFfo/T5vyAoqEhsWC4JICj81wMmJnGaPrH/ZTNJJE5b4zhyqkdhNXINzFPuC82O
+wtUI2B3+s4cXXn/4T+C5NhbgI79Qw6r3CZEuK3Wvttxe0MO8oXTlGlnyLJLebsFLMzrUw5JMv8l
KpFse/xSAzOxLrvIgCl61J/5BHJrCRiVipDLZevzMUkpSrW+guqQjAtRJhmZa/EqrW+Co+gal9hR
/Rbq2PD9U316/uuLL2LqUBm7p0/I+gRdnq2KB1YYZ2VchqWDKGgqK1fzQJa09Jsy+IMK8PZUoF3e
knk1ocWObZb/F3AbYBlTDTQD10JhD9d0rLeTGXOfI/kPSaCH2bIZWDHUuA9DtN9/q8H2CfMQ/m+x
dMBuHkq/ROlrUncoYIrB3LSrZ2JSUNCv5v1I//0qkar3tMc0YcID84K9L8R+p8XqTjlADb952yPU
9mZS13arRab1ghz6Rap/2iG09VUdZieYySNe7pcEfFeTrqgajJsdfZ48reNruTRA2posqyD+LRXZ
nnwaKog155pHQcLKgxCDAT1ntpqaLA3XsIY5r3xU0Gm0xzfU7ZxADQyzgJQfzoUcod4fukVN7myQ
Cx5/2yeCVyNOB3qXL3F6re/a9W6cMkuZFU4SPO1Kb/KbwFiH0x7hJV2eXa/MCKfn92460YRfbeBX
NDwft6xJLdq8GVm9+wT/SD7jBFBMPtQWBpqs+GicaOYCkZLPJWJ2OtcBlzRtdEe5+VSzm8KCeIyI
tk+EHmjQ2pR2q8rZ7v9Bba18mo36CyTr3AjBuB+bxWx7L9l6RSV0mj3mPCHIR7Gv6dFmuTP5H+pM
Wmoh72Mze78NLOnIRX8tim+Ga59nEax/L72y/tz7SdXoFP9e5+NmJX/AbnfEY8/ckslj68ay1dfL
K4SMbWWt3Eu+e3S4iC51PNjJZM3WzQmSqgZOVIwfWqFCap7S93nd4ZIbwxJpCQ0td86nNvEzt+gk
KIW1QduSU1LyxAw+1kuilkCtO8jI/QtVEyCgAiYgehIQq2svVRPlKbbwvP7Cz1jyCYf8HoPg9H72
tau9PyE1m+Ur0TyuPtzDWjq/W5zMw3RivniE67MIldx84741rk2/LNyggpB0YFqkuE8y5Vt1HxH4
Z++8S01FaApArNJMvqS36nuceeHE2X5i4X+cnXZ32ZmCW5RHtrXm3eCkXEKVQsokecpH+hkQM5fD
LO/g22emc1Pt+9tXmOL77huJu6+MwFUU1HGVALOBCitULfYWR5iD7+JcgVYk381Rl/rEPajjpXzq
1wbLVAol1rPnYAmIq+vMO5V4yCxuXyjUGPfMMoq6M9Z7J+S+H/t8B9Ngr1F7ZUTgGhadJCVrm1cb
FlQeE/eqwC3qgcIp0XLY0o5gUc1N7BDIc2cVumlKvQ1pSVKMHPUrBsTwqAGQZQ1PMALUEh1wyGHs
DFMYmaVjdiAbgnKvNXZ+U+8S+31KxRA5sJ0yKD6RarTxOkVX6ODujXuFBITXDKLuBRmbIwm5oAKW
QRQF5ruRpxfypFt/1XQh5gFJu/fqaOG53NCbA2bpzy/ZimXKtvUm4fNktNkaKWOrGcaKfbHAzkhj
+thhrUOFNifIwDwhofQc3wtg45UPxQYxhwu57Wc7A8G2wCHDcXHt7zHR/RnN8d8373AyV+CuoLso
KswAPca5NNYa8x+dkJpJ4XbZ7Sn6m7l/iXECLO2ltNaL+2qfCUJe8gV4IpP8wU6ugP24ji40g+QL
NC5NXSLDGVylBiC+jMd7zjLdF75fyOQWEL+LiS2WVx0Xr0GKskz7J7Y51PcRHEi4sZgrOYUUdy3a
BXxKwOrUPUFo7UF7hYUjJrsyORTgg4bTEc9YB1Tex6bqCzh5H9xTrSRhO1e/VVwDw17oFM1PAchZ
C84dOpUBgJ6phJOaevqB1GZZ4MC7dO4P9tZkdALhGlbFB8/Tg/Ha9u+bcv7X47BPTt0y78GCTKWf
Xx7L1IJCIoaDyDS2yQKu7x6SAfzwGyH+lTipxv0H1y+kAHqdcgdqL/Ks6UEn9NNZ4lWRbo5h0aNK
ZXX+FXpPmq/zm190QxZh+cI/7x2K7VITOIBM8Fagvq8VuPZ04qbFM8cevDoRHkFbKCA9mNh3vWTM
m6ZCPOW6zQ6QOJ1OjKKCwLOgv+agBi4KJzPZs1DRQVipZS4KRvzpBit3EfbyaWrD3Ff3PQP49GGq
J4N1FfQ4LPR13h6XZti7TxgAcnw2omD1mfHrGVjABZ7tK4Q72asimnZi4nRAf74c4Zt1PMdwCdqm
6g6Bl+L7Tqzxc4AXp1u3hyMzImGSJWY8WAUhVrdf3gkV9RaX2HmQ0APNNlH1RDxKofnJHVj3+Akm
NjYfpvi4h9gX/wx+Y3YINt/WxNAoctCYiRkWK7Ubsh9+2BWWC3agsqAbxaf1uW1MZIvqKWsejJl3
pfGZCRb2CP5+npxvJfQUHj4dvPmFRFGUCX3NG6CwtorPytc3Zn0mnaUHlp9uPUgzLNLh84Vl0Dum
Qzeuji8RMNZN+7lm0Or2hh3GYCjeirdL/f9XSgUm1o7ipHV8Vb8HrkYCMjBx5pTfLInR6UpJB8XM
aqy7B0oNnNDlIwlimGtjplAagJATvLDtBXid+38AFMagXlfd7CkBq1pl/krBFIJuccke8eoKI1T0
JW6z/fJapCESVENAq9TNR8yobTlzZEeyd2oJpEzMuIpNYTxfY6W2H2KLWHJHNFobcR+0gImYugIM
GYL1dhFJUavfXNQ2CZ2/q2REF1KZYUYEVAjTMtI1UbT/GPjI6PORePhZURMhY1QGYQdMWt/D3YlN
nigz9BsZyzT2f661CTfQMzAfrHfIiIp85xyJp389V1ja6W3X5j1HJXD3+DSOUezNMtdHpqKauCcq
dtQmJEHHOpeLW1HrDQ99LkFRVKpnI6xmv7VH1PoZS5thJyhy7yQZLrLK5VyjlyLT4WMnqTTB30ro
IPkC9QtmK80lPt55B3E3sImYZ7NWAqdrVHuSmwjANFk4pxSGuQJ6R56jZNLE6tp+sa6Y7Ls9FKhi
Znaxh/BO4rKvRmAhxh5sDfW802Yc6PlZxoQFdq8bgafi6WK7sFt8Oifzem2qAKBcwBlFm58HTFQB
RZLI56T4M4uwkL4jny5fjczRhNYmLSpvGGkumkdzWWxWLkWn7fjEIKJ6RNj+TrXs62N4eSr95EEp
zqh1UbHCn0cNYqDLUaHd2cld85wyyxFLxyW2OEX4F3E622Wwl0GeAnG3ZVd6YLuoAiqjoxrWgyPO
iK5IV2sNAZul99tRGdD5OXZ7l3nNjQIWJja6IDNwT7cMllAe/h7Aq2VuTJJMb7lvM9hAbBpVV+uI
28YTp39qiw9wXqkwKfNGsB7rcHmBRenvN8FKKPDG1Vgd/fzzr6F2OlhzkMBFKS06hF4lKHZpDH76
Z214MzFHKhq9JKfiX2iV/EqESNxD1N+c7JxtWvrNsoAJS2aaNgHCgR+0jfOuibaa1Nf3DCnr79uu
UI09CW5090RlrKbnIZGhJT6VWVj1UVQwh8q1GTMdWHCuASLjwGUqkReg678sZ5N4eoWVpEg4jIsZ
tmwJd8N+Rd/3fzkKgusM4DzesZkNdT6gkg06pKHKRnqblBaNCrzH1rTqGTck7+bbGKS5Un75KtD2
6RWMjWsj9JCDcSwjNaGBfeJT34bToC5QKIiHaPWH8kyH8YBQ+4RoM1opfyd43CPPZmqAVAHgNwQt
cPJkoGXHlvBknhGcC6d0cMq+Uhi9jkVL5fXOzjNUu/M33f87OEs547OyPCoaKWnM7TNP3fK+/aAD
OhDjvDtmCS+GmQIkGJ/cf9YdyujGhWvo13az+SNU/6UdtesjVMdp73ZIwI1VEtKyrimxWzEiy/yT
Ce9zzL7dvXkBFdELxbQ0+b92PkNW751eYGdJclM0o4as2shUYZBnhpG8ICdLEbR2OnzDub61hX4g
qDBxTdMFXEccS29hizisuFO9rGdw4pONUg2le0guZvpxQGc1NahE+Q4dvA5LjROQb7WosbngCkBb
Cwdm88dl07qVhxNgUrK7FLwj1B+pLkN2GxgvKXpF3MSrFLbriKUfrxCojKqah+UWW3KXmD7nFavY
SLHRzNJ16ZhdoLRrZdIiWm5usbjFeXzwsblzyFoFiC/L7BVOKMrZWe7YruBtTX1tMjQx1v8GHSbM
IQFWNyll12avRjN9ZZ+ClYrPb+kq+gkvLxkEacRHIa4WyRW2qDAwLNMANYyNQq4B7l7iiiSuNM7A
Xj/Fy5PCnPLXH+bXUAm1D0W3/AEYirzncFGMxzvZ8tVeOwRQX99fwR0vfnPWc3oEUnj5Hq/aXf+a
if66pc8c4H+4JI86giSYhIBvsSWGBriHznl86WGra6uqOJXgOvLBeNMij7YZSC3X4ipZuqafKdMl
fXO0xIxup1cVPuDfiej0SFBjI30sn9rZPwKRFBdTrNcqeWlh9YvAqzJmHSt89nLMEWt34gofsza7
W0FOH6crJApNsv6G6Sm8V0ulHCJAJqMhWt12ajBkKbO9+lf21vPsx0KqAxa1HubbZweHYJ6r4FAW
x82zMt1hM5Ba1g64vrqo5PUxgv0WLeWV+bLMuC2fKg6WLxnnqlc9VTrh5u6Z8I4//X1gqOkXgeVz
YeeI2jvA6sjExKiPTiyugsZDbezCW4lNu+TAJWJqT5E0LGCQR1WrO/16g4c/gBYVanJ2T/ycfZpx
HK7LUIOAW+/ae1h6wcv2IY+1C5XfYat7XiRqoGftx7NchGO15UT8FOOkXJncSs7HARsNlsRg637+
mw0mbaRfUpPQg/E7pH2QCq9maY6qooPHM4mZyL+cb8fBOdnVyN5KNO4fMtMXaiLsVszhJlWJ02bT
yRsuqAbQJh24IunmUgMODeD4mPHTwuA62sbVxrwsCJAI0fMZYK0YGrEnCcc6K8EEawo71UPgGGHr
nF/6V9Zlq7vfKVCkxTXlLD0lmTfG4wKLJfpDcBtbvbMSYbUzSpXVTm6F+9anwS4HdmyBALCDuL9F
6OLKKdM/reYUHcDKUUxTsOXYOmjeiLN0Jf0DNEU6cXKmdndaoWgLTpUHiXHFaCFZROID6AoWlKdm
BUi3avwyziNkIhJdELlmYaTR5AGOhFAu4vjKK8Vf30OxftwYJUP+OJtt3D3TACqs+T2e3i2f5iVd
GD2AUNq8kHFTskoy8Zz4596AkuFAnTJJWxvpPVDfaTDgBP8PbEIiznbcRRJKLzzKbA9OUIjdkUUh
LNumn7rzEtyBXrQBgTnf0PBJb2ZTnh696nOIy0dWBeLB1259Cts+8yiEHaEcV3PDJMVIZ0oz7L9F
62SYIfBQuGDw+7WUT0c/8wmI+oQc/S42wQRSJ8UbfQ3NugFX3pc32mf+pCt+934QO5ZsXwtC6TUb
VB5uKV7N3HQqbFSWjQRXarB7wCzqDvlkrZ8WkfvROmb/FDBYnYo4tNTBde9PFUTOdJ6MG7KM+zqY
5A+4/xZSzCnYcL/OrikJM+Y6iRLsTeXDMCaLR0OQeLdrPbNVQRG3kP3x75HueLqkRld+sW+PGMAy
60jAkKjAK64tcoueB9lc7gd5Guwe1T3tAzFIV+m3oKlamgL1u0GDsKOVRgGee8fwZhjOc9gWC8PT
RlkLtQY9WfW1sMM4NXrFA1D1xffp+pM9gEcbkOUjq5SZWExVB2HKMsQ78+yjogXWJ3ab0BsHVZHd
ShNMZzmTlHLN4KyKSXf0FeAZI2MRdYnJhlZ3X9mU5JMgW0gVkRrJadpDUWqjLSVcXzlagNUyrLLw
e6Koq4E7mphHflUXcqkzptFRAIFjD2AYQ2vY1AKCx8CYaWyqT+s8V5HK9C+NrJ/ZJNtgge6R6T0n
5u81+sblbrPGyKjBFnLrlFxgmtkoyUnCHtsYeW5fLWWu3pvL0lkYyqdSNGs/YWEwZyuvVIVYhUDP
tsLQbZiUpahtu5H/l6GuqP4oFaQKI9yLEF8Do1gCa1W4axWdFrOExkKtR8foahr+HDKs+c26SrI9
yt7clHWXhfn2wY9gOkuihb3gx70npcNF5/rkxNFxsEh8orc9mHybznt75NTsHTu0ZFGhqZy2xx9I
PB5ojbb0eNz6hsTXOX2VtRd9kN3eKXsQkPNRIpLS+YFBd+j/J9nDhzdzRCNihYnEonQ8+ZRTiIQd
x2/IiYQGeDX3+nMqk11dXgPIUe6ek3c819lLwUaG2/p+4EFP7ANNRJehnf3cm3txSXCPtVyqnpbv
YyOuR2FN3Z8I8V7gxDvQDGYkZbL1dq5lG1Kep0LTGHse+p3yAzZFU83/CWwTaLGmcad5T0KrMrD7
1dqALtw1rhETrdCat3dhjpJ0w5cwvgKeYuvJo6FFzUac+I42mMWLmszrS5iNJSZ6RNr0swSaBBVU
eOOOLR9qKvBSkmsmsDaiT7ih7g+O2G+wu7c8cX68MdwQSCjqvWr5UdYa1LzvBR1NFzL0SAnGzZNl
9wdEG9r8u9AOFr2z/PHujeLyTkjfhAq0hQxopzjj9kKkbSBUs/UnxPHaCi8DDk3HVpJDpn1y0UaR
CixRhPel7w9mQL3LRCWU51ed4PSugaqZlMq1C9NGYQyA/Nl+fv8x4yCIx4SbiYSpYq+ycs9l5RIn
OTWuPoUkXe4YnbRK4uBkln6tp9OBMSLQPar3CNRKcjaUwBQ9Ro61UinSFvKPrkNBtx5l6LcPL1Dz
w8fUEQ4E6ZTmS+j09AWQtJ5XwUrlIdrVCK+swKANCx1iKcr6RNvxIPEsj0OhYNG7PluyLXu19b0I
QKC22pKBfo4eVc2CX7pXp83M3pTB/RvUyeWvwF3N+KGQPiuDebtuR7r4GF71ANgV6epcWtzVYxJT
MKaaGLZOrm3ZF0C4M6FxuOGHXkULRlE6j409LI9RJ1bwjEmy6ZpTTF6QjC7v+RUCqLPJiSI9vudf
Pe0XFXaVKsblExIAK6jO9b/0eERgEz/Sl6RjSIUge39jHggB9iEAFZAlhvJe/4RmCX6smxSa787O
7mJGX/dPdOL/zqJumYqH98yX32ToRe5xcT5D/o5c1l+MJCVJ7HWjkBSB0s8SCEe5Q0M/4qabZ69D
/WsVBIzYphI85rReZFKB6QqPy0/B0wUPNTZjTOHQi9GUY4vVrw7nkgDmTtJCee6LhiZd10NjrNCx
dQ/hmg9G7uElUJqVeeLVant6utx1NH+YTd+MXamvATusYsqsxkloiqP4jZg4g7Wk4dwdCPF9C9Mh
P7j5yFauk5XbG8NzGjJSIkhur1t3kBmwwXdocnSoLNwH41rekf9giiYW6qR6YYwvPpIC4FFvd/ab
N88lZoHDUsn4R4Atqo/McOBC3u7hKCOykwLxMpGr+hRRcKE/1yVHz295MKBDq7l/vDsSlEysJMyY
oHr3qe8NUwCDNA65DmnSUcBtUE+Mfw4hYnHYWk8AH0mlH8XOFtt4ciWoCY9Q+1HgIwQwBDl89lE6
1gNKy5zgy9MDtdJF5DZ0CKt0bOK0Egf+ZggjPlYmImtM9l3mzg7nK95Va9QWDJXSAxxNzW+Y/wel
6Ersyokkm+JdKdogaIO9VwtNmxqD/oq8Mp8g6G6vhGQUlgCpcKu2blwPlxbEQZl8h3NLBxvpbzOH
aDZ5SjKVKodrcs833+iYmSQ8M/zv/ezYXOfoR485ROOXYynPtgp3pHf46120fGA7SFbp8Ypwp0G+
WB3ou2U9uaxywVI28dPonCJVpFamX9wGpnTqnXl+bPuaFT/zpnm4uDLdYAEwbYc1NySz/L0eehxD
hMyQFAoSOCBVip6Kauxs8/rMxpDbq/tCyxTbOVe+zVGzpMnEo22EHxcuZE7BoUjxldFCH0Dj1V/z
RcvErIztZN5xVOBcpezUMfLgjzuzt2mVJFxkv+0C+vNtyT144SG/mwh3zmTsC7N4CjGEhx+XE7Fe
uJuWxGzCcZrMaFdBTq6QMLfLCLfnx+ZZEH/uA9EazMUwwNCuIV6MlchcPiIhwLyWB1UZejFFFh0/
43KfRdEjcITaIJlAE5d7MLAuXXxGxeexht5zVeKEE3XH1x/6DmJhjV7TOudsfP3ss6ZwQZ+cTyA5
+LDg5fKCKjEgfM1VyDpgNCMqved9zg+9heuihbF+Ex4mocm8kJVGWW0jwAOX6MtCpu2PcT4cuxhz
WSIuAU+nzqrq1cdPns33AkThbDZRgJiMuqSdb+di3tCdI52BkranSJK1/24UHqXdRny1Bn2++ZLE
prHCiVRgyLOG+YgH9FVt68N+9Y9kOUe1YmV5phWZUgQ8StcKypIMO2jiDRa/4p9soaYscUfiTIR+
rnHqBxLkCgR6xYlTdS9jwMYcy2GX/f/tC+77o3pUA103WwAac9c9918IygeMIvG3CjuFtHGDvUuH
6hrASRuC73HUkdVZVJATZ9iFDsyXXQ0LnbxxVhv/Hv08/UMpZ/fx21OdD0sX5T8RIVsl5X/BhAaS
y15kFjpGQMOuZ9Av43FuHQmR2itDeHYLJQbH5RPkz0O9UCXqB9YxqZ5TwJYFDL70O4g4pgtWNye1
9dKOSa3YjfLFXUEBq54dfZB+zC5vOD+t2oRGtFM5Thd9vII767zNisO5BTJGRyjSPyAuQxUF4f+x
lTE0hhT+Aj6UENHF8s59dLuKOgNugkcT+1HHaYGCHuJ38EgvahyDq1Hfb4BY2Gwm/BmF6FRK4fFf
uWhsbXAlCg6cBnesivGU8RSBbf+8C44jaCY0twgMIqw53r/pYI7sqQsHcikgfcFBsoIv9w3jFf/i
X+0DZtzuUUReX2MsqrMBGwzX8hRyq0vyh7kfIZzXN8f2OJRUIk0eRzF50joS99PNZgsTnC5CyrUJ
46rG2/rVvxMbEg+BigotTpaIAd988DLrypJ+tRX+jHvhjVJsEsV5VYhA6i3nKlk/1u8acJMg2sZE
TcAamT/yLkY+4L42rBqUfGuvn9ZZLp/UjjcJP80X+6nwWgCekFyf/tJZ7F1PkT/jcD/gQfDMqVrX
SSk4Z6GEtKMPUHpHYRQBQddEiFklnfaMLSPHa+kEITW7vJrjKWFQgxxyAoO1JBiBMgm1qW1Lr05N
r9sNWxveg/TeMORo1PVqCcYYGL5jPgLhSCB0ruUyL9fqS97WWfsdYnSEriCYDlZrubE6nFw8A2C9
IlajIRJpnO8qnsL42D6BY+G8w6Rv84XUDHNBo0CeMTWHwjEonPNtaBjqzhNC4BgU4mi0xLMVlWyM
RWZgkEypctBtGiSH/Fa/Sw7gDkElMv1GzIQKn9EeHJaxYXFEVkGBVpa2rTm7crV+WiVIverG8J0V
w0Bu6JtWTxrnAwmtoT6c/jdiFGnwEVquE/WM2YoK/s0Dhf8oNcle4LndPyd9196Y6FhYDP9UJEfD
0nQ2gGSfFCEjRsrSTHOpUejukgGLdZFsYTh0CfydfuJ0PD6/hD3/KnvIq0q1wSw1w8o58MisSRm9
VaT12kYUo5/07w+YEtgkEo+eNBuQFMgjo3u530Afz+w7qBnrFd7pQW61wFbtpWfjtN9HV09JUXsX
Ybs0AcIsMeAv8RQaJdP4/5QxxfUG9VLp31092BRC+fyHllM3V2ghuMQx+iRyK/2Xhj+Y5Ggh5GO0
wHAba7/QyD2qU4UlW5pVxFDkArM8A9GF2OTgjQVT5OUpdkdp0eADQcRWgrdsHHMJ5+VekLy02Yc7
rqdfbQBiG0ir2Zxl4XNBoMqp7ePimEoqnf38NFVi09EKaZPFmbfrGjcXVRF4Yvwxf4wyrzXmetpu
LkEPfTdfCtUGdXxQq9nYurtPevQ02yjFiZs/a5pXJgrH51Sgsom/Wxhn5GDybvhgpLZW6uqrcagu
VMX8WZzg9P5Xp/s8holWEvnHeVSXwfgTVHzthguIlifauMHsgItfZid0WuIUfLd4d4EFhjlnQ7u/
vCLgshuae5wUoNTsULYUc3p7Zf7b2GVvZk99ZUKbEwuSzoRHuVx5FoOxDlkugmhJcQ3hHcDynB3L
TH8d7vy3w+zsdzm24w1qX1qYglR5iBpK3m+l8vc60aoubgQh5bUV5BAAxOvZuw4QW38TLSjsJfRO
orbecQIZyqa+lhIVhhCnEnenTyh0/uin8sTkM1eJ1hTeN35GK5vwEugqNeIhRAbLs1g8LgRRBmqg
JPg3hf+CVQH5g9jma/UOc16n1yH8TyYEqx1XudzKxWlA3Rv3HNxQB3UqsjD3PKCljxjMpzsW+7UE
sluBoZi1LgB3/Ieg0M+jWfjpFMLha0siPh6PGFNDmmXqT0nhCfyaJT5cL2ma5mHxQCEejJnWuuAG
zWRET5+sf0G0n6eyzLtvS0PsqtwNn47HxqeJ0EiR2BY/IFSfaZUnEmjYGxuI5VJSqYsIF3GtUDsz
kReCPGiWcrLI4VnTcKh7h74kbfZzleEXMOOrYcjH52odQVTb3iSuqqVgVxTjVRnac3fSWdRbwGU4
uynGQdQCVMPpf0HL8uV+TP+3IRVulOIW0kHDSYqtic/1KsC7mXAMWf7B8L1uUlS4FbTuZEZ79dfG
uAUiSlcdUekU3jFeQSmf90xPkT90PR1x5UUKSl0iyIm9Y4BokQtlspE9cixA3WH7eDNVMsHTPm9f
EAs7cetng1Z4/TIpt/Di0U3WJ8XCsYThmBrR8aMkrSHCK/U1ZE65alBQcv2bEjowbpCe5CcG7VM0
5l9uQ6NzJ247FaquhRuebBJ9P94dCK1ssZqDxyiOdRsb9mjl2ilfySosDp+EZqWmytxkiYrCjBF6
7+1xuDSn2TPnngDGQh8LJXgLHGoNmr4Hsj6LP9aMt+EPjiXx/SBmV4Qb5BPEDX0uTefbMNBUJ6aI
EfmwNqpum89OD4XSZZ1qc0r16giG5XMBgxfhsniPLKwZ1/uIMXl5N2a6mlZyxqcBjFkwdiyyBW0W
T3JFbSL/Kt6yE9JlRzVI1eccaouPc+KjTgo3/+A3QvIIBLNV8ubSHMghsQjzeNTgzw7U5knb2A+X
GSo6yYixXlcGz8JbTBhBteQm09NdjwRA/yRjRjTr5J8W7tPRjMGL/g1rgNKHz9RBxNq08+DfI6b+
iBIQcc7LGfbEE0pbZLnwV5Pkp/CkCEIDWaIAarV0lJ/woMV49GsVYyFWizQyK43X2SZDTI5Qo3+H
BQBUKwDgtoRE8kTjU79caarXLO6H7caybHFdLJfI7hOrX2esonxv2Ut+hc/toFBzWabH31ln93Ap
o4Kl3ZfMA+RXZQXQlH9aHIj4etUmWJhEOyh6SKlANp3pGIFR/AejJQL110kgTTylJAcwmgPwuZc7
p1lY1/rc5vZoWLFpoRLSpf3Nkt0Gs5Fg3v0RaxfbTszXEnSWErl+7Mp+hAVlI+TYxgybxpf5UXQL
kryU4uEaxHAyoX6xAkd0CpwjYv1tqqoU/Sz43D1RvdtrZ7eAwxbNwr26XDxkU2hCpr1FgYF7R0ap
jVT6ebXz+cv7Nae7hh3yJYJEWIPcqYSIfmK+y4/V6EyWVH9ann3y2+0XGCAc++2s1jEnW3o5jV5M
VZ/i644Ll9xwQ195cFJih9Rho/KZFBHcpXiNj4UUqEwHNB8xeR+zFmk5kcCYFgXoQ3T1k59211nW
Q+YAHKs3/DYDZMrNgB5tpwOEQ0XMrCN3/Tj76+FsH0+RZr3/8Wh3djoA7OLuAtyT6wvefR6tLgFO
o6qj4VmaAnF8JfRq+DeJnl16Ib9M/TvwwMaSCxH5TvyoFp2sfK14XhfIqbAN9pMs/NVzIxBqxpc3
uftr7mlw3S4ghsgX60rfHeHncdiuy/N2cKHn9uE2aF3QuDCivUt1H+l+iSmwZLXD9egM2P33Vsat
5V1VMeK6pY2eqC8wWytHUND6U20qo7JBsXXIJ799K7pL57LXLIz0Guo8UudHfr+0DViqUSCjDKyC
MxlpbTozK2Fs4yD5rNWBz81Ob7RqF+zW2CGBf/TzKQJ52pG0DLCwgUUVrgNNzkgCg/HE81LcqQ4h
dJLi4iuZpHOzXHxVCP4c/z+J+dUPJ/k0WOF4Ck0NrW4FwxA9qL1ji47XL2oNT6aHK3bhW+snpLh/
tPpFnhyQIphIhFkTM8vc2ehL8CXTTUSPnJXNo9xXvoH0qBK86HdUyrLZa3Ay6J9RmQpv6oAqfGi4
b8h+Vrsz/x3L+UNeIR1XLwrt+7A9XBmszyRMap1FjqKHsgnBB5DfbECT/vBVadNZCCZAKie13BbZ
U9Y1ZwfKIT6HAHjKRml57MaZYHE78c8lbTcWlqt5bXuCFm5yZen24GkOKc63LZQLmTB32yOS/gQF
BAaYlC+ZlhcVPf/1lWgRWpjlwvjyw/0HSM/NZ6diXsjnIxR+O9WB9rEuwasO7FZyEzrTmJtYLDZp
zVZTPMelNsLHYZJ0PgqpkAcBLSaZweUHWv6mgST97Hmm0ifIiNn0AxKt00RzNVenfBI3NUKheIPy
G9j5Xtbyr0KbpHd/MP3QRwi1B11fU0l8eWiiMA1lER07T4coBDEdZ8DexNB7m8tH8uhje0vT6Mzz
ODCNsOOqkdEQJ7JRiOzwE1to6hz30aD9l1pY6Bhw73jik9ZIMON/Hdj4nWI6TPlWO4rx/Y7xJnw0
dhQIvzwwZj//9BiL5XdQ4NjN9+oMuXdvjoFBQrlxhyDHkDTEhNX2YJookgNbFL0TXk9r5qf0hQYY
GHR2gunzsaBWUKo5guqZwcPR8UoRPldMSYdOEZZ3rtoQvksRT+pZwJQlOGQfuGlY+WYzxMkgjise
KUvZ5JbmKP/9YfhnKOR7g7Tvy6GGXsf+yGkKWLXk3nmtXLNeqHOIGf7gqdIBF2yMbWSPqQ+CErRI
w8sn9qgojF+ItTiaDFyjF1NUQd8uIq0fmgcvrW5BacZkqFbDJaW05TBkYPGpqAu6OkFPWJ/78eIx
7hpaXm2tBAcVXLRR6jc2cgi8jG6Fuj4/l9rTnhFCUA9eqBcKtfuSG0q/bofSZ6iQ3bxex57Vatz7
vVrILL/Fu47ff6gjCnWSd5Hd5gX3EOyYzKYxIbfRul3Ix0icyZzTGe/BjChawXf/IlM3FJdjxQEQ
ytQ4wizv2oWm+wFZ6hOa0549UojIHATKn6nx0U3UPDXhl/zkmqvnw4dyT8wHrtusl61ErT3cCnjj
uxGGM/7LRvo465gyN86L174Kf2QQh4/ZbzZPhNxYx747mPUotQx5W2dqK1wAM+n1yewJylHPBvD+
d9XXeQSRRYOFrqqWMJNuVCV1DXHU8YK2d0wQ/0UIAbCu3qsA1NrYbvWvjMfSZumZoOrtaut3SBuT
O2A1XF66Yst5ATzh7aZNA2qWL4o9GXsGu8SxutpSkRAtwqV45bz18mfoytJFKwJQ+JDr9vOx/WuG
2TVZPg8ScVMYOiXi17g/hbQBFU2A7LyfNW6JoeyypHDrpchmm8Mo8G3UTEGkACV39twZJ4qQwlNj
C6doXe/7RWiZPaPL5Pdp+w1oqbted9qpEBtZKDboqCf51iUCs6PvoEJOrPzs0Atoy99fsxUo/gG8
je66kU6X7eV+r1kot9YxN/m+yoN/sdGGaJoqonGzLzQcq8opLMPyNEfPbIPq3O94SnZohJwie4Zm
ZukVkMhkGBIU3RbBFtU302mScs9o0mS3Q8Oqbgl+KoSOScTd4cLjqKnSbEiOBuymUZ0kSiDWOxwP
7ZlFzjDWfpdtuW8O7p66BdMkwoIjSbQhngkm9Qsgn2P8ooRcne+6PVWfuvAyVLEAEHHtKHIYy8RI
bT4J7FUQZnfSOxpdjzJklkbcTTqbXpimaTggMYbk9J+E6nXwa9paLY+MEYOPC5oTMS/dJmPN7CQp
wFENqpJFPjV+3tT0Evsd9nLBWBwULOT70/pyaZmipipAhrqvMjSj8O0NfMzZGF5x2s99q7LcanAy
EjvFFmrvMRiMQ9mXwAJZ0aBmWPk7RYZEcXBsp88Aq44Mj3kK7W7upUNUi7eVeFcini8LhJ7BVzZw
1PceBSjdaq+NmUWARKgZ5ehXXNPNaX3bD7iFLln4UlcpeTwI6fNOFdb2cFKtZIIlwhVGmMcPvMDC
Rde9ocfK9s1dCg8u8qVR64npphKe50mgV+frr2UwWETqzvaeICjX8E7EL/8bn8oVKsz56klbPAzp
WhJ+j44yz6hvK3N1SOwZzqC5PwwI+6+Qwllm3GaUDwwnv4gx7xyTEo8LB9i+FtS+Fxci31mvACb8
tdXr+RHSJjFpVY6NJF7WPB8ez5kugpeP6w71OdDyjZ2qihg4WXhC/m0g8aJPwKS4p7lyuhgrUHVq
brJ0RA0Fzk1aN2wQYzfBgKKvHXS9gFYadVMrVBzqJYxrz045+GNF4BmEabNR9DDSMUDoc3hA6veP
7c+ov5e6yvVfIaftgrOTxZMIkXsM9IlyJu3SH1Yaiv2kFnrLSAUuEHl++jONltzafMqld2tBjb77
DSrQI4wTcIl6IZJWx37dh0pZwMU8obpaXlGgiVENO4C46nuy4LB1OIOU47pcp0VFDl9ukbzwAxgs
y9J/IEbYdcmmmD7uwWsyu2zmpMcT4Ep+SScpBEQpxkCIHXFJq+J7xAQRMgCJ81fE39GCKBA9eeXa
nqVmQLLi6I6u8tvqED7nNH9VIgg+jUQNZynw1Q+zBksh2hVhGz82t+Ozd2kLk8eW/d7dFaN7Pezh
FWrr+6uHB1bhP9eSuXUVu4Oi146KXTLTVsAqpWeEFxqhXUGJVh8U/QuW0mBjgX0HJovIqi24Gcmb
dUdOjBHM1aLRGsTIhnKGLclo5o5qZf3PZVKWx2Y31ARiAvO76Gnt4UORLwE/yhVIsw/3QeAK8ZC7
Z7TR1AiPxL5W3AbcPHeQVAeXVW+rA/FXhxp2uQ38JtAheE7nibVvoZjnaEvILeOXwbt1MXnIPC0p
SU3eUo3ZkYuPty9WE7xCXqmbjhNNco/kNAiAN3nINyeU9+uVdn9iO53Af7OCJgkxzwG5rsKXOiql
5Y/4h/k1bYw3utwP4wnhVplZ/nuyf7+Af5G0x23G/XxgQdGC13SxuDDEPeFzgG1Qv86otAcZWcrx
VC0Ngh+EoA44Cdj30GukyAGeDyYKjX1fwhpsdqtK/28PRARjMFcNUEQ+qq5ue4MfWQCd5CNYgLFS
4GaRjyJxpEU65KTy9/RmKJ5gbK1A6j2zkjcYbG7+Y5pNDJu0KWBoZzKQI9YpsQC9rNJtzmTvlWT7
/w+//1bn6GYf0srBFCc0sg8bEqvAAx+EZgMWmTLmE54vIrsGSJ6P8yDYYdpxJ8L5UFVfiFtwAP4w
MFOA3PHoOYAqZUF3n8+AZ8Hg1nQbqRiltg84/xPFn7EMCEtn48aJjjd86zDrlzlwLV5S8EkBLr2Q
A2NJlAh0+CJb+JuyqcUNXaiHHXl6wBWde4OG1KP0saikfR9i5ZdhwbnDUGw9cLmUZ20NwzT5QSf9
FM0u8AUUrrVG9FGLb9dUtGsBKjfWCPyHH9pw8f+uGbef+GdQM3pFD0GzqGY3EuVUuy2FZ3gOaLTG
BB1/XhEeAYEXBAiJeXDzoP66m99XbPSbG6oSe/olfDCTnKS0IpauujKKnqOKpDSjMj1R5W7dllwC
SoDmdftOCl6vHsifT5Eq+/s7d0vKdf/ZB3eUQE9Qi0GzVh+PZ6mY5cxyrPlZAWYI2SkFO/x6Qu2j
8+E17mZDy2zl7XrdfTnhdDUAkB4YuzXALxfHwrkGRNcIw6GgGBRjpwOC/WVr9FwH3MNkdIXjc3kf
T4omUBD8JXlhcq8cy+8+wqO6rCtMGTWrYGWlZY4Mjj9u6oYAFK5UqfEMhCumAK5ngY+gkjrLYOiY
DOxFOAll9SvZIajAymJa+IULR9WF6yt5YwNdzOFA4yG9FlbrUwvY5J8RvzRb0l4wMwFM455Z/fIj
Cr82gNEzPyqN2wGLf37XH1s7r/AkSYJ5RJfD5tgTgnoR7vY9ZdoASWlL7Ldphp0S0Wv8gj8WhiO+
bs6rzLPzYVrxOv7Esh+EBmJh3zPefa2vMgYwwtazlJmZB/YqaDgiGF+HX60L530dJ2GwEbEMfL+q
2n5yUcwpUoTMkv/gdEOLmyXRy3TJKq4FGwlTUez7XnzSjWVtaghymhbTO4JC7ceT4z1Wy1hyIwZx
jJ1RySA15U8FKoTLob63Ac9Cfs0b21Ilgu4uGtJoPXFn9ymtH8KV1FNDdpdW7U+AMHaQ3haLoo6A
dHh8Rnu44RfMk0nWNQqgp44/QzpE4HcItlMWeVH2zK3DIPnGgvGRBp8tMXD92lfP2ZR1XhzMqIWX
xStYPHsQFhpGbIKGsSi9I7Voe0vneHOHAAFo9xowoDu6+HX1TyNB5TDWJe+JmGBfgii+NOBS5+R8
U9hUkc2feRIpQ78VhIGQSHdT0UfkT0yZAW6clTwapA4srmdUfcUVRqMoo7mlo8GfVGaYLqL24TuF
uEsA+zKuUlOsDcJHMi3VERuDvFsY63Jwqj0lYapuc/E0ZGYGQEy7yGThN3qjf8znBSOpFf5E2Hh7
TnFBT4XRC1SVSfpuxrcNbGoZU944ZudFeqmStJwcbe5/HuASdI/MbhTcAxcJIgZX5UVrkKlpPG1W
LzK8Bl+LVIJ99webOVGnfULK8jT9iIo3EiIRQhlmRyyoYlC87fnGUXzRoOfyVD/CLhxJnl2n6WAd
Pl3swNnJiSK9I8vMoYLtTVLicNpqRWmAzOWZrsRabuNJCI12Rmnpv0VPFLdAS8iwEQDG/wKDCdr1
pNvlwbxQyM9eBocnfVoFDDGTHl5XFziw8wxWj9KEfcJSLNeJw6Skgc0qi3njgRZ1PHqi9RSpg5Ys
BxR7F8bhU25AOmQEBFE2FFNMMQ2kguNWVHHFGm8ad9lhR0LrIewfsjyOnOE80YGZcgfK/zCIG8xT
XQak0vcoxzNOewGOumfGJG2EgLnsSBNWDGFU4patKitv7Q8ZY+AI7az7IkyVTlV9QLULjYEvkcYu
PqamCSCTRotB8FKokXHwdmzywOFBUUTRqzEGajEG8vrupXGHZUF3CZt/S6sP1MI9VKrr4gG2fy1z
v9J2fRDSjEmDXpRgxw5W+BTS6XJJV3IyKl21ACPtfJOcSgp7FAJ8PwHwzLB2uhgHZSh0ziStu86F
sxixcgkAGllEC00E5zPrv3QTC+rfPrwbbuRM2uLMG8FEPDYWAd3AM8ySgExpyVqU0Af+QFTgxhpP
Lmnit8ONlZFCosvvb38gQKWrhM3syyvgGacnaYt4q/gkU+FTE7aTf0//aPF+KM+8qRk7rA9YUs3N
TX34tAIkL5BF19IiY55J3MyqDqRlL3EPjRQFPPoCEYXDpenSCZRPMI4fA4NMZZRCxH10bTbJyDb8
4Xh6ugFyNyPs3rPnzGfmF6MwFZqmm03ZgT8ArkEKJ5ZMKq5IFfxP//9G6qEHIzw6/OA5Hnhjjeku
S9NZs6Dk909rYG97zhWXx24mDqFm1dAyvNG1LKPz3Q3DBQbU6vpTN2uUzcMG7lEmBraA/3jNcbda
+XV7pzRM7jew5TZmpJomJkXzZlMajmUFh0cdXlF7bgvIBL8jG+A8IbneYXqGDHxD8cwO5z5tfNOl
Ubx8hayy1amsPp7N4Zq/GDz+xpwAROLmGXYKXjrUQ7J6hc2if6KvDHbIhRstaT5sqmdt663FJmeA
U0bawY5K96aNeUzoCyPlynkLEN7Ve7ctbQMIgxmkw0AjlR+51Fgc423jtUjvV4aTu/Mmta5p7ojW
XobOpOcRuLIS7pR/4K1UKXqADnSAJXZhYN8WinG0f2oTQJYV49Nr++1xEnRbJHTmikNpESVhcgBK
xFX9Qr78AGxnZs+zG1/zARDxSVd29QtDIbIOxVaYniV2eaCATiYzJLPBrK3z/eJWJzEJxx1AZJ3a
paLPdfnNJC7mUoiIxv3T+5qz86IYspMOgEKbbrtDKY/M9VZ6gdV8hlNt5oa3zfGaC/xBxIXuZm9u
ySbtgq9FDp6PzdHIdg10olFL0rHtZE2X8oodSnu5LEzZr6AaFd+G/qIiBzapkmb0yzn/ghJiESiW
jDNU6L2sGHmoSYOv/97jeJw/C+RdCtznGFDT7b5j2nt3rrh7VPm0z0m7xdgWfuE3sIE+UP3FZ/s/
qpiD1rtINxEmIbyD3pE8ivF5HrkKW2EXPQu593GFLeZPNUZvOVMHOfjsyXuXD9qlWsSkM2Gq/N23
j+wkuEEHh54fpc47QzYZnhYZOOUqvVb34Ecz+BLWoIn6EAtk/Q6sHIS73wT+ws21CvAI1jRgBBkl
y3mt8U/xIkWeHv04G+wGBEGwA50wCvSUN7w5uM0+VfdxN7JM0EPugXT1RUbQrwzfZmvH3mnGxfQ8
Oe49aZss+zPV8dod9SxIfTg2TltLZssxoRr62tlK6cSpc7MmiSclqOKan+kGW4h5nLkcHlICgvaE
dV1KX4G8zH3qdf08Y1XR3OhcEzlHfnm/wD6TQ8xcIVw4hqn2xRYA9ja+77V195TcJm713qiRVGMp
aLoSa+xldUalAT6Av4Uuuj/T78HLhK8vQTa4wD0erqhr2eY8a6OGZXDIi7JysnhP6Rv4sB4cxrPg
PVo1nHTtZbP+Ik7SSRXWz3qPvjHmbAQbTaGMw83bnfkylijlW4ujATR15vPxKVTohA+4jZOUU4vX
zIF9EWHBQBh/YH/uvU/OiUqzu6ssETGIAq/OVGklCjtS2p2opEIRAsEXdqZFqKt41Q08+AsTRWx3
TI1jkHvIPhgDdxmT7hv0kgwfjz+hv15sDfRqqY7+q64835hwBIhylVrHPgKXo/j0J9+6qOaUO/Sv
2Vqf1SvbLzhRfFCa0TN2wg7jJDwPveBCY5RCH7nz/FkP+Z0JIL0pxluKLJpuGrh1qNTh3ULM/EhI
P8wHXYtFsHFibJ3mgEYFy5CcFcSfW+tWxq6FadMRo/QNKpP+wPxs12Xwz32WhkMnHcvK4u7mboEu
gC+zBzcQJkUdiq221IhYhciYMZcn/onVtQ4gg/QtAOsyVRHqyhk+/V8IMCVEx0p+AsQcEMq3k0DY
GkVtBtndiurob7tnJ7DjmLDslJBRwOO/dqoE7mvG5LoCuH2UcVamE9RRTUGc0jEZZnhvtOuWdp2W
9gkR5ZwN0lQo7sRa77l6yNRviUb4UEMBCHZsUprGGwvSOrlB2uuPXvnLlTm8d1UTBNt9a8xOPqp9
SXZ5PMbptLngMl/o2a5hdOnV+SovzvKx82QyFnqJUw1l3EEFH+D0p/V5B6uAztBc62tjmNUJKuG2
wNdCoKKt/PxZXmmDc/JX7eJc7+ixQl2m5S8/N0ot+dGuTb4eueX5wOOQzru/a7WuuqdNK7MPNyZF
+Mu4oExK+OpNKLKDCgD587Et8OvY/NbReUrweXhC4bLpJcQ8TtCC+hygPXTOLhFG0NrLnH3InwBC
srUOfyqMqOHJL6m34mX39WQXlyGGUyXNYwb1bQBQffxsUbc2UUwbvcH/XqXh8yjMo5rzNyjP9Zvc
Ua3muV+bqvPW0Ccb5o2mN6ois3GW7lTa+Qw/wplSlra3R5juhHFsz+TLnxf6tD99CTgFvnxS4Tsu
1pe4cD2lZeHaQv/571B3fz2UQpFNgERAzwi9SnFVhrYWAsCzZ1Fgoper6YdJGdnnnq1An2mdHlNS
Z42WUbe4K8cdKnQFusqsx1b3/sNYEkJTRylkucnOPrCeW8jgMBdGZT/qcyQaVnO5Q3lCQHI/aGZ9
j7z7Z23k+zqOtKHekb6w/rPn/A0IPxNMys8w9FtF5t8HFpR6nAIirnKx3aLIWMDpOABiGPTVD5Ec
JqfzpV4echRB3zMve3kH4nfukwnVDcUeMbOC2UMF8n0J1tbPDkAc78RLpN1RgdAzTaUDoA0/fN+w
D4bNDsWyQnFIIT70u6diPyd7W1Qnyfbx3sGMY48LBygEQM/tE1KMZKlqgTkPabscvCmtSbRy1zsI
rzonks9UBchb90Z4VqVmRSimpHS1H79MghbTEdX/YGfDHD058yeC+J5ummV7TIpjqo/EE2WEke3W
ApHs+ggd2Z2FxkwOWBhNbMBafNsQKBkd+am3NnGNnuGGUnCcRuEz1jyGjXbpUDMAZ0BwEEm9Y1Eh
8zmWpVi/+qs57dClsDMsv43NgQtIQzZSZAx80I6HiVc3mkL8ntp88428o7+qjJZG5Ine5sFbVtVv
V0mBksxkZZvYzagGkF6X+6XpU1TQaMg1ThLQIzD4maJm5UU2ihrjvwmZVfaiy6xbfAgCdOnjn7YG
R2e1AwNFg21ikauuY9xNxd46af27b5RKM2R3CcMBAOeI1obaB33q7KYAHnomb9dYl59tDt0qJctA
RTSLNijzza1KdOj5jD3RqQpYz4QrCTVCeLXnOpHJtSdZQ/KUAMiKP+6HZmK4w8t65zkalXUR/THR
kwWuMsIH8rkcbyeCVS3seXFlo/Mxl6riBXPlqEuZvnY60lr5UZiwHdUAhUT9aAIQr6V2d4llaMa9
+QFKLPJGgbtIRnvPQq7SX+lAZvG2HFVo9lE/IjM75eQMoeMrdhKvsu6KKhNmE9ik6g9T8669moMY
kxIxJkr9N1i8HkiuCk3XfHWh5lOy3ijoY6AbJuL3MIzv+gI3HyWUns3/CE8gYsGIP2Eu9typCam8
Wr73CK/zvaANs+YZs6W/0d04zJq53n8hxdjjXd2JRT2357Pe8nAIab1+os1GJz6M2i5/xDOJikNL
XSc2+U2Cr0gV7tUWAqk5jxG4UOTBT+HEDAzZESwJNSnOQieGU531TDkWBGFjpQ2xwlqXkIEE3DbY
rktnM69lhoU8tznnEcMVjMi22d6mJNI0Jj3gjEPNkrmY4D6lPbDDVkr0ug5MFY2rkT2p2ovgLlym
K2sDmbEyURzz4WBo6vBF4ypVLXWC1QWGz6hZkacMEJsoom9OrSDh6Hdj+aqA4PmbiajHYNGtY6Bs
2zXmzIpqCkFoFSwiMfcZLzgWGnht8BT7iSEPaQQFYOun62OHwJ7oNOO83NB3k9TCKjuFaaHT7Lv1
z5Wwmn8/JewWOjJbiImuai97MdH4YMsRdSR+My7npntVbSuVGD+UF5TbbJzXbWzW5WVopVmW7JYQ
u0UlK5CLB0SYDpNmoXiVnILjWcputk1LeGgpqxH9/K5UhDNZKcIHGTN+v9KK73jAUXkp235rGB/N
8wyu9u08yUWdBYOioe6QDc0GZW787jvSpihRDK97mQGEtLAqFfKM/SoO4bBL4u3IL/zRXhTDnCBy
DUdHJ+/g+CSq4IAwDjUT5PXefrHJNQCLlJJdPQQF+sTgMEjh7WHrPf4qLF/JrtqwQY9syrDkFRqG
TxRhe4qAO0WMpMhlOZ+MgS/7yv7ktpcitMyTe2J6hmF1pCVWelQTz5leUvnI/Pz5icLRgbEb1Lbc
kqlaLNOrbnNUDtse7SmsqVRg/uKBCnbVXw1gdDsTIo5P5Tl2lvUtgwOeHBY8S6fcId1y3gWm3Dvz
bEUhT2dhG968Xdm1l6hTdA3rx27MCpJ7FhvzFIGovzrAlffcG0RIU+DAxZ372wqCMZ4suxQJsslL
xe0KlfTBA3gr5kDf7r3lXS/2myMZ8MyJ4XXsehzrq3t+F8uYt061I4kx44f2DKhABxJBAhBMsY/V
l7TDEiq1+QAAW6Cfj4RxP2UHvfcNYx34FVbVHT+/NMB/J3EkUG2ehcFr3N2hXwSYF0HgAeTER96X
RMPdjONw8rtav2qbFd//mlXglpZpTjfkwhGLJ++WeqwkFIrIun0to4v1YyKBpiTIeSleWWBOz7gC
o7u++jZfX9Ftre8TcfI835mHEwDJqaMeysDDRt6NRt+dtzoPoJ52C4szQg4qlEtVYFAmDRzywZqj
Htxp2vt8T8qrVcdUPhIIlo9F0WVmdP0ZUnUJCCdpsWrmABe1HIA/HxDFcEi5hKP8S9L4iyvITc6r
suB86OGzc/HUaDUsba7hYFYKvInwJbIMTAP/J9UuIqr1MlDzTRrSuRcajR9lAqgXyOeaR60OsefY
idhybRtxJHoyqM9PeQFdtDmkLtkvV3StNAUIBpYmvwUwV6Py8xXB+Pj//mHqBj0bo2hkP7Olrk0X
14ysYyw9iAD/R3y+qZ1v6onLAfwm57kfKpEzukpbwFoYfpHMvJp57IrcjbA75MQkZoqjNx4vRQSf
h8YRPaEwW3JWoVLPNhyTR1cjj3PHFjMxmbw4dh3wyMfteKgB8ZJ5cUbvafY3Y70x/aMsf/IhwTsZ
x3KW6MRAjYEFBCBY5FI/NcTQ0+6T8s1Pt1ouhtO3nrgBWZ46S7AjPWOIHyHRQ/dPFo6EMbfOF93O
TUtpiVOupwL3+J/yRMlMgqsHHWQ3RXRi4T2KgaNcW+2kH5rfOpXsThF3S5RriyKMcXVQa32RoQEP
13xabCA6Dz6c3i6rxekaS76ouIXubozW7qWzUrOBFMknR1knl5kYKYJL8Ihslf9P2NZvPbvTJVye
VGBfc2cXEu5ILCYnGD3m7uc6mFtMtPzxAtgYPtRElvjAX2OzQRa/LjaSaDOtyu8oRxG+shCMq6Ti
4/2nGtbRA4yGwhotJhB2ciWmRi7Co3gCqVMoD20l+05iEgKCveObvwU0AnL5UkbtQh3I5ko47qq2
N0ExHC6DsnGrjVrT2gGwJRSasPCt1njzhMidLJYIeAHVgIiMnV1KI8HsFAX3AG3Vhr9KVX4065Q7
4aaa3Lv0zJpcnyZZ7voxyI1V22J4F3bUYbpaMSLRvXdfP88spxD7Eo+k1YTHAEOl9aw2zhNH7zkZ
zJEw/ys/X/VTut6FdXsiCgCi92NiQCCghYCE9WgVq8D1ggl9VSg+/XQJi26Ao/qY8+cIq9ib+LEM
O1Lo7n0wWWoKBJ3JQuwJe07eF6zLUxgmQy8YktJCVcKRpL71hWzPaTssbyarpLKSmbBfYnbEMGwW
PmjYUzyalEN+yfixClF+MfwLS8YcTSAZt4OlgiMAz93O1u3VyF4NCTQkSaQZzxn29tzxqO6TQqrq
nAyFNUwuaFBJUyk6uyOoI1izkfWaqPiw5oocxzhmniOThRPH1az0B1YuibHHWBwmQmrEPQXYSsHW
gYjueyCJpQEPiQiAVDEjwzJHMmYf68QcCsWqCJe9UPWEmdevjEbstgtbqvg+fBgN/Ur9Q+76+N4k
ED5VB8zCLmc+82omk/rAdSpJZWr7QxlLbt/pR8cSsBriSDtN8XAiYSaqPzC/hVa/aokb2Xv40uD7
VEy+kuZgvqgG4yM41Gl0rqK4wP0GQ2b95EvCgBA26frzYOeKNCXHIWo8agecHEgivhkMYKAGm7Yb
kmTyPtOZkQOdb98r7iTrw0o+ocYO7p2B06E6xWYyGduUZuLj9g/bilw4ESlUTRyxzdNpfAOo6wf+
CCdLNAVhuuQqw1xQv1VTO+9HdIZhe/h5ojV9x/O+MGrHcXQIrKYr8S7H4UtvG9JhzsFpb5KPi1h7
8vTWWP33KNc+mOEcHRdfM/eqEvtt1//uSbA0TKcJaR4+EeBmrwiarN6ONkf4cXG5IZTVnTDbZRIN
8oH/wzKogqoB+hUyUOT8o1D+t697PMd/IXLvRXoaM+RjNFFLHngQq9Kj34fNKe2iUA5YNeZw06TK
VvI+gle2KVbpUsYSi6L4BKXrulYmn/mKk6nssW6stlgbJ2EKEmstI33B8QG2p8+uFxeiutgSScXT
ueA81OIfQEq2aIHbJmdJveZaU0GRakHohxDYeePgK4HRxZUY3m4oYe84KL95SRQKN2r9EASYVMAk
4CLokkPNqVq1uErZJvx1b7vx6IG51Wo/bGjibLy+ErGGiZ1/3WMjijltxeAZxQVJGp3Ov4ZCZE65
I0eQ4yKQhK2ozcz18JjXp/q3Mqv8mTsU46jC/V/bM3Sub/kD6yaC5kvJSIvD8byuJx0mgv9h198l
YPvm7SwClPJKdQlXS8Rekye6zhlxK7HoEx0J05p1rvFzVJ3iTw0MFle46A8mIzZm1qgsBHnQ6tUU
In6y+kaGnjN4JpsGSIdJZMwbU/ktW5Z6fJdvME1/7zeBUyDLKeAymay4hjdSw5528JQ2ALTjkX6p
eTYR+DsBQUfb7M6JM+SnJO4lIw5vpuhRQpmbmQyi4Cze61a38IuiD4Y4U7EgGaZyE2uzvRZO/Rdx
h5K6UnrMf+Jy2dWUO6panZQMhwNNsd2fc7rMlZlozEbj+xjPSwLeYwIKtfEcPGNV8qvvLD6+EfEY
vJDj/0wPzduauPFVAUr1zmck9lEInfbAmKGgPS7EpBDqAeC7GeCDXQLGimnhpjNXvrVDF9H+8+ji
TErhc0pX06QqUO7cvf2Yqpe6Vn4s6XBr7g5mnaR1xC8XkpRHi1TWEopO3GmnionOqB9FySoHpgA/
G5OKyUgez74/rnIn9G+66QM8K9FPDGd67+NlODPmNbwDeMOcyKdLd0iplnbEP3DNZCWDvJuo5PC8
Ew5ncCXDmBXHiNvjTkgxsI8+ITH6fCwLNvDZbR6kdpW6zkzX0Q2tKBM3wY93sdMtGxPcEsQzVxQC
dq0cej3Fe7vLisSmSPC3m2dRucDloUhx2F4IbDj1KFsLBYecqvPVrhVZQ5zSLRj2jVCO7K7OD7G/
34JqvxosvsK16lUZElJ/dzRcRmmYp3LhMAIKubI1S6Jd51GWpl2I1bT3b7iJFKR/psq0ALIvOxt9
6iiIDjUeKFb3a7Y892Kdlwk2j8ORwSheluWyO749pwoWsX/wB5/do2exW4qFEQcUigFdvX3VrYK7
NAlx/psqiszAmNMIaXCgr5qWWdU/bMwvcW85B7OQnYhx0DU6FP8HnhQc2zBH3w8o7dHgrMK6M9gl
gj8PK0Dud9yue0mVKd/2CeW4KG+4yN9NlGR4c5KUotA7Y0Mk7DcjZ9kIzIItJJ/6cabelZ2HT2GS
SolnwdrkXAc0H3pbMvZegYJaE2Et3EPrLmVAaKgJzbajRs1yxd998e2olAGVbaIOjM8BHeRFUJDN
oaUyKjLxCeRuIABH5F6dtGTMaVJ1oCiRzXPEiznP4lPtpx5tZIcnaGwk6/S2p888+QVwVTkQLPfN
lXWWarLFrPwyF3FeiNg3kwHs9EYMEblQvaKqwZSYKC/pPYzU613VZr42a477D+aI7sYhhazHMfH7
GLlhkvmYNgx09yz+WaObTv0Yj7JI/2VBxK/osXrk4hA8EOotKFT4mQOPGZcpro4EJAA8XeU/PCHY
hjtk+TAQd4VKRXfApv9YAV1FxBV85hJEzLI34ArvhPe/pj1/XWyytVIi3VPa8DOY6hD4gArcoEdo
1M7dPxWIAX9wLEajTyeQRPqG0KHGfPbWU60Ltt6d0hukdZ4sqHuAOYx+er8v8zOgBxpTW9jecHAd
bdOwUcNQ8CauCsjD7sBxzL6nvNgi+JR/ByZhK/lxg++CM8DQ5qvpDorCqeEvmFZgD9AbE+eo4BVB
6m1ycaJfpnUrQ1C1HjDblMW7y9mQcXS3oVDmAJxTFjzRdpZyvJKyycaYj0Xb6lUj5p8guO59Il4p
IJ0wurGXsKmIxY55duuATZ+1OLkENvIfd2KVVD6c9wJSfAPlaQ41H00BjF7NBhAY0QpVqOQRiDlP
ENttbWuMDQx+oHJFKvvvaA5qTXGLjDBgNVOTPDOSyBesKz/QCZWTPm47WRYk2o2hRAKskzyqIX8N
UDQeOxQ8ViOW5vvOZevyQq0FSWqlCb/jat3LYVoxKvTnQaTNq7qIQXPs1j4hXc/FxHOk6ZJ+VIWO
DY3jIZotW3U5SK2lIZGXQm9MxsmkslYafaPfSt9UUrI31XiB7kqGWEWUOHkevS8yM8eJGFYkWDoE
Y/GTfNXUtoXa3Hcbyv8MXL+tY5gDShdpkG0QJnWRl435w7oiny+pY5wif32PsiQK1WFg+UhOcdyT
tSO/bzOO0MiVixSfdHceyV2N8/q8WWyoqJIqhamb0HEurTt9qDt7vdi3iLAFIq7XzZhP2YQrNEWp
cQSpcQQNxtsnci/BC0qWAIWvtdXHrWSW167A4w9g78teyBFGzsj5V3BTr/OiWVVCX5b9L7zAd+en
X6r182aD2LUcDENuM40Q7Db+jusay05V8yfyHax2fuQs44D5JBaRQ0XTkScBnlomD5cdeqshmHaW
j92H5Wpu05BbeF6XEfv84kp3GKu2PrJujwaDwcOvhF9Qho4BeBl8nc7PZN0p5nF5mBh9z6VV06lt
HrRHDV3lzXkooESRAY60GsrA+xUy72276I/vPxMgm3r9ayR07WJkgI5ZiUFTSCDItZNN9VKLlHN4
xo/YIJfXC/B61cBhB0Y4Tp0tezEHYlMMNJ1psfLqlp+9B/zUTQQYg39QsGgydCyaXEBEMwF40V/C
O0XdIyPmVfCKrOXaaDsq67pEzfT1s5yJl/igKYPQIUDH+IdOLKHFdXuHzR6oANNZmHptX52I/Psr
rbfbwHAVzX+I6dDfN9+cHy39nVKbvR1Udzlcgn+ThywrNfPJdVpKISFQ1ZFP/W3VMrocIwHGryo4
OrjXH34r7TXfwrb7ZsnCOnJFXqXJk+WLXhaEeYdUpW9zitYosPTG5UOqjucw+k+0sDwOXyDoiVgh
L9PwyPURF1/nlflW1B+SAAb8fUHnhnZJ4EROrknCRI7yk7bP2qsJ6q60qmFvA8CMCwa0kCNKdhrm
M1eKvjJxGdLmu8wDQ7+Mqg0Ro44HHGFk1D2R77NXWIWURjv81Iw7Nvi+a2jJn6OPgR5MrASOa/LU
cCXLrpd9qEglSDJVgrESkhVJabdtKUYHA1/NLW6eUyXM8ia3cLZpYt+VMYWzf1VhlbdOkkXPLL+F
DhW1mjCFt3PhdjxnGwwpM2d2PFgy+CtM53jSd0tHZBPqN2o+tGDIMbLomW+oMfFM7BaYbY++MVsa
1xDJKjHNUte5A1NmK31sTVo1NGBYHnAPfjLAmz5lqVoGiKdGqzTtN0HtnmVzLL/fDoIcEBupRlc9
5cV4+EtiZgWr5NwXn8jkvm6YIgP7F4eeyEvg5FQyB0pXPtt1bQo+itQpU+fUX3wNyF9il+cMtV29
bkbK+K0Zmdkwo72fK85QWZ5bIapnTm/E95Js/aH2pQZ/EkcVVS3pqnZviIeEqf1NIwUn0y/WZar9
Y5ZF7/oq0zto8Gie3Ijgtfsx0QhiApAtMr+FslSABWQey6isUFZRqXmnnXeb9JUv3iYsKUtF2UzG
NOi6ATUjYJXNWOJFZBcPKMyKh0sEirN0X10FJWrIUImQ4LhMZUTX9IlASVedDxpeMt3Rqqoc8h3R
cf1Sor9D+MkkZVOCu1WmQpHMwnaeDrgmEWf5+u1a6w2eUaAHxlSV8wiVcRNQ3iaD8IaEABYxSreZ
4T8wt0NebQZah8TY1ifWa2BdCO8J0n8BN58PhT6/HwiFPv8dzky8a7GvlhuqoyrYyZPaHYKl5WnY
KAVr1HCNA3au6EoywCoq589eZftE5SUS+KIUQIWS03CrtKjGkIGbBHFw1xQ6ul8deGmDlwzH+toK
jD7o8ym9UzNvPbDIiawKd9KRUSREETm4Cu0uitOSZ3i2h3QOGfHSwSGQ6sUn0AmMLBoM1dHB38c3
0SEwtBXDJu8pr07eVl+ASErowKIBVV4LFpwd1SawmIivVinNB4w1peQ/8KDW7uIIsFobpPlJyxfm
W40ZiZ4+qNY5OkLleVUcKawqX26eYcdUYfEFhjPoXnNLaKMn+DqU8DKfIe5uk1KqNQiWkO4d90dj
/ZuJ8iOHLhqaIDgazcZBWEy72eRea3rFjRVjjwdIU0hE8cD81ppNP/d7wI8ARJz39hjChrrkymuQ
2/37DGL61J5iv7RJOMXBioWpo1XLF8LGzqW2CdNFvDXz0UFd3+m0kte4lGUWaFoBHDXuUNIsVMKe
62K2J0ywcBUHHY1nvQActUHlSDrPpX4bcc5ybImtwM96dxWa1L4Dbg3BZlgVykLzIKyQJHHBDvm/
J99PUJit/k6SC3673eBAFSvHdWRJAfhPjUBZzkGCOMrZxuMqw8jwCLSGn1pNzCBOQaseBUntR4oS
5IvOI9z0wF9XJVUI/qBHsCTyV3p+p+VX6h5M1GEBaaPT+YYVoYTwk5zBnzY8GorJqlwfwhdgPCft
ObwjZQhXuECPx6e/CbtwJq2hc5tiqcVKOdndQ724EKSNx3jC1An80ItD2yKe5M2i9jCL5ZtZjVZK
0zYzsmOHEHMZwEiJkvfD19H39pUqIvito8kKi8+i7njk8budS2YZVBRYWvDcamLxnmMmlx0GbKla
k9EZfO/BnxYJphp/bWtT7BKg9njwVwCOQXpxar4wWni/5iT/XHVJdaXZ8SNCkrLgbn9tUhnNkecO
ge3vA6A8Gcv5KvrZWj6pxhg2H7lbvZjywVZHOSGroPTdw7kqaxL0cy614qY36vhz5v2KS+nyicXi
SzYnoolnvEDefCRzuzgOA7oBnqeweLNxdokNV1KMiIKMJVdU4bHTGnzR27WRJzCe0Fxb5lfQaDyh
d6oxxZCBX7nPuX0hScj2Nt8rt2YlWdZNXew8Yx8ONPlzbqCu5Txlx6FuaNCx1MKtcutEhk24/41j
38rQ76bVaR3vxYRT6ZuohzILCKvCoAfdG1K7M4S8gMO6LV2MVl/xXDCaJ/5r8i3TY566S3ZKnJpg
9X8811ypikjA8cQSxmnJ5J7aexxNRPcHddOxh8oykAPlg/Z/pRnJNY3WTdQvaK74ereXLjMZpWi9
cYVbgxu2nMFsUP1DBO1HudnCun7QHVsgAlvmgegYELLQK27njOUINXfk4FtbSHgynN19fIYALuwk
Rj7XVgp1t6fPpNtYYrxjWfyMRgLcejNGJMGEHC6RGrutZdrovcT2DPX4J2yXmyoQ/LeeO8VNiZXR
UWnawKBtPikMPK5w7iZwqaKroCbOMIz9QpfXUIuz+6XbnpeB9WijtxXO4gQtWI6u3u1sNxLXGBUk
kX1VTDKNz5ihj3mQ4UL0jQRr9xohnl18BuiCPzA6uwv2kbTrPUSg7JDooK1lacmZRfcqvcznXEva
SthrwVssbadYPb2cPAP1omctULSmf6BNaxxmqD+ZvQNSctd35SD+PgzQb7U5kbSQqUhJcMI9lF37
ff6sMhL1paTAcrrXc6aeJUYcv/dpnAlDxByMZK9nkWj751ev1UeErx9EmTl4Zs2orHNeYIXzlZNG
JpHdi3UacF+gU1+CtkJ9B8jB88RoisikGfwRJV/vP6rQ5mFxwu66PD2O4WRx+lskye0UxV93URcq
gJvdgWJ7Bje6kADVBWUkX4eNlf2/pJFOvctush5ITYKJd/nIgdXtaOhyKJ2MeSy2N/k2NZ3gmMAk
55Bh7zi9/ode/AMooYCuFQQ5w1e6cFyXGD3i7rc5UoiVkZzSzu++cf3h6WoHE8SpeBxFJPYdpKdG
GW3qXP6ZKXvV1kpT/j9JLPzRzoRk6+ArEIFK06TejiHRvkk+58Pcwr4SWxy9MqlQ8glZ3oECzKzZ
tCIBowjNG0nbmp/tQNZ1dj0lOOgIzfbPQROWBRgsB7XnJ2SxyTjRhghPyVwjiLxQT53lpOA6098j
/hiG1KB9bsjsNtMJ/Ulg1gbW1K+ahnTEZUmYc5a2ITQsRd2LfiODD8zeUl7fetgdcvvq7d+xNOti
PcIxU5XFlUxklkArY71bDDciS5hst5ux+VSYBLL/nBz3VbRWqJcqJpNFIeo/30DuLYRA0X1gKs9z
55sSWWl4QGQuwT7q5E3r9wO/yhBsTG9Swt2S+Z7t5xrDVjL6sdaln0UjlGEhO+A+7bEkTOYc5UR+
b/TKm9FY2joUrS1xHEXfU4sZaP7/N0FANuzEDnIFwRiOHCMOD/KsaWjr9SDZZXjKXja6dl4qZLdg
SsyZ0sOqfocUDuO6NnYpU367JVOePlROISwM4pm3DAnfo86lPZNrwkFFhXKVGIZU0kv1PHQbW6f2
5jUU1oJJ0JhNEHVBfjOCpQujW73iGur8li8xphT8VjBaaRA5ILK1bGFJ6n7+M/utIPCPtXFlW3ZW
bkK2lycYMVPFgmNfQL/klRz8XlSEuucNFzCmvF2aCoXc18P1VYt6lbg6FlAC3IFcxhFWVU6LkNjF
q+ujEnbAKgv0HAoh1aMXy2v8G7HUPKlhnZviTEq+cqg1/Ffv2d+qTYJgjE+75l7GZgFF/P+VP9Fx
2YtWt4dRe0RhHHmYnBD2ynvxLUNX+23JlP93XAxI+WE2aAlT917Ism6WerO7FqqnPGJ8UWiZvY1g
K3JfJYz9u8hbH9C1jgmba+zxn7bS+RT+lRRmssZiTlw+Fn0JTYIOaJGNdO0Lm0LZvX2zweUVH+u5
jOnIzFMmY5dU7+820fMDvhc4VWf4aAiXhiIDn/cge2EYmu70HPc+h8UvOSQvwMpofGynyMOGH/Gc
72pVfXujQZITrcTYdAiAXcrZcm+fRiNppdQhx+256whGnz1LAvtJ+A94HKhcPiexBfff9RVU5zU6
NmrrsBsWETJ+n8x5agIga0CJ64PNfNnfYEd8kTYSpBhoEq5mIqVzxDj35zuBKns7NzirQnwMDy6t
bQI+LxSllJWYuHPfkx5FZiCh8WnRTA8CLyROecE4lT6JYE/ICaGeQnkLmCLU/9/Wbu93wsf2nto/
oJVeKwEvnhcqW0bmSp3I+r4ZlEqJCI3X3Zc/yBmvsskKwnrUbUpgn25uMzYbhJzZOEZVFzL/e4SQ
x8YaMNdw0FGyZ/JJY39/JI2s1LD2Tg9iaPd9arw9bKa2gWGBJTaNyvP6iCCK6NGADV93snZdfmzJ
FEs6Su45S47zC85lKLozQmMWrWIKmaeOM3Eugx5c5YFTzv4jxSTQJ1T8MavqpNCVA21Lr6WL+Agg
2kVT8GSEqh9Paf/SvFTTbRRi19AXSCt+Ts5CNbdK582WCbS0h0/g+XlC60+G3s0+L7XJkjX5dMxK
FRwaqNNy9PB5qPVs6qO7/PLYkoaU3NGXhBNENKXF3pkSjuzg5/t3sdgRpveBFumrVvk3AjKLRXxj
DpGPeFHdgj39u8Cts1MGy3H0lPbFWM2ebDwUg88v5CyYCsEuC/V+5bpbZMA5WDWfOCrPSUN1P42Z
kV8hGQO+2CPZxlkZc/3syi4hVdyHNXIxt4e+kf8iqxTdUeVhisr1yZStQFVIU7FWX+CkRNKUBRJO
dTFKK4H4aFgp1JRUGECO2aaw55vrCemOYuv1W2px8+l3wN+RMBuX4tiJviOxiqViO3ItssR23RZx
op6u80ojdyPjEr2tuFGf2cYKzuAMDQy81AItoMxvA9ljpyfRDyM827qljcKvZTQeOcXFK9jle/1k
yvsYpLNrLfflxzi7cxouqxwYYbuXhq5GryVvCRv/EK6iKewdKVIq+vAq/FPStqCWlTYRBWlymKeK
XKWxBbRhsbBl/qQPTMJgZz9BXUNYp2OtyKJ9qi43oNLu3mhbZIf1iHEv8iqsq9R5c2hxUgDqYtLx
NR/laZwCW7KJYDsWed2eJQBC5TBWyvkPVZQlcvCq5aVskTuoKkMO0OZT3B7sD5vTMPCmF2fuzTsi
ikKo9aToVr9AaQCF0dE0KlFtB1FryjbnYer8YVqSZ9Vg6MiA2GUO6+RXkJpJN96Y83IHOUXvI1Tr
cVUz6DIUeEuhB4olhwZvTqWkbkbuFnZfMXTL7pVKGZLyoM8xJvYJv4DVGbtnCRDjlibbgFrQraho
pk2ijKOSVHCZbHKGWZw6yVpODXznDt+SDkY8+OmS2S5SYhRr1C8wsArU4Kd0fP7ysUH5O98mqvpG
yCieWk3SQE00d6JirXcdL7yxkTNwueRS8h/bw9G2w30zdwlH9rH8yytlr5q5WUGwMu40DOW05I9r
IluG10mhH46RSS3bailfPSDrqJZuayTsuHEB/EWsn9rSYGQ+K8eliakmkDe8aCFQCCcIF0dnS2Hj
Tn79rxKpqqwn/xOBZVIKs6ujiATuqOj7frRcP4HpoF3O8yYq480bt6qzfgzzDrD+ddO8H4TbWTI7
YOL//MPsywTl9agKH03u8T30IqPFWL1G3IQT4jn9yYtvbWpRVXl13dbUhVvXZE/S1hUBJ/kg5XAC
cNCNJrjBL0uU16d6y3T5PCpfvVvPrjXIdOGqltnfMFcv8Fp0gISUm3dX5EfYp9I3vCWPJFVmbnRC
X6AoECO6q9iRBfEulGPYJE2/vOgk8dkE5oq1JofBkxAqWvVdKwa0Fn6a0EyETGsIPcF/XhdIvLc9
ph5Rz9k7KT3/o+i9Dy2CuuWQT/Il3yt/e/7/oGgFKktpQEl5CG0VRMMsFNO2Xt+j3ec8x9LEGF/0
PA3E5Pkp32eYGaVH2U8OlgM6ztjQEOukjdornlq20y/OJQdnwnQnUhkxAEJkn5Q///HORuwJWMMl
XhHpyDmNUORglZsT3y8+BN7bbZLav0K/L8m4cUNHh8x6sKCV2CyYwnzwjOrOJD9oZZVmb6SdwTCj
+/RoSMMxcf+CHB7+3BofnGjGbx/cWir+Ltv5QRQHJSFEVk46v0T08skKzAzg/bD6menLB/H3i9/m
63QT/tD0EGOvJbZhV9H00IuQedfjS8ree55+c6UxhDO6pKw/pleSUROJxQ2qtt/bBMr/QTgWw7Ud
qbBB/HdAIwBp/cBKGncOVfJLZi40VUhdD6SUX/F3Vablue5KY+A51uJxEduXqkeV2yFznIocw9Oc
nng/nbZgVknnl0S/uGc+/2H/Z9D1PdhOmw2RmV5SMlkyWkIYOEGbahxKSo4lAKhEsI0Fef88u9sX
7IIJM+nTNhzMiZP60tzTM+jZaKyNM1GqPDwcU8PzBOrHrCjak4v0TmC5Yqsa3RLWeGvw2U3/T8j4
RQHHpAix6v631zGK1vjIg7ZHM4XaMdIsstshZl0QuR75lOa4SIquMAfvvfBneGanyPqbkdu/CzKv
5GjRc7NQtlM/rUpt1FfaZsteylpI9HRZeTlZ5o/kuyQm5ibZl1zVbHLGTI+qJDe4/BCXkr/DFU/I
5c+ISaA5NGzcbA1p+Kkv3wFkdiHGpnj82fRiDGzZn7uw8AbmKrqH0pBP7hkPJNYYZ8dLhk61FSJj
8nSPECIBF8HysAKwLKfZmGfqhkli+EEj+KJNweVu8JOYqwNlQMOPnQAascOf3u4xVk3/r3f3jNyh
5xJ29zUQxvvOwOua35ZKKUAJuhJVQOlH9iMySozdVuWMXGJO1yrr2IaFTZXcCq+TXkzXMg7A86yA
ZLLFxm37pH+ATxsrMy7fgLuYx5sa9bFHqqlbxBnANBC9SFWpknOiIPAFWAQ0NzkmZZkAnxGJlelA
1QkwLUrfCksp/6lTsOZ1UuQrDYllZBvPBbRrl0sYGGjAg4QnnYA4iE5elDSSKdBWyKGNaZ6tsDDQ
c7SbLbrfm6lF8NjYIv0vre95vR8OIxV6G3iil2v+8soEW8R5asVUGpTttXYV1ofxxKQCN/3r/0mv
gtOZRNim0JwIY79K09P0ffz22ioYNRUCbmtwq5pFChAnqoZE2KVvBOZUSpO0T2F/owj29MvCuHru
+BwypfWc2R4IzEvCcG38JkawD21MZXPhCi+qURT1o8iis9j7QgN1xKDp279F4Gw8t87WRe5ssF4S
3sKIBC1jux5aMT/cmXg6J8yn2gRbzjTMEZRAHGK3RYZE0v0A+u3WhUgSz4uMm76cq4KD0uyIdk5Y
OMrv0DcGCgp5JmUbwlob7NjRSx16XwF8Xp04YOsbQKVUDiA+TyaKqfUVvAknVrOJ5j+GbMoXd0hJ
AodTE+63J9f6o2M52LU4V3EqsK89rAHseEUG9eGZ39toKn+X2CwuqXa9n0OOPCxYAJN9JwwWtYF6
RBh5dzuYBIPIcosBfemvhnVPHZu80amSf6AtptqCRiiCGEQOZDXifRQxieY6+0j0LWPWJgeItDjs
An5kdNrdX3mICN1uZWE1VatTCgj52bTg9ZUuYInfsmgWSZ8rYjyAVdZXzehodwCyrUwQvyJ21UUw
PBfYjAYXyl5q0Se95H7knMUYnVpnHYsrsEuovpv2fhJd1pJJ7pyf295VCxUPWlLc9ydE0kEXe9G0
RHEgGSsyql+pOl/4dhme4X5J+GFCPJZOQMg9lcmklUxIUbW/6MwqFRDzIt19ECGVbqu9uYSxXcOJ
BMtQbR9xaGGnlT0OrH1NBo9FYwfSCp35/79DtLSU8glrcTQnb+6ueIQ2hOAV671CqSynBYeI4q+8
qQ6N4trFVQZJD3GZMQ0nggYTwWZu5AfO97yZB4T0JjL60GJk+H9obXDXzkM3son+4o3CuW9c79Wy
u8Ve+BadO2uuEh7Pq1bhX3zxkw8g6nrQXMKsb/mCj+WH6jf7EMov7PlzUBfan3+Jsl9HlOPHgS8y
UpyRyu3HRuUg9ucCxXLxIZwQTBqkbWJBNh1oH2Ogwxujb/+HLiXbYGVR/hWBMVKcBt4r4EfVrMCl
FZbt6aMWt3cUKQG0O4uOHMBXosKgG3MC3nkF6WAoQFCTteruC7PnwaCOaVCRv4W4wHlNn8W8Ce3c
ZIxrVWRTP4xqZiQb3roINlDx2hYPZueZ5uQgnoDptSFeG/LIB9W/2tWQzHikbqhFho4tuxj3orSi
tbQ2aSvaDKRT2zpvHPYY9xfQ5dVTMy2FIJrnxpcAOC8CTV8o7nfkE8fHY/15niCkN+w93/483vfC
7/ji1tdLtq1MQfanHtaOk/w4yfrlVV4SKHy/2vL66fvC5vpmVTahOlh5HaP6Lcm3rWtH9QmpIq7q
4CKt4YboGuYgFaPY9HuK1I3SRYjcFLgdErucDgYCwRrxPIhpl+f+VLyWEwQr1bOZwQTWAHrA3eG7
74LkDTDkPGiOBywD2QaJ+K/RtKhVxMVYajaO3P+IuotIAl4rFGL9AhlontwJbqRbh8rFERq+7BoV
8uElUztZhSpbg70h+XKPXHEnvq3DEA4ObZHMoVPpuFuycGN09hoewWgejg4otjV91Tlvv30qguek
MTzBodEVcuRpPalRbbmT07iPnSBF5IGwPMN5E9JpD4LiAuM0FvBTTdLK2liJNLYYSZ3ZHsOlCQUX
XDWDoNQz4DDDTamwnBIr1oa31oZ+JtMwX3nzuUMpHvRHqPn9RmfcnHO3lwh1oDD90iI+urCVqRY3
zIPqP19WwWYIoCGAX2D2z1/UbG9v8CW1voVL3nKYsoxkVNEyfiC8qUgbOuDAJGzS77r2+eann5nz
oelG5jcvyDlYJ4EnQhxS//h4Kw5B0PVBA0XuhS021LXg9MYeM1l9gJFX2rcHhfJOLUflf4RTJFzd
9r9ZOBMvTHVe7WyqNPTKizEANKlVQfqipa5LbFPrC/9jBrwnEoBuRlMkeJLYfakG4V/SatdlLfLH
wOq1n1DkfBCSC/O3hO+9Vgz87cedyDRX8ipmKarxhBT/D1mb9Mk0u3nicgpum33YMOY3UvwW4Oag
B9daaf0dpSQgKnEXjCIyPAogCByQ/qsmHaJ9dsPUAGtvqS2SDFSbk3hP1iAU8qBgTxh1849Bhnxx
q/hdHZV/p07PXpDptmb/lIBHZ0rVQccv31qv8tZcvfQE1ZK8SjteNzRgXxSuY6jpmpoPD7xIhHYi
vdmQHzgvQN9YRfAhr09bhi56u6MAyWSEpcR8cjDGtCnbCKV+Q2ubzFlBeD+pxvdY/wvc30Gic2ue
iWFTF/j6rmGpFTzpnrAoP/a/A6vTjieLkFctXmS1raZ2rr8ViDRC1DdrTFdRpAz6SLY/AVxh9yl8
XVUoyls8hEOfSDP5GoUfLNA0yR/6usbnE/+LJCS67s9/Lv8Qh2JKl8md+BD7FE3Ep+y6SOmaSBO6
i8kSMmpO4GvCPzecW/KGZydmmOdhLvSlyzWrFsqM6yIsNDOI4Gi9khsEUcSZVdf0HtB8DxEyPsH/
ckd1DyBc8HMHE0CH05Rip9MwbZUMbTXMXuWmOVFyUbAI1akZzmIuC4sGDhXIZrfblbHTQ1yUzCHY
ovmMXWC9dGMbQ5u6FeakXBdzzwwRuruQQu4Y+HfI2LkiszrMGGRNVQ+fC4ZpXVpqdGL2hCUlf3vM
eVU7cCjrFIwigsnn1YJ1ePmzk9wddhhAmP7m2vtcSAzq0AdEXqiwfB9oc7iwbFarrqJkUInpfzB/
qXSzXPcTolN6qhM4H4BCKuRsGVrg9I91cAnaXKS0zzQ1PwNjUcpNHuyQouCgWbtv9oCfA33yXFHe
YNluG3zJmRuHcsj2Fg8M3UnL5qmNok4N5r/b4TJJPTXT94bHi1HxXgLi0PndM2Jbi8KwAk2Hw5KW
BjhLxRguH4CQ8M4CVNrK647KKWevpBh0MpNknXcHTEqfUnG1qvWU6oeIRM7RxVsviH/AqESiHSh6
8PTKQASh2OIZ79OJlbxtVivK3/sLBCqJnV3ddhcZxhr0bm5hdo0Ya9h1XE9TJwRYMCcih6n2ik1f
/8Gb1wDpCzxkwI52M/g1VPTki8ERNeFz+3TUg9QBUkY8WYyEiQJQ2lm1IDjJPkHIbPHE7Rc8K0bY
MTv54blIJ2Tvrqizmb46FgmAbNcRVOa4cvchFh5dTeudGmSI5smMguuqWoqAfla7ND4cDoaqYbJX
3fj+d4rbTqAdABWt0bLXzhuHgtA8okdDMTZGAVQbIYZn2lN7DxuOKwYQjsjJCX2dudPdelEr5Npo
CbYMbRjDoiO/q5ruZwG6pNuaRhvjnFwm9X4bMyqpSQRK7hZyjYYqnbcB/tOKmAl1ykFXQ7c/KbxM
ZOwKOw6xe+uoS2KtsUHnRayX7bEsZKmUge7k7+jWtc06+f9Zhrad1PBNq+FizFelUBXCS5ASIN48
FNMGxGwt3+5F4ko0N3hotU68sfuD3Ss6DIOoFjKD8ZmNWHvPY1XOx+eFPISXKAH5AdAT0DsAiuga
OFLYbSIsChtxlRGHo0xNBnNRsX4HKfH6At7RMxz7T7xlozzJbFRyoydO+vkPhc6EJCz8rxdrOpMa
cZ6H/tg5pkuzMbOLokjWaxhOTjJ3+SXTJz88wJoDNEPKKri68X5Gt28tzvVqSC+kY2vYYOrBFVtK
l4wqvYVew4SQb2QCNEMB7Od+XDKh4hb2P61Q6sYmnCAT+N2iUTD3Km8Od+D0+fDcTjjy8RMd+l0f
+GU6rmHnGBEZrYExqcb9HeZS7M2DCXSt6xK0VkzOzj01aiXtPV00PlQ4Khpa92M+qLtP1Hlvcfgp
6oDEzJsIlbHwOgBXfoIofsYNvlQrxeh8wQAI88JPkmJSDQlOnOc+FPmgjNRk/4UGAYB7ssrlsI8k
G1H77rFRhFGR2yFyXF0iLKA+3m0UohCgdW4ozdtr6/SLlzr+whFlfBiwZqWhQew+8k1ojSBonpOw
C4JnRaZ1ZlubDpooBZtegjjMTvwZ7nL8sM/FvffFW8FV6tZVbkRIyZLk7y9AdnrYcKXNYaFWlOZt
9FglOyxJjazUmO8t4Ik9r/Y8KkiBqXncyrNKBE2yie6V5OcZ46ddXp4Hgx8SmiVGSsJlsur46a0c
ubUi+zW1c7JyZt3z5AtG1uZmS6ucfWXsPHklhSBo7mHMVH86F+k/KyRB3kxXNsBHlkjEfbKG3ieN
0WlWg4OrsGMsY6wg87mFM6jlIbZtv58Peyo6StNbm/tvVweJCLiEXOd+AKc5EIyiM+MjpPjg7pHI
/IvekIB5ren++R/iJZwrP/Za9ThmMgSB7ngxmK3sagQIzeWZYqp5q5IV6dLDEGV6stTNNhhm+MnR
QZ4e00JjZvNZuDuJXKZFf2ynuVK1mtT/jAABo5vDfnK9yIeqmlzUafok/lGuJ9VAWcXgPvBRrlVy
pxFseanZBso7cCsTlPmw65pyjsL+nkanUIzjj5ye00WPEB6Y7kVIPQ2dGWDeduPQFdVYCuq1RMct
1Vd6rHmdu+yiDnS+sftPvv2AMpDYHfYOjamDG6YqtgY4ooFx3zxPtlD5MZnXQazgi1+eLA6DjMzI
D+nC1vcYyQ3fKj4iphfLXLj5Y5UAzWghLMcIAsF0hwP4nenLuDcTlzg0MpcDGNO0gSwsa4+6XG6J
Eooqos5bsomlovHGApLXOUWefzIKWEI3/mxDuw7tLLAfJFfRNTQ+yGqL8MbTUtn5RY7fdvDfSG9H
UI83AC4RztvTYFrlGABo7QunwWXeZ+gl/w/JWoiUG+xepCRxVGcE+mqhauwi+GEBEBMlR8lWcWIj
nZqoHea8X08UWsqNIGOaFNY+HxXBYxbN+JIekG8olEt2uIg+xcb7pReWTZGarwl090qEYjG0vuSB
RflL69qQ8F2SH88/Q9r6EFm8PHZCUUlLLodJOoKvxNrgID+zY1t/+ZrVY2pAqUGkRiinkTgztFsm
ooU74w8pxWDEmkaUthugoKngA55SodXU1GVYGcMfaXucPXiDY7jkKBksIYSE6rcQ58Lx/2cEL2X4
cydiWBRNgS5KXI+8hBQ4d5ixFHfKC/bUy486HceYEaSfI2ZuRO2tvkxwGiOuMEGTnfOeWy0MBO0+
nseDxhbU74llaCEtpXdfSbLp3jAo6d5uaQXHhOcO2SW5qRe9NITTxARValkO062vzHNzSrqbJMoq
SUMfP38uLEZddb4O22CFYtRgXWhwMP475JOo3K8EbsKro127OvNR08XfNvS4pEOKwy/dowx9TCAB
TCAjMJlm0WSLIF4QmpyLbVtiOLi3eW8WTrLHmQF4uApQs5XBDielAlVoWfVGNrxrwDlk9VYPM/me
vLkSMUpGUkgT1//qwAr6VtslXp3GKnpFIQLAv8ICYq8CA+Cys5p65vLrM+4QTiUkuK+00qOjRvQa
jcKUmByNCJfok/uMKK1Yh6N5ZR8qTyLqxRUQV/inZSKTiR36bjxw/rW6dXL8FlKxEoO9rjU3aWV7
sEmBa8NUyctxcHFpBqF/+dYx7ZpchupBj0z/e9Vs5NoYOI9Tmki98bl3TP1eVCgxBa44WCPv8H1m
CgGHEJ3q9gIrPZnx+EZ+Nd56OdwraWRufuvuImW7HBPA1Tb6dVKj4myqHd65O/r0IrjXWAN76PmP
TfotQL4bfc8DmjUbZDpW07IxC7PbBhMrG18rJroQTu7jEzZSt3u2hgENg+Mg1rWoD+pKnlfQ66jy
GRmKrw1B2l3Q/55snG5EEzBypGam1J4rrvWEMhCc2Rx6dvbVTswfzGLYBHxy3k1uQGcsemiDxgmm
Rdp6m3VC9VUmz07jza7VwG7z6H+Zy9/BCYtowIvk23cNoQBSjWHCYUNJYp8SPd3lKfb7r+TbQ96m
QwS9F1HlerZxxyfJlBiZ3tb6Fs4Rku0yke/fH78hIhAk/j6MuW0ndgUNur/xRUelgKJas1qASARF
dNz+4vVujidGBivCE9GSi7iJRca8HpsMahS58zYIMWeuGGNN6ctHiGgLfOgUXOM/a/IvJWZzQR2Q
VnyFfGZzcOsd2ZOTzb5bH4Uatcen+UYSW95+ImNSmG//E0Xr8RnMfZb52nTYJ9zT7Wk2+ZMT59Nz
1rhQ9amuGVc1/tQN9kyGJ/TZMI9C6aG0RoBO/yQtAclqZlPV/3i3YJD0PLbKV0zVmzMI4+mlJCff
CVFa42lO57nP5Yk1lKUZnm1GnoP6pIM1Kb0OW5qweDD22Qt+usEYOHflnUz6AV48UqEmqYsfvbPV
vovERNiKmk8fGW+qCWA6oocZeqDfkmbEkQ7V8O1gMCpLIDl6DqeRCVNcUW+nETImup9fuk0uW0W+
1VLXw/E37+osiWHaQjxyZ7y5D9v1egjxVOd2VGbkb15FNPSL659JwhzgBogoS4hL6CfEmnBMxbn5
tw3sEOxoGfpLb9vPlEtYjYOon+X1AXVVHqYzXOdRLiIZwySDziRPvNixR8ksGw8tKpxDO8oPHLEh
eZJmYBFiGsr4edUneCyP1ADzFT4FKR6Tf5FudXvYPg0S+CF2ZfWx8kHHzZ2IJNlkzxBQhFdU2ZVp
sJardRD8KruT+QaQlcaXDLoi+eb29xjWd+Nj/RzYa/3iXDlA7xLmAGXsNV4zVKuMFLcFXbYTSiGj
fUdEhOuWFO+Wm5amA5GBp7FQlMHAqMEr9pfoq6wkBfTnlMORXCS3+enUE5UYaHqe3MTh8MAlFm75
LqVGCrXC91IXS43IXGjpRCCX4b0oSYE6Bq5G1oH7NTXiAWouoQscLShTB11kboXogKJ7/h+zH/QZ
J/DzJXTZDZekpryHeSMw9YcCpPNMBchQW6xMRmNDETHuHMSfKEMZRCW7Mb4NuakzIw6B2EdtXyoh
H4MZCMB4zlYe2L314ZX35YWkAjKd8+PRHuTRV9UwpytOyScCmrI76hq0SRbeNJ3d1gJeAxNPP6lE
RMNGvGjnlIadHTxfxw/ODGlYeEI4k11AdQ1LUVm1EHA56nWa5CjMIrpaaFMi5OhS3rfiG3DA3qD0
xuydPnmelip54OnMg2jxoI+o8n2glYUVy5NbC2o8ggshTZnSG3aG7/3XWc9llkhhgwIqcydxCaD7
KKE2edotK2LMefGaruGD1I7eMmcjdTgzcYSgMED8r5MT/oXNeu9PIbfKvxMk42lhiy7GozJq+eTw
8RoGO4XNc1fwhVffLukqTDqRWRf31JPoghZcbObSP1/6Ofr+kND/7CqVa9MT5ytBu8XAhCR9ULG8
/UlGmG16I/aHU1/vs1QN5YhvWROPDEZwdlXL5vH9xCn4WQOPUiiWzkbDJxaPRlgLSCD1Q2e7pqLf
TroXsKgw6/mBESemSGpBXJWCUyo1drG0aMOu/aba/nZcwPWnRKwy6/GleIQnGFOgtS81zsgts+2O
6MyPw3wnvd/sLz44wR2zCdx30QHTJEvi2ustQF9A3HGDkIeQ0Z/uSFTj0t+mkJVFGvUWUoDZMK23
D1w5yOn4eEJ6/l6BezLvhTIxqNrGtAoDNw6PQdOEpud1G5lHRRqoB56T1LBmAtpun2P577xWkoet
9uGssSS/kktBvli29BfBbkkP7WL2aZBppb29jZpHOqLavq6ZbAebR+jX+Vnos0ZJdk6MOwnlNuKu
c/aFDL/khvr/ZZelpYOfhwkU8zlelszFBdLYULGqT9wCQZdzUileBXDxtIPXQt6qVd1xuIt6iB5F
1bvsBemZxW21l5YBk4F0ggl2rqMTy1z2CVK9fVKk3px3JxXtH7i/CINuxK4kaoCWz3BsHiBgNn1T
CLe8d2rAFlbm6O0GMMN34UAkzdDx/+FCgKImT9Q9K0UU205yqD5EBSSsJGVh1M+4sIAcoO/rUfEQ
BXirT8c7Oqq7gP41WXGMsSFhpRWYziBG3QLfWNJVksBw8dePpxA+mR8ogigJRzvn3VZ8Z+DTyUJ3
iL5Nk1TQrWU93ftvSDrc6gG8RTsCPRnW9DvMMMignhDiHRIpgB7WHbVTDZFnfjAFthEp/W1i42mc
qZF7yDqnGxxsCAstt983v0oa9DfL0FI7w8pF15AS8MSUCu+9vgaKglMwPbdI74AQXjgAoXXYcJ5e
nm2OG9tZxZudbiPYjtitU4D7XJPSKRLOLd+xSkf0VPZ4Ib1bKoIqdUkY7Xev6JN29pUFSbnvfusE
Tq1XwOuMEml8nQCH/3L7An9iPtFcHRPVtBh/hUJUOIkUn09GmnScigxEatQndnezCS8wpWP3UQ2c
WNP8UGTfYYgyN+QI65Uj4W/il2hzOHmIc2BcvKv8DG82mE6RD+l1UzNJzK6qYwBv+lCzgoulJBNU
B5GPNyWZpp4UbgkuVHXyLvzEyQO73nb0tqiFY431dUGqcjPjFV3sYDtDY40zeRxCQqO5+eVU82t/
XgCruLQDGGvhggmKfeKWdS9W9RuNaAoXeIePRmNfYvWosZvx8N2IQAHXAPlRCTbFnsMjDNaDsOFy
WfxHCwKyp2dZVmuTUVvMaL3NfwCBRqd/TS/yd5p30mPoQFsaBk+HDmqLtIY2J5sIatMDC0cruJDl
vbFMqFz/3VfFB9kFPtBLPXCyfTcOuimHZIJc4+gDeRftzREyxVlvQDbvcO6cO2nqkPj3+LM5YcuP
PoZM4GawxNMK7W1j6ZiQmKf3YQqPIuhvnKXtmFWnKaQRj6V029l8jRCUOlUoYnMnd/FYU4u8rD8E
sy88sdOTUsWzA1m+EiPcaJsGCIpTzhw0yre5TeRFhaLBkv3ej+y+ZFligi7qdLKCOMzeKdHHXZow
wamccdF/31bjOgppWiLgupSkYe0W7rAR4UTZUvaUN52mhXegOxmwVuUfpnhRfrE8iBeC7BqVepeF
4syaT/rnWjW12zLOL6dXmBlvlcUkjAo4qeh6cTz8+9GSpN0k/K2IkT11QeU8Blf6rRZd7VXF3AIV
+WdI3SkkztynaK38dSQBz9/nvhlKgFVMTGNuUQG/Ur7dMSYqKQXxjU+IKR7zSg3gOiRQoh0C0A8D
fdykhG5aT10mivHhHPU5qPmtwFQuOo1zh98MpMcqb9lwwKsbfzOXLd6C3aFD1kUGXUu7DJ/EVmrX
TpuKPr/XO7JtdrWrLzldyaIzeYW5UvmJTzCC75RCANLuYNYOuasWF0BeTFw0WS9DLZgpbCBHuz8p
DhDclalWiTmsCPNksevB1VDO7yof+oMqTmP3R/NJq6kAQy3sJb8vOPfC5k/ysKyDNp+BKE60oNCK
wylZhtT716r+73KMk+3rCWISd50U0GTd3sKD5OXKlbnD8zt3kRUrqZUhloPbmMjWKy8mVS/N1gAj
vrHYT0zbD5w8E9zfQGgZ5XsWDNAHOtI7hBpyXXO7ZKXmXoCCeEr9NfVqL8rDYXg5e4bN4iEP8Fe7
gkh93KxFHSh8O7jcyb+gdd/DOQfo9MrlhV0B7Xm9XFq/4/RdHq1PuTgQ9KI3nBsCzZFoZFE8xFO1
dDeZHKRfjkaoql7IwgbJ+jsPPKwNoSR4rTpI9fOlh1RLudOlFF3sJp1rq4ZJ6yy6MofPS0WUcZ+m
DwUteZLpGDDFf6fsPqDjqYDgP0iI6Lcs7CguCAQTtUShOKMKmIsaw6oLX1kLVzl4VmgOpY24HZ0n
Op9oi5xQh6ysuL8K+4dYZPA/FkYt/s6x0VjYoHuT55+uH1Us5eJNdhMYUqgalnEm3oTfYBxnyatB
lLk1ObnMxND9Gt1LmIPpe4MgkW9inppR6qkOFQYomwFN15H7H2BYt7mo6WVN66eiJmCYeP6Rtiys
5gsMyK+5qoWg71L9NNpOWHUjdrs5jrbLuadY5pUWWaISLiWGWQMSKtzdtpaJvxgtSQsPXffd6K7F
hcMVP4MjFvEN0/Ic8L/b/H3N44sriE/to1c1CA/77FKxnG0Fxox0DmPp0V6l+vJTjL64atbokUGS
ZtEoB7aCu5hTy/hEUOlbw8iNrik0MSffpDvEld3vhrmTQtX1LrXZpQDiybJ34/fN023h9RatWJQa
q+WWhVpltLmtUUHnekSRH5JWFnpP0tw387XRcjWMPM/RhQoIsmXZ6ldXs6AzjMF7VwPuBjIhiWM+
oXcW2gsvEMfm2G90N9Kp2aAJNDn2uIBGrysONkFMIgNN85I3yf7rpIWDU/5NL0WaX6veKuBH6kvb
16CFtDJ+QBh+eywL7saSGli6cZdmNySYS7KbBzXc1ZA+JLvYM+ZHPCIeOqC9v3tTZ5CU3Qz4MqYe
/vtAEIHpFXgCRTQu9VLt2PdEhsYsf3MzCdcRxRAVLJf8Pg7ZnMSF8MDiaVHmcVsu85oEApebH0pP
AhBQWHEI5qnov5Oda9pQjsQDQj6xqBeKv9aUmaG1B0uRdbcDccl9SmCslXT8L0hUAiuvveSQFPEb
8uCr4eZRb0AZ8fDT84T5atbyp8V5fm74ARcc1SFk9RiOQ3Z2SkoksXZtxx92fUQVa2shdumQplQz
GBRymcyT1CohTPoPRjuFGWEPU5cJ+6sfQUVJXO00AXQuEb4SujFXEfKLKLUNUbWb9VvSKMrU2snr
Pj8eTwQxmgFrQipEpBKL7Nloi1An+tWpWutwLt4/8OEi54Z3YQ3e071LnqfrlHwCdfH8XBL7/ZJT
H70ivIU/eKXjh7HCcOnZjXbTnsqqIIgj/ASQct6spGFjec+dYWeSM9DF024GRhu0WgFP5vfzc8oP
227vMjc/3DKQtZiEjkKk+ezb8JID9FJ0/mM/06YAj6tmNjkC1dUEvsKENgGUy5AYUZeNpC0EVSlR
4l/wefYUzSGm7NKl/o6LdSOqu8SimbdPzWf6Eeg9YbLsVxnd6drFezMx9dGUJ9ujnJms0S8B6fb8
xbdQPzIvTxbofJEIESpmggr/QsZfVTuTNJxdQ9H2rcfCHwo/m435lxQTf4wMiG+k3bwymR2m7NTd
Ohqzf3kUUAIQ/FewidWn/6wU6ppv2uF6vsieihoguSS4aVAY7pmb5b7Ww+NnDIcnqgH56KZqPOJx
xRF4Cs1QmBzeLNMqbzZtKpdjjy0/GM4i82sqNkSufCIN5j+5fpdS58HRFkisoQGU3mzcPRIUxXm1
H3NUd8UkcMVym+f4bArykF0GvLH1LVARUsQ3Nyr9Yr5vYgKskRLxPjd0lKxuPvZg6cPJtVfZdjnb
+3ZESeCkPb1QLk3bKkJaQ1C3v/ApdkZ8JIHjYkjxsBrgJ3XsNUzRv2ijyPp6WGoyR8CXTctWWzX9
B2eIbsjFzQeBlGx0k3eZrHNc6MCJQQY3LZDpmQjm1bgG80Ysh/OkoTWuoTq8sQIjAXCfcqOj4wSw
x3HELeE83XWkddOzQ7JNeALmzjXpWBTZ/kUTes80C862vi+iB/Gfm2qka/XBxC5OWqGY+eHaKX/i
dqrTgRyU3rZ7XB1YMcZ/d/ted5emvfazKp/jx2mIgX2yMRfue2c38ej/zaUk3zdKUFWYMlorcRhz
uKDajN9L0N5KuitorY0ExUQ4go/xoqlWihp8JdH7bW5aR+R8sbAR26eG0uZ5xDBlCXZr3kRVpbNu
4JBw69SxMrR7UG4QsddN3x66WPqt2XBSQtOuZ86249HwV2Kam3X4Fa8TZOZzEukShvuQfRl/KvHn
JaM6EgIF3bex5cq7iLNIb4+V+HqVPPBUhL3s6dH3ti/EHCEC2ldxz2aw1T1/Ht4X3fE6eS14uaBs
kEmaeL57bUE2NXibpgyKjmRECiz+U87Jsm0U+VrZAzJUOlnVuBDx93tya5D2eWHFKRE+6DTQOgus
5+au8SeC8MTtarV6FK/cHTbLqMVFgsbkVd3EvizzC+2XtfejTD+8VRVxoNbiBoNOb+Lng+NxzWD3
fEMLmdLhDMGzgn/aFSpgoMTdu3KJ3zuIuNmceFb8xdo14GSnkaTlOIjt3NhoPVq3O8KLF7iNjAQz
mh4v4gylLmtfDp3mG69cEdILoQYlnyvcfznfMWpTdl58XoNuOT32TQ9GxBzQAqTVq3N8m3nbe56D
AIF04egnP08AlFiBb7Jn3ztrRSPnO1dhOgENJzcc1A9CTgc6sXogW53a/124Cx8fyXmbnDwPWPmo
C+eKH6zYYkxlMx2xW8tR6qPPCd+rAuE/kJBcJHyk9EFYCH+p0sGFolMCWF+m2C4TAxTn9h2g0pFw
U9LN0hAidf3wrhXhWqjE7S/K35DLncfSUbtQ7BgMsU89po57htt6GMLh8QDyflTvbek10eSJZPZH
V12Sssr9i/7oNIwioi12SH0gOoFpwPCY9GuOMCYgTYx4/b0SXmscpw7ik9Tn6jYK4iuEdwGaYUhU
ZMlXmeaNpE9s9/UsOXs4/zfbiAFjVJPAoPF/Gag0D7jDtBkyTVhYbCu/8hdhoFVQHclXC96tlEEo
uEISiNlMSlEWK6jeI/jq1A4xYVGOVEJakfA+pXpuUXZmbXqhzc7Ws8h3KqJjg0KpIQB/PGDfksBs
NwZ7SIvbOEW0h3Dt6/aWpObZaMGWswwJujOWU9ODSEYWnpLhKEEcK1bMbHbQa7kxE+eHiT/PQzxX
Xg7ZElVdz2i6Lg08dsPwggtMTy/MMrBbMiNil9yHlf4AL7mvmN0kNIk283G+uXat6WJVDpCm9MHB
nmfvg8xbPksuDI9cI6PGOCJ/pE45pTAmjRpcrFlKvpnpfzgB0qqwFJUcPfhe8e9d1weyZDblZ25F
ywMvEs6pT1bsVEhEF4xLDOPuGB2lez9wULG1X9Ts96SsToaDzjsYyr3UZ2CBxcTGIwPy1R0FgoTK
5ZDkvLcR/uexPLq2uv5Xe57NN4MlQ61OvlLwpiU/AVM4UKVW1XmieSHavAjuq0tL1oD9EUyXqZel
OYu61omSmzBo3HZGXDdtep5sm6y5gvEDZi+oF6dTQWk/EeNMwmWEtLQwwlQ3v8iXvQhJfvkWBj59
3H3HUwjxo7rJRIyiDCm/uTneaHYBNx1Og+LsOatl6klUQ5P/4KRU1fUwsLe3acXK1UZB+nFMJX3z
ZqgPUfcOwLxBJjfnsBEwpCNNF7FFRhZo5XPIUZOAH3zzOGP3v/bENuIpTO8OZb2lky2uaXJyFQOJ
n3mccp9wrf6Po8r7E5OUJdltguToTMSULEQsKL+iEP9ZVeLh4S8lx+AxLRnQuwhBDglnv/dEaiqV
ysKzc5Hojqru+Kd4Y5CEXp98jx/SWWgARBPQOKHKVmdO25f0UKyg/JnGKQKNAb52xOfiUIoOjRY2
IuTPd0nHa9JVSP7XJ/O+eDrnB2vlgVD6TsvGaWWuq1bw8WT57BB81JjJq1dm26sr6Bdu15V/IVLW
ZbvRE+FJ1889WThk+1yEaQA8cw7OYSHVy5JQdlNdA4LiaPmZutGA7yGA9gk3N596zxxLS8DAeD3i
2I/eFAKd9LlAIDH+rHqkSOUwkwBWUjWfbbNNM+qU/zeGqStdJzy090hbMCpYAk3BJYyFxGejR5Qo
6iAWPwXv91XIVWbVnJhtw8Dz251tmaMEKpQhJbefav+ZlYoyZ4kuTP3YlHe0T/rkFAZy5eRuK0m/
1uIEGfcR5blx92D1OwojDZHS9QGKJsmsde47XSg0Yw9ik9emF1JS0CH80LJ57p+vmI6pSXBQmciD
hx/ux3nsNSk+oSHjAv3Yibxtkcc7W4FaF9ZenNjd6RdGvTcAEMg9MlxN1MrC/DfVCfBNPk0H5U52
yXQwk4wrvLxQd7lhvyXv7udT1aKMlYaAWxKkwKLvpgbtFw8RPd2IWI8praIaveMGqt1HNWbSJORd
9/ARAsDchf00Ir8S5xzXKdFZmr87Bd/YyCA4ILwA3/t8n2B3G87zhOvBsf/abafaMQUq7LUuJ8h0
nOctSgOM44u8uTEU7D0VEzEif5UabtIg3N1IzjVqHcYma5Yu+PYmUrMzIM/ZzC+T+aVTfjnqkOO0
hxzYtjkoEQpDzqwOTTDW00idyv6elIHQ89xjBmlrlT3OdGXB5fIKqmNooaK3oZeGeAoCaPDwjb+Z
3Fo8sCKpriR+VgY8ixJuN4fmLf29qW+2TJP30Z2mSS2lvInM2TFLY9T3uaicAJCW3CobWQsEAt7J
dVbNON+UOBpRxFDY33pgIzh9SCf2HroqzZp07PSC6HK88zBBkgvGSIot7a6FM2BfQeVeqRwuOguI
jsW/gleuRMNyXJvxDGEpgTseoslnXa+plIlHtlKxTjIPuNxlGZyMKbv7eYNPh11WyN4tNTulYv8k
MMFpnmIRyZQkWJ+PybSfY+AHuk/uvgi4qN6iMKG47cBPM2AE7uFctJkOQYHu+bLEV50Knk+P8ahs
s+5aDbpEQaldzjB63RovF3SlWjH9b3rnIulXbC1Jg0JbOlYWJxpPmrEKGKWis5JcaYHOg/e2eOA6
u3gqEtWXDJjBj4aVXiWQ4gc82AOYfgbkZvb28xpGNeugoUr2+zyV6ZU2s6EF5eHwAjnz4LqskYhu
IbVWAl01W4/CLPVBaYu8dvAms4yeM60pmuH8nbRtmomwKmYJSWdLKXp9zzu1k34EnoBiOtXEmUFI
8BtVMIesg3DViwLLaYaud9bGzy954+N7CNF9fzHErLRkow3rI5TO0DlFVCc3QEYQgI2XsW0wCLVB
WyDT/oOZ3PRTW/m+LoAA5YdGZ7GdXsbHzDL2NJpTEeERQDqTCQFySkeX9vAaaRDhQ2Q3lU9b556a
DFl80Ml0o+f10f1TliWUA2IoOcIXGKdj9FV5VVJVnjQ1Avx3oskteLBgmx/JrMl+J3HLGnF9HoE7
EZ4w5Qcnxs7L70idyAmr+55eVS6UXvkSixUug/KaE8PtHH7YYaucy03LSXdAVkPW3N32tilQ8EZ/
AkYwCfqKb4qmJIKi5ccTjmHmPF3o8Qo/gcFYdYdLyOaLffQ98K1WkYE3uLul4QM9LgyX/4ik5HHP
A6GWkRC11tUJkRUylnmU0lJ9uMpYFY+9qzFlS1r8ugDMjcM5hgdm7p2IcEH5vPG/ZthykILVoSA8
PcPACUUoQx2KgIcR+eDYO+QO6pFSpDxoIiAvkVG0MR4thTuvXID9Y3nmJogxLMJDIx2TfFvU1icn
r0YbpLNkjjNcii5a656iwtaIDcoWhZDzewO8EIE+N5LYIq6CCnXvMynLUcGkclRjYTcmPjxxrkt4
2M4VaXzCek+W3tw1fm6oNhIBDRn8LJgP4lxupo5fWi1T5nvzsfqcWeO9c5O9yQ9jL/46FQhJ97FT
HKU4VVwMolVJsURhqFYZgBZZp5KCiUqAMVGIAaHS0jMw/3J3IhezVS+QIKpB5C2u5Czs7xCZ0NII
Gt2nGJHuSmFY9QAFGg9siDkA9TJB2VC+4T1tvA8skwcbXyVdgYhSCofkgd4q6wKpxjZGny/eFpxR
yPnSHlzHwzXwKbhYJAY3IjvsyWcq4MTBG+Py3P008AZax+5MZD1ZWi0W6zuBKyRbujfuk20Zajx4
FYX57gjP+Y2HpmUE6EGyHHwt3wLCsaClKxqv93Yi5SHxJwu6vXJm1PypR2VE+iOYlTiXdsYys/Sm
AJxD1GZ8kJ+bvOOC8zQ4w7PSPG2yfmkcokYQmT2MPiw2X56MxV6DgXAPXY/78GrSPDC4wX/u1kxb
DemAnbl99fyYVe9Pg0phtPrm04SgwcQ198gwQ3irnYJu4ALX1D/xxsBqCSOraBpQWMF9esPqZadd
gqkT0638UNK8On40vnUEzRUm7c+vzwvuy91oTPXdGTpo2W9OwFTwFuAAI/pyaw/IBld/zNcuI082
oNZMRrJf8A6woO19he6g1XJKmRIiBFZEST+d9itntTZ8mmHXIjedH/HESeLHBmGMWGDN4HKuF1vs
B27VaT8OMinuB/1puqP37xbnr5Sv3vwMVIaERqlCD3Z0tiDZHrcKIYcAyXx439FL1UQOYvHR5JY1
yU2gcVDQPq4+Nk8xHBxn/u127TWtcqUsLLWzOEAaCzQXqNTzHwGndtQPxJ2/gaMCt/XVCw4I2dtd
qbTLzV+QNhw++8mZTFGpyN1C89F7jO9lT6UTvi1imTWUbMBtVNG9mSsGpLAmaU5fjAiEqUlAmcaV
GLLzEhteUUGbiiZZ2nxGyAezcgly/Wok56AbGoPyM0BbWRf2Iv6Kqf5sHpvsaRPpQlrBU4aPy2zh
Zsajs8IhZ5JJ2yOCml4nwasOtlG5zpdU7Gx2v16uFIrjz7e7tWtPIawF9qXJc+/7f9HB9AsbGuJ9
Vh+kOh+pnQfkZdNrlWUGI3AMM47hxwYJIWrC44vFF7SjT83Nl4eACmrbgkO+qdkJtSnbbuiOU3Ow
eqGJNRoHdbA4hLHCHcg8BioI+05S3QHundXyocNesH3I7e9cxy9VGU/6EZpOOuFW33u+ALK5CBEm
ZlnUB6rerKKfO3rZx3BgwEdsyWnZGngTMmIk5bDb6aAUEakT0YpumrT+iQlsl+zHVkaFNLaMMP3j
pZoi6RR0DGe46EBqMGZRpNOHv5THkxqdh8T7VHwOUx0JwxJat+ElkPIbn8ZxAuO163M3PGJpPYvP
GFFOQKDDjqt30p8j4m6uUs8K0C6oxGuNdyWF7X6n7JPgo7tYy1e59x/1NK4Ad8bouboE1yKif1DR
wpSMyqSnLjR0PRVJCto907Pbak0+uZeM2EI6ri8yvwgdM4AeP0CH9aoSctc34yWMYdTimnMzD1tb
JBIhRJxbNfogL0Vj6Ai36HzNlYD8EZ552xUvv+USCPMQg7erLeVy0AkICh7+r/7mf+4Mv23dkOit
FzjwZqwtAIl/qV5ZszBsv7KGpJltqGigNRkpU6NIIm+JeJTXMAoR9paB7sOAM9R3eCPm/GQO9MvF
wuAYrTWkteZEMwOKupEu6nAhZxwlJfoKicyUuK2WKG5gkKTfFBuyeUx2N39F/bsvE9y6tDLDANwx
mXP8fa4ZvKN8FKZnPQgQo2nBRckL/YJglVmCcZQkm6scE6RumdG9uJ/1aJduvKVtKHnVhn6vmchv
9QPnF0QczAtazPgGwvYYWdrCA1LDB5Z+H6E9xa/r9eEDfAb/nXsVp+YD+zQgv3DzqF/GV9SlfCE1
2mtVNIQm+sosKA+RFzNNNZHjlkeICIONNcLgyNH6U36904xdE49OVAnkbNVMZO8Jf81rtQfHjsGw
vThbrY03w9EmaWDjlswprxsZq6UrHtT9SC5jXXoil2IZfVdmqE8cA/ej6PCz5Hh71qZ8RB96aDyL
3miTmHvcd6lHTb28NpiUBNG42xYw2QRb0luxWApy0TwEixl6EUqIQev6FLOaM+vKDDrSPy+dPfKW
rz10lSenakrdfEH3wTMV7DNceCVuxvuyY9zaalGAjZBn1o6XkMT9oJ8DGNxs7aW4loNJVGwX5ljx
LuVDGDuHYXTN/6cE2EQH4vTk+idZ5QFYWc0tsy3/3J3u//v0jgZP9b91aELZlXQnoSmDFDYQAdHe
iIVPsM+zEzNZgiih1EjIHcd1qj4S5lvtK4WpFreGnwR/Qc54nJEgKKMWkmosPzeBP+2MtMVUmZmd
lPAVF+iK0e4+nFpvjd1bEPHoSJa6+f3x7noMKC7SNMutMW/VABkppNxooaT9jEF0zHihkav+nsU2
xxO4qMEENIAj9UatMm75TGbPMnyC07hBfUtZf7AfCjLjFBzV+F3tuKpWrrndybk0uP3zK8A0ffXi
B6QneYDQKZf7rO2lekYFMGPGzom3ygNCPOyqRR8sYpMr6P4EteJ9L6iOR8d40Jrip71O1YZTxJ11
zv8qYCiMTbUQq/f3Ij/iJdnnXJOha/K+QjBfmEt6lDoCRmLPw/Fe5I7iaYjIoKVr+C9rfTAIwJhk
4uZg93L5jOejehfidgzrP8HwW9egVLea3xcvJCsNAugV9YNNgIKQuYop3Gm8gMcOuS0lVyPVJy2A
KUeTrrdNhm6ZV6rjjbEPpuSMLy3XmFTn+Uz/xZTsyAl0d6QVG15nHBlbYZAL6aakt/tHMcmlkpd0
sDxV9lxRmlTEHJUW1TU7SeaBCF36X53ovf7ZO2Mc2yeCAIHD7R2EdkR6wwAMVYbCm2HoHyzbAsex
Njpos2aBmneVWl+hXyqtTZxB71aqU+wSWMR0tywVFgoY+vaL4Fz3m38UPs0j5ya8hNgBAfYivPeP
iTqb0ki8Ebb79sojOBd+X8QQKg1n8SFTlvsGj7jJ587C+QrBjfUYQW0mp10B5rZTxbFlnumKHjiS
6Q63fV6ltRV2bTUpKXUWxA8wvnNlMEB70XPUYlEmkXdZ4tFhiERiqvh+e07ClOig9yrTwnfucf6o
iKk24cJSX/pkJDPlNrFH3l0kvQb5pfSo2At1JR790V7McUv1txnSJjleHw/HDri0R7QukMYzLQJO
dDmDjRX/WGhUE717heLY3IIcNyfwD86lXx2sS3Og6wE9UkSm29D+hxP5VmmJDSCkluddtsvvZBQd
DR5k6lHtO3yRBDokeQnHtSb4gO1StViylzZlv377eqA+g+PW2fWlbufAjJ4Zq1/NHrTBBcpfsQP1
vgiR1lopCQ1/bq50OnL1fP98Prp0Ew7NC3I8VnNywyBhh3RcknW8wyKRLQTqqVYMkDgdbZ6kWWDK
oHyscE0/rAzFSVsCNx0IX6yqMi4csussTrPA+dbeNZwHYw/VzHvQgO1Soi5yJBRYGqcTqgIbHRod
AFx+gRU6sGQG97MkUhLYLvMcsJjfq58Sq8X7uq0xjic1IPqEpDDwMi8IS2LgPlHwUTBqdUKbOqdn
Dyt0t7/dIXwtg6OxTIT2kTZCxL8HpWIOAkm7Wn2sF0658Tw6Mg4/REWGcIaujDt2xBjSKKXV7MIv
dnsUdvyfWb0nI69tk1Wyod3/VXLRkGyUY7PUriCjZGB6FP3xCpIJM4X0ft3He8D1sxA/ALkDRPgg
cPZWJmPkaRB0ZklaSfrr1wV4jo6a33rw1zfcP/nOiQexRoYt2dRoyYqfGxX0oi6WNoapD3XiZ8NY
D2E+MCvrbcxNeEZGgfzNwI6s7Z3HZL//X9FrkW/7yIMsydfNko6tkvpX66FMEXplYnr6vZBeMAKG
sU01zoQNRim4ZH92dEZjX1Y0mKtX4Q7tIPTTQT9KpUcAdlOptnqNZ38hPGuoAgsXKa+LF3jEW1FZ
3KSCjbMSO8X0qDaiwNwxydxwHbrjHBpmpP3v3QGl0XHXa+NE9o47y+4OtUQSWUNshyKzz2UPh3ni
LDVrW4gf1opYNHnoX57DG9lDARcZuA50SboBriYJGZPKQ4V1dNjbMh/OZuogk3m4f95Ry2dKYfmB
A6BPe0OfWUFTkTVZ3lQQQRyugV/TzVLCkEpMtmN/i4dzcgXKqf2ZpOpGfizTWVXIGLFjfgZ9erLO
JMPkI6DTIfjT3xxTuIqa0VWkLiqKXzuxpT7oyT7BtlQfIKCKAc/rKxEvPeTLcA0BHb+16ircAo+Y
MX32hXt4PlJ2popc70z6Nlvs4vZNzchHS8r0M8wq1/VkUXzOzfR+t6/DOPpK26WhXDg4gXnD31+i
w3dALAwNeyS1dDgAf6IaDy0Tk/fEfRk1nYuL1Ly/v60c4RztdDB39MIX0kMyyX1asRDwJsGQwLXR
dBhadfgl4T3qUa17FKdIFP6BftKlq7UjiWw7hQ3rB785P7A9SM3F9V2GK73kweWcIyFAVGsQIY5i
haBuuHQwdXb3FRCYy4/DQkAEJQ4OLJjPN1vhg3M6wtcE8huBrjToi49ORUAT4mWmuFf8qXCuhYVs
tsC4hz6dW8opPgy0SynMCTM1Dvn1sRj+TxoP1GEHmLH9GdBCglbdJzNp+ZprhIonYImiL+S0UpiO
/Slaz0Bg2gI2ZkoYAd/KqrxRtK3kOVZ7tzPHC5uoZLbGlqf6aGZAUNOBXp8y6DbYC4nhAQqRj3rW
8evr8j3U/I3jSGa1wD9grQ9pADeL1ukeGzTPYkVaOigf5PvsyuAJcG7s/VtdfNfTntfD5o5RItjh
rBfdfHebK719AzgMeQu5qNk8m45E5r5igQDy/AsAVpG8qBtSb9KwUH+005txjTyVCR4ShvFBlNGk
TVVQGCVVJvitJmb11VzUElxhqYrCwecpR2MPZp+tkaFo86TDBXexd5E1L3xHiIr88U8CmzrO0wyw
a193mrzC1Uxpj/q9ipAomZ7JdNkbrfyryS+9gZ1Nf/4BvjJePZG2qVMmija7GY7N4CLZhTDsD8pB
AChzcaXkQqFJ6WAxDB23H4ryVl9pjZJ8UTk7KEu4f8jpDzODzsJpmMVvIKNizhdMPh4IqpxB2b0T
jm2nXGU90Wy9Zs3WCd4J4gh586eUoFiucSDC8wkW7DvGUpG3cf8zuHbxZoUi/22L3yULskP7M9T4
BlxA74it0gWealuYfeN7ujXMU2JY9Tb20ETCdptGd4yxkmE9fAKz7zMjpAaaEWt9pXSw6tVSk+zs
+5/NXvpn2tWHRnMmmnU5o2e5Payn4QBlz895DgTJXvVUwXAE220Up3bESw+rMOnuIEPMLDubPzv8
1CFIjYUoD6BAr7tpn24RppsG1+bgYMs7AsZ/kxBCIb9dIplW6WVQ6MU5UcyNZKq1fTkJNJ+bEUu4
d411lacb+85iDZlFo11QCqomXw+H7OwueXxJrhzcWNOYEN5f5z91hu7547dT7Q0loMDYfyJ+LhG6
okRxbB8gyHzmXKUG6uIIrLoMKbe9kM+skrdMIImzTKFujvZWBd8dw6+vH4zlZ6UJXgWJsXUCplJN
8Et5tRZwfb53zMQdgYi9c0CxWzOvzgh8FUgX4D6kyIe1tboKFJ0r5E26Br17aHQPF1f1sVauqMAs
N5es5JQ7tjPcpZuI82Wyh5gSJlxI6PNBSlpZhfOxw1ATKh7dIANmX6b1NqEFLbdeffgXZVvM9w1c
Pki999lwvL3gnz2VrEQZJv7jMIFXt/BBiVJd/9OILcZjMRQdRIGsjNmKiS37WJxfI82SR2Qcdy2W
qiJwKF35Im0gUMgmxtDHBPipGSkqUvEcYQxVfJ6C27tmGOtBdfRlzEwe2DjlF8q94S7MlpO9QB0G
r9yShvsGLANmqVy1W4o46qZ2DuuoEYXHL9LGoOFyYIJpq7vRK6vbYihGFpiFoxcuRIwcM6/7DnZ9
q36E3gKT8dk870nwxH5lXZhEbNCn1GK3igDnDOe0kSvj7MUl6jQFlxA+Led+QCqUwccZ33prpWKa
GvlKn85xkSSTZX16/tJ1NkJKUH8nDLezy9ocwXTGz49nFjt/kls6VzRlXJ5uwF0m7KIni90g/T4x
wLmwwk8KHgyw77Hfu44+u4SuiXjotTK05O1WKTpyDYfNdW8Y3erKlGYfqfHHKrr4rOdV8ipKqsGj
fY590t91VHyaDcOk5WKw7MQ4RQxGKCjhYIzhbOB6YJJcU96w+jL/ywWlclDQgx9/fnA1CK+eTQgQ
u2BMaEYOGK5Jxfrmnh2lHUbXHUKlnAoAoZ+3Qu+o3B7r5PzpYLnVacEW/tLjy9UZPbHkKONn59Cy
Isx1Ps7pssX4OipqgoCGX+hNJ5ploMiOGMr6tr7h8VX0S8CDJY6cMC3a8uY2/XRcW4eQwLVPaN2R
W0Y7M1ye9ej/odsRS4ole/Zr80f/Hp5IDLhVcPelzEY7m/IaQ3Dohpe/e096neM+0ewDn0lmGZza
yKRyLep1Jlva8uu89kPWwaLL9dAo041xu5gilfsRHZE1VOpKGtA048NPQN5bbd4ieQilvBaQ+6o0
VO8KR7QXiPK3b33swrfPngkrjpfPvCEBq1WuLT/Dv56b8dFL7OwnOoTzAUUbmUP0w1r3znfflsqI
FDHboCmEMg/6Q+r64nvWfC3d+M1pqbcs3+hMzqQ9mVNm+o3u9eXAQVuKjqaM16Ros1mTI/5J+FQT
YW+zJRSiCB/jqtrxvnbmcSYR5+RO8F9iuq1FF7QXf6ujpYABWu1ri2yS/P55GWDjPpARLLev+IQF
IvCAGHEhwyBus3zdnmF3WFbKeIfbqhpImbSX0pESx8q3XwjV6iFB0duXuBcqBapktp2MVCEYbUYC
Fyb70vLmYHOPsHkTQKAoJn67wr+e+WLcgqUYJBnaHbM8jtXrP74sQld3dEmmLw0+M2N0U3BMzq1w
9Sf5i2Cgst+H31kV6e3rN6C9rOwGJlu7h+3LeW1BjwSoQbvzthtVsF2q62c0AeEDy6t0wPBkirDg
DKg/mmJFgeHPApOfXb24XTid4m1EaJIneiA6wvctPJ2y03jhz96P9UiAAqrqE3WtRzhxcF6f9AMH
8ST79QRqPC7aI5VwKQilTtWAPxUK7vMdUuvdv59XeANesPe63CXHZ0gkIkTGwGJKFjxlXeP/hVbh
a80RgDrWKpjB5azP17r4S9SH8XERi0l5exDLXjD1cht7YjdJzrjWZzbJCdbEJtH8OXfCIyQEMoWJ
4YSYn3I2db/QprFEbsZ2yFYLfGh7/cRVow3gbOJaPeTyiCtZR5FZryxqADkakFIdlNgR2qOFapoD
Wjn6i/ynptLXIEysI/PZ/p71CjpbiKSWyEj17PkAWz/v8v0m9RubHJ7Oi3ccp4llSSaStLFIhavz
eMQDoywAUU8Vs4CkRPLW6HSlLMp/uCjJhzZpGdHlXkc7D0QYdrwYLEuxebYNzz4bCGqnzssbfiN7
aH6NlMJRQ83kUlZybBj8wz12b6AWY/WOlOHaga0kBULm7e2qgvAeJEt90lXm86cSk/NHtV/KcCHQ
16/QFw5MXxz5nYXKZBPIBTT7f6XhijCJRq9Xghz2j7mDZPT0epEgTuqaHZbYR+YiNsWOQxsfr3ZE
5HpS/qWjOkQEn40yzocAavUC/OmK+xex9nDwyKPBKSSe2wirLAqDDle5ageA4IofgMbtGRL3lIT4
MmFhC9/6+ZvYTEIEnFTMefkBtzDkhME0rWoRNkHcONTTSirFjLs2v8y1DKDxd0N/UTuEAhZ52qBc
W0s0PzlatXx6NeLhhy2D4pLd32b7/8YiMz6D8pR1oyJOVaYytg2b7z4tYZj/bMl8s5+NsWCd+kWa
qDklqo7tiEgURwXI/i1uWZHFcqvly2jtr2GWQVGM3yHiQBqKlWaCj6LuhzcHwPNAVex9FwPlVh5+
0DZT21VZo6vZeyLdJIPI7/s60Kvt3qbbfGUa0h01s0P+EAFa+0gKAgZ2LLfjXJ9MfKnQvhE7PByO
lzGBhcC3zAeprWYn3qV8IgBsdIjcF8nyApn+5eHXlGSoniVEbQRNHr9SRI0846108PVMeWaD0Zed
D/gAk24Ydh1QOd8Y84MfHokx3tmdNjECqFmz/nNPaMxNZtv43iwioZBU49SPJIaCMMUwW/1ingxT
l9WrZ1C5AdoFEtITyMbGF7x6YCtdox7fpQmACnInXFBIuAcliSFe7IMmNLy9mRQKtY0TQ9nFEwpM
IYg3WJykkzfqk4Z/e6wgKp8ZlhOVGmro2HRjxkmOIm1ek449ijDydRDslKP7ToktjMabjQ+sIQ02
WelHf3i3SPW2GF3HKUAFGwt4IDUK+mScWaqn+ZDSfXcpSSVfWlpsAbnWIr+82fRbSbxtvtWQ8JaJ
eA7qV3QFKS8P96Ly6kbXhHz7E+bp+nSrGtki4m8L60k1yaOJ2OMdWiWPP2dOMyx6GqmTQJJMkR4t
sHPhKvmn99mkJhLVzPBa2XR3qOamkpS5LKpwWdYa+nl9CyKPwQtgD/AldqssLOriWqQbmVA6RJyu
94aYG/loVbTc8pW3iMUCyLGYwt81Ndt9AbtAF6lDqK9sUe8IaBayHoangCG9a1LZHBrj2bA1ScPG
GUEJN9Gr1FEysZyuEavtQxPlMenQ7d4vQiD/jg6X12mZSkHY5t51Ov4bf/J3njhvkyrMe5Nro/Lr
DEin4BlD3Oc3J7JEhE2aT1divCNEm53yAUhLsrQSVarc1utLwa+mLIHoPQmGtx22vnMb/a9pF2jG
7eJNJ/M+ogqUVzU7YaZ5FAx713Zx+aghxrWpCVNqg42NOZNRS5AVkAtzZCHLs5UaKT59r6E390wV
N3KXcqAUx8BRVVwA2JwrOMJUIjLtkRhRZ4vJrSju6N1MtrvH4bofrRbxUOLyOP9NI+EeAxsoZKa8
RGg9gBHnaBSFhfqT1qxx5/pgsiknBMIvLWHYDQj8CCa4quv2YaBHciCK25D96XjIpzj6vgClRo1q
2ZunKSmqXjkatxWIRBhCItBCIkvQ1TkScNAbrUCX9ptMVqaFZbT5PwYSAJDDZkeqAwbVbrfFg0YA
D6q8GnZELsUSfQueVIu0P6XVgmRy5MhFrwF/CLC1YvOOoEXVSvxsy8yQUqs6w1ZPN9xv4WCDByMM
QVZN1N9xc/rOoNweZfsxSTqUfLv88FMxqX/wZmVJaKcuX+1PJvjvKgUAlxNZo4Nk7tIw6Ua42HUv
Z/mn2PgWuCn2XD3ZBIjbNOgnXLJoKFC9CQMgL9IUUAZXzRvgW2o6KaTMOndxqBa8PbdqQBOTFkri
27wKozFoO/SZoyzJIGfSxgvnm2dN0Q0qUiFMOA7dpO3L13GvGCxVGsR/xuek4qR+qb1hs9Umfj82
F7q+ljc1jnXd4SAd8YS7HNKQbuYj3c52NNcbMmojJdSSur8HHDGumZDwjQAaQ7zfs0SO0hR3e3yF
UUwh8/W5ce9ztQPANiM3vPrDVmDUBGzlyrSs/luKXVQ1aPP9QOq+157m9YWkLcIXGXdJ0U78Cd/v
+VuNkXhfQzYDD6QRqk5KxycfLkyQDZsMH3BXlJeOGDpVHRNCaSA5mrGhfZpa24rj4YcKFi2zYoYJ
GYILcUIUwvaxtMdik1xvTPvIeqGb6TFY7UIIekhfGjPK0F6xEs4fhiBjjRW62HFV2mPRhgM2oTKp
2U3g8hVy/fRnPrMLCTEIIcDJzkIxkhzftgD3HvfyQCAQcKEt0aZurHTB4pA0RI4W/fsUURb2S4Zp
dIOFkr01Z17jlMjU9ijpa7iqn0036Un8HLGjod2qPnnIH80ovCLdscPr/HOUkF0padRAoZdUjO02
QV0WYLAMfN/6+ZlUf+IxaDjmjBxmqERoBAhfkGIK8Jesgxm4uhvM8nMQtaT/xavsE0J/BikvVnCU
FDxMlWaTECSOleDFuMbrZxRPhT5+1/ZCqVlclctu8Jc1BBJqccQgSL6wUJROpNVxbLauyxGuGvUJ
cMmlXcue/biGS+RbxNbfx2+lG36qSttIqOUuy8foxvW20IwemdM50DGFxAz636m9u8bRaDq20SnJ
i3fb6hbxg+QPdMnCFaK6j6wsSdN2Z9O4lSjOJXnWEJJjNYLpnL2Pw6xcNa1LDjnibShLUOxWUrlL
gPBqfCFxyvuhKWH2qEjbYXEIuRIvu/hy/khXwxXgzp+/TVZG5EgJ4DtE0W+V31IG+mPPbgh4idnQ
o6ycpo1XDCM6H04K7BbQJ6+yZRA3Dq/3Du16blyYx1gJ5iUdkJWG+PK2s6+DHL0GrEKO3Krb9TUF
DnTn+BJ1E8yXf55lsgLOWTCvyBYSzfAidNxmAR9qVeVU6e6K9ocKedJ3/0Jfut20nb+0M1wbWerW
NHoTQ+qKha1tS7bFbulUdOwdYrs0THN5bJVrco0AJApvJeGFZTFgxPEwkl3qc5DcSJUveSXZW46g
OSgkccHF5ioWxIFxnIddSOe5OAfBHdqhNoA8eBaKXBc8w3dBgDEKW+0yKicOXa2xCkecVPrUwMB4
4x+08xI/rH3fGksQdYaDZheEjXJYr0qU4M9dG3gbQLqpbmLX+rnrl5fuMmQG3wPMvnwVMoFUBQO4
JwJ6tqG9+d+Esem9MdUDXPWBfetFF1exbwP1+T1jfhbSZX11TSlEzizJpBQg5NsC1XaH32Z37YhH
630jzu+5mDHhCpMvG5zRBYR1PyzTlK5J3TVNrl5XVFsEKmYzQZ0Sm4prFPLlr/0RgR/3vcfvEUrZ
KY3tWDi76wqDlRez9OxWY8MKuOqiGAjtkZDQZp+Ez/he4pZODytKlZQ1apziMGzZkmasodkkZN7Z
BqyuQgFacBHA054RIcvcdcyerLXG1Tf2qMv8/GaxjleeRnZrs8aQpCv13R055Z9WS71f7qme4zyS
U+7j6Qi40hkuW3pa17Di5eOvfbgWiPHbd2QD2SCM8VMCMr1+gYj27V8RacTIdpOQ5DTG+bHbQNGD
zmLRJRMny+6aISuCmpseQeAy+E/Au9Fb0PznuEGo5qnOGyvDhz5s74DDCu5SykzOYOYOXxvcay3i
ocuM3CMZmSK9EUIVNdjasFb1yFy+kUrpwKhMnTLRRkIFrsjvs4eD0pqBld6/f3racp2KBPbKQ4jP
UCpe6O0qNlpCj/Hw7tze3L8qt/y3Lkii72ESM2fpqlV/Bb/7UUeJ4D5MehBQHtaJHilr8/db00Ak
eqmZlDktUykERHiN9FkkbMvjR/yekty7NDFLmXZSUfSKXo03mENvBXPM3hCOWR3N8IiFmLvg2fh1
CW0MqpuGGEQ6lZekFO9ei1M0ZTV9snbiB9gsoiYV9cFC+Hp/guRmi2c1RiXKFyq3qOU/53JwBgap
7WoFuoNceNB+a/JSqfdEMCuEgguwkeBdN/UoxYs9lYAKry6Y4RhJKgbeMyan+HHZPgUyTsBcz+Mc
hLv3ilrLxseOGbt++YqWldID9M/hVsMaa6+Rj4zgywhgbKItPySXtiJ+fD08Z1lT0rK4OPaPsiZN
pF7tWNTXjG/7DlFb3BfJFGlgaxb1Gg4gVTaEzSVtbB27RU/PWY0MAnvXtJr/FAfDjOJi13NXmLLo
7GNvs1t4Gtfxf/h3vplUA3DXFBJxPjtpOZ1x9mp/eICpgzhRJhHcFGJutRs7pxFV8JkY37g+8/TD
THcqyBSz/eqkZ8Ub/wnu0ftVrG+A9h/ybT5VNUKSb9T8rrXb+5dLNvb7x6gZKujdfUuews9P6kmB
CoIvV/3DhyUwMjrkgPuL9Mv7jyCHXa8FDyJLl/7j9JcjEzSk2EphYxvbbXkn2KTNlX6EDIXRXNjp
uhAcyAoDk+6mRpPjtrDQIsS9hAHcQ3Hn9tBAnR+OykZ0n+jDVRA2VaaK/6WsjPgDFN03w1cGIpNU
ZtpcvDArpl7Hp/dAhr67+48NSMRTXlfEMMwDDdi35B33ZTn/IT/eJRjQfm52+RztOLuR6ouYYLIA
/lB42oPFA6qEsXTomyDRgxkW4/Q9oTsFapxZ/bh0Bm4MN+5CO2eqicY5bThYAXNFF1PIkwiFbezo
CZ/dIFcnigfO8PVJQXh8s/gBc8pEy0kuEoVHgmm/vZDTbVPEX4bgndbmORpBv3AYU/WSMRq1mitQ
EaBdnR2UAy38pz42y5q3dSCLJyFLk+xIR6eq9Q4lhxQ87IMIMmBxNNx7oKeI8fbKyYCd+Uv48VK2
3kXCtW6xGgnLnbDiKiGqblPaTWfgbjryJXqccAr1Pi6jF2WRrugjL3QVieAfYFfoD6uCL6XmekbW
c0GrqLZfvd1oE5O1w/rX7kwHAO1SStGB5WsSoexpgxUShxKvvpGIjiMld+My0m9lF+PHGRFc/Szw
ZBjV7EP1YMLr4/d/6d60rUXno2YiHqHWN2VF3Pw74hihRANqDOzq1F6OrNWURyz7v8U/LpqpjkN4
76pfdS19HLQUQM52hd8MJnOYWSEAU9+z58TVy3x67WXHA79c9DpsWWo0uYZHWYtep/DhIqVAFdjL
TzpKOsbYOpQaoxar51GfC6lAKkKSlxVVPvU37lTqhkaEG6333ag3ZE8/boF+sqp5UMKvMtsC2fwt
I3HOSuhShk5aTnyWuXhJI0rLCXw1fDthl7y8I2KBFj/q5wjJXGEVHAEK0jgpYj2l4vnJtdDfRfkZ
qhjd9ge0cQ2091V+hOiAM/YKNtdF+pkj+q3kON16Pwk1C1t/UbAS/SjWp+ufLn1+3sz2zLnlear1
KXHXbQVlq5HK4eDVERpOiEo2s4tod2skmBWD2nooeJ386touHfgypEU+8iqUvF2qT9wnv/EPvyn4
58wEunDfjoqn/zFdxDnuGg0Haflo/tv6vP+IAOWkdwxTS5UjB0Oibfh5zmVwVpAjoKPnb24nluLb
9ruEsgnDJNRVXzEWe+o53nPALlqroP9KYrSEzCISTPX7T/Uj5DfrtvcjCcOV0EvJm0olcEsgiyrB
26JK7elOINZoKEd9S6q4ZuuN9kmXDt6lbTRAOW4wL54XlTODi3wq5eA0SVe+EcBoiJcmsyHP4SLM
XUV9yCclU9DEbbbzKb+aioxjRv/r0l/RtiEKsYbEIz3/txLFkE6succmKualnouO784syY2Ez48d
uUuceg5R8d2TLej0d07ZnQT1yyVWJPs2NU0K3QD2hx0jk/Zrl6G5zJRo1ioR30A4mPoW8Edpec55
oh+kC5w3ByJp0DXFMthboDINssh6ON6TR3BG3hMYaIpBeWHdUBHBJUFynAUpGhRtXI1+E21LsnSB
UzMqrQM/XtX+2jBNJzEstqsg6GZX1k3g/si5HWW5+TnamctxoDu6V6FnQSLRIkEqU17J4rI4nNoG
XYstunYb9vZ/hkil7NxInADFO8MtkbdN55G0JdmmNXSIV3ETV1UgVAQHPlqwFfgxHVRJ0Ypy1uup
G/gXK052VgWVCZH+QKNqhpFeE5+AmYrc9HeUd59/rW6d8wGGzppz44P/Ht3z5u2G0dFHfUkrsqP/
HIvIRmyq9QBMRTRniWGqdgwEw/SZQIeaKb0dlJiTnRQXn/HgyTkagWSOmYvbhN70Var1QmwAiTEb
VHUwN3ZzRmKS8WZaCi8nHzIiR5fVCf3k3LoYdg0TDAkgSYGSVXyGBu/N/CTPDs2P6vp0pHucVbIb
gaweUsyFHsYYwueVqFsO2bl8sO5t79lNm5ZVGmkJX5kgsjK2AU986b5VVW+nUDOdM+0zASKWmPJv
6GBV2SwQAtOFFb9rX1V0saybAfFvwNn9+bvpdYn7GAMs9n3TWb3lv+KYWZGvco9EeeN2vXJbzMpy
F/VQEH8nGUzhsD3pemnn5ScBlMpXz3jcNShs+Nwsu0r/QtqglottiQNe46JOQ164imeTWHNJgQKp
8kHxf22/uyMws83X8rPGzMQ8mnDILyjkOJuDCK+SCW89wEEQ5pNwXKjh6i8cocDjBWDvniqyH8Dn
CN+I6FeF6yLBoRNeonLM9XSnD9hU7Bvihu914a9cGau3elmxeWcECyCE0Eq3dK0UrPGfCWDFxVUS
8XlMtc9t2/iG+KpcRazrkLpoiAwqKc6PeWw/Yw4zBja8h5B36lvqL4dsWancVnkdLdGjQT2uGl97
QRhmOgKFXPs8QDvEXWUmUqwPuSHcJCuJ0RYzSKMY/SPPDNRAGLliZby0tt2U/3a1NunQiVAcy5sc
9JGVlJzw6GxO+oSgGLijxb2E2X7ZOPtTSwFT+uRpbTrNTxIifqOWicttOv4o5Q+DAWZLIhDRpkx3
I6nHAQaZG6oiSys+c2+g1aTxQ5VIf5lWemC3QYeg28RUZdDW/s+O7P33cMSJHUj8lNLk4zJditK0
81P3vLJfAgAZpQCS3oNwBncSdayUWvefgOuxmRNFlgSU4Q3VQEu1nJH+57gLa2Gbhs/6FWmknDKg
3CEijkZtwTFYTPT2Okn2g97HA7bNyhrwu/Ffyz2lfzKLxeHQBgnL1vuNdmxOgbdVmVirj6wYOrLl
2n6yl0U58QwabukYKTmt4b0AiO1vS6Zv9CDQpzPImKegRuMX4oIW1fIcRB087S/9keH+yfIyNNSv
WK+pOVeFm8n1NsNlNtdV1PrnRcI5xi2EFPAdYxDow6qySpq1fReEfPhDJTJG3kl9pHxTIO3hqfIR
8CmHaRNCme2SvKtIWaUegenN1R3G6WnC+hk/X7JpVW8ILKuNuBSJ+VadrdyajUaxZsYn0qzQUg7a
Bh4WRgNl5fRGTxJLoSMr7EupLxPJaDHT3wwBSmIm3IbaAkrgIZvS1T6GhXwJ93ZuNPrYzzAXVgoq
P0PF13vtjZnAImkv7KZZ/qYy+D/cKHMx6+UoNb00DIRX3hWVZB6FuxuibW3REcUl7avqnEKpg23w
G8kVkGkXHCX0HQL58Rg5F8CtaN7ehxNV8uU4jZFIwK50gDAB3a2OZ9bnD/ypaIR28kbhPd9vTOBd
gd85dohye90hQPLhrmWju2NYeUG9o3EFJJQaVB/qsUkMDkQOGALpX6puvPzW78qbdJ+NY/qemWq8
tDYA4TwcJCuX0RH1MVc9chFGqFaojRmubg3srzdMkD+BQ9/cBArHJIX0xlAZAG8YOJ3/Ng8DCMj0
HfkROO+piHYhsxm+L8SpTq6i5EOlr1wQGEwIroWMPksxZtW/ITaXC8rOz1CrEXLK+JKlQQvSoD/Z
YvC1XX6QnQXbjzrbUF0H+2ydNkeEcZCYnj9oot49Kntutjl1MUOBbdfWb+FyIH6IkB1RA0Zmz0a7
OMIyN583pwjMopJ/BMXsDpe3IFgj1cVGj9nTYxRGHTIFADnk8k2DBfp23pJcuvM73hnVgX+52oBV
c1NUbVEbgv9+jYx4UoPpLOGVAbH8x4gjTweXpRFUVOtXrxLqDqRUDgOSZSbKbOC6tIf3vBnrwrA5
dreRQF3KuM78lJuWZovDWUiKx/4Q0ZcZe5DCibBm1q0OwODROve0oHUWNOV4gQKCHeue+nWzNTW+
CaBaALL5cenpOVRrY82txC/tivjQf3gw8cX4McLGCEoEQr29OInxl0oayuZW7egPnVTWMGog2F2f
Br4hD0bNw0oiKXw8joDc/Qrdoh+4nB/dve4zQMugYjxcuNJvdg1LhpggNftqNkt5+0FbjAn261Jb
RnOvbzSHeqDYbavAXyNXgPQr8vRYuhP+uz6dJ8Dqb939kzPQbM2NsNwbxAznKezJH2lPBOc7MPzC
PZC3VvV6BXk1N5QAC7/4VpACPS1SNu8ofQxg1rCWifsGt8coUu+MnjrHHI0bDW1GgdjZUruhsteX
0O1c8ZGY6XBUVB4zUTcqBLXAMWgbAcTQs231wfUFrqRktD5AQ62NmhYQZkywmToCjIvkQTKUeBwm
DOKzYHxXH3mkepyPgyhZeN0g5d/iuKnjao6C26Y/RQ8tnuDADbxAdpZ3l2OVRtC7h6/JKAkkxzWk
mb2nt0RmeJzC2UDDvkXllRE+zl3tCgHyaih4O3BaSI+qKfwIIEq74lv8Qb27laRS/8zQvwUqASp+
my7SOQMlchIAkht/a/ONnTqh5RMZnEx//SgZLXPo3eUVgxun/pW/Q3Irzjanwq7i6qBMoyhthEBP
yW7gWA3N1Yji1ryh7nBnsPq4mFDs4DxkHY63RLyXi+fdZkJ7M5takySkgiCIHSaoLttHWmCk2ixW
gGukMFQr02Db6aBEINHUl2Zr0Sf8UPjoyXhqc4VufWh1BfENkTMn+BcA+Tzdmo37Fy6vis87YEh+
jHsln2j5eOibN/4M58PV1FJoYxk1PvJkesB9O/uIOsct1dHAqFi1ECCJ/bwLTOCi8dyEy7HF7ql6
2pmR9CGoGS/vJFsrsOUXpk3Z12Xdn8X6o/48eg3XBmYfCBO5s1iAC3fyaDNQO6CGCV2VPbbKSMVM
c4caPE6PHXkr7uTGzhhmWqgfOHyghoaCjmMVNYCJY3omiZ4Z+6HcNWZR/jDDlB3kDTGXKfuYY8iE
y4XjUHpGx7mdCPKlBvabVVAtsYGPX5EqCg965MGs1XdOT/8cneJh0WjE8VvwI7I1IAbnidsAQq8f
5CdfZJnFryAQmeVhVKNCNKLx0rymH7S1DcmlVNe3gqu9/LeudtXpnGjRA9hPP5eyAmBhJElnG7uE
DUmLPcJh+z2Es3Ye87401+iVMFpvP1c35W4GLhRmC2Ap38zOsrOe+AxHoRXJBCT6HkKaU67IP3zm
5uebJiBBgJ6gSBPAjn5C2HWrjD8Nyx8gdqD9lZ/9NRtC9L6k4xbFDf7dFCWv/SCK/FvJUXY6Kmup
qqVDviF8r1YAScc1rKvanjSSZWVRecUZqzh1P5IO9rjTi3SlsXtuxFJlFvkUBD6MFB0ePjVKbUdy
SX3JOwDkD0iJpDRVh56mImgLEpwv5jILRvHtemYBWdqXuyXEA13ufD0uvWBwYHK2oLzo8+BJN20O
pvhbNngds3LEb2MG3/V8w82vvY2dPc92cl792qskdxhsB70ZZAOLdrKjcOm1xldK6qqTACL6nvrG
3LhgNxhbUms9DX/XvoIxkA7pEavQqLcqugfCzV4vzCPDf0jnh2hA2+NMcpnuTDPWcOs7S75AETLJ
yjzXgEjZLsAeqjMnXCK9U2G95ztDoP4/9SWRI5+cvO+0bAD3uD7vI8K6GEFrxuDhFnnUSGwZFo+q
PH4ZOXZlh1dkFfsNShANCjeJ4EC0msnUdsC2TLO0TiNrK99VQFruwmDjC4SGVLOhds8m5J0ajiQf
PZcrdChAygndWt9gGOI0jngvqtNLyiReMAOlqwG97NmyTr7oetXvDxAhQkXF2Zq4N0pKUi2M7Nbc
1Dd6VsLCbF6N+Uay+0/YnxPUG/XA95pik4MYqJdgEuIFJaFIF6g+xd8GOVczBG8GSwsX4Q97ZyqH
BOquza652cgm7i6pQpIJlIi4mXiNMOKtdEuY3MH+QTb3DxqyFZUZYkK6BPQRTxDwRYpHm/kw3GUg
CQG8TVVraU+fKQKgQRR/6PQQVkeXRhz+Q/xd80AxO/lOr8fmOPMDT88i7Zus9VDdQJbVyRmHyNsB
vvFIy0hMCFHVgeKMnBH/4CBCaDtYN2jWqOdwX+x/juwJkNIUEfR4lF05kJLCa9jFkZ6j85dfobqy
YBJq27YbyvPz5oAh55RR4BvpBNodXwxt6ToNB6KwEci2eR7YtZ0qQaYnubBpvinzpzdqrUcN+677
EoymuKQJBNeeivlFmNsTC6gVREmnVeDqn45ExOPwG71RvZdRWf+ti55lUcQYML/VEYgo72o4j0IN
W98siDtaxEoG/GCXJwkiK5ftji+tkI3BZVNiAYH2bSunveyvHovGasX0AlzGQoaZkehd8XRwKfCZ
5+I34RMToWkRsP1LMMszEsdP1uCTTrKVqrRjv8FsFXZgtAdW+PQ4S5ItqdBqZs2Wthly1ZzAvtgR
wrhFi5jyQlpJSfsLRUILh8SRPDtU7uhst6pGo0VUWFKLTPkGvGxnT4S/DNtzb56fPl7gPUOw+XEJ
qF62xriaZUTzLBs0jSug+WONDqdAkN2NR2pIbB5LNyfsJNocQj5aU79KIHHCpAocPXAeMRi7hOl9
2YaL5Hq6YxVcqKLpoMyq1qj9K4MZa/q00ohEp/QxOSEC0GITq564K6KY3vyV3uenWdNo+l/R2O6w
WqsQeossFJyNNw9/lPgSbbizCrW+/7jrkIqUmZLMziV8hku+VqR5ortBouMAt5BGlMF8waw53p4x
cp4R0VFet+3l0A8YqatkR5XTVObtgeDHSAzS9UsDl9lYPrMPy02igwu2rjLkjyaP0W5+IWvcxcyj
3AC8/g2ykayr3G7eJWsAJAodN5CXypXwAlnEzHRw2AfzpS0/yqZt1YKRmMpDJLqIUbapbRUO23b1
51ux2qUqGKFxOtQFmaN6UIKzGgM8N0Ptkgz04sHTDPm9wAgpQqX7xFamedWMAeTlHi9cBRTfocEK
cbBOcVYUfOBB3FXc3XEq2uxH3nCEHTzd4yTn5DMC8/jac/uCmCM2wI50O0JSVTFkL+TqzqVEPHcT
3S3NkORp1C2AFyeY5tG1rFGsTy1+FPH093nWfANJUeSVBjy5p+mCwiNx9HrJ/feJVIcNj04ctbqf
OBpx6pBdlFw4gGQIr+gcOBnVPQNFTWUiSfe+STC803uwWH6N6MwqMfzIahSBXXU9i6WIcTYBVqNx
dh1Yh9eS8B5ii4BFDfSM7oPPuxZxs27e/NYb5rw9jGlymq3APZxuPdKTwWj4lOzOuE3MnLFMkMHe
tgGP5FK9ICL/n/BT1rhaETDixYbo27jwdS8mAailOpZ5hajyz9GvrDLkoqvJ0lyDobDteQZ7y4h2
T/F/Nn3jVHoEux6r0u6cfX6mJAKbMgPNfpBxO4t5HII8vIIlDxcJVLQPkbTuGbaM7uDUWVszjGpp
w7PNRD1rLGJGFm+p3wtNiiLenBqsxaoOzL1L2vuTKBlu0kbwGllrmKCr4q9PfZrSKr+G2iNl4cUu
6nd01AQzBWVlOx1nYgE2IJ2zAisnjwQazx+uyB9AObk0grcU6FcheMQV8SATe3KCk1ewQFrVmqtY
kRaFkjQYDsLJnOinVbVM/AbCx1UnzfzeQbIw5xvYwBuIe8F5UfZpCKTCb1XpnV1JPknM0HT+6Ixl
iNDI2Y1Dzu9wRIpQTG8XvBrEah7XLGlI3xHbeFAxGEAY+6VqHRvNpr03xkRpkn60LT0Qraet/GI5
zjhrSwjIof4SaoANbruLGrouLSqwGE60nA2nHN2BPJWeV7PkwnN3UQccLW/s/UQfhqqe+jZtVKiF
wVf7rOvw0PAPA1H3QzTcwYLzzmADORjdDNPGpdZyb/wlOUXBeleexVRouoCuAEfuNL33YwUlpIHm
YJLUsXCI7zaUIwp8eq82VKTUuIBc1QxMJC5hlZl2A8v9MBZih7G5r1rBCkrj9djHvOqonoQ8RbRI
dA3iXy+ya67pRIuBrXGp1oK5cEfynd7k6IvzKPe9uI+Y5ZwJjagjLPzcCLIe0TrBou+CvjOB7JUH
Fu0PZNqGONWwxbHEUKaznJyt9ZrKOdOUehF6wkcSp6aGRKPMikeDSM9OU0i03lrcUA8ZhNTqv+0X
/qzX1kTP+HRVqRB2mv8f1p+XsSxTJhV7eyqahamfce6hyR3HF/Xw7XUy++ef8uZABTlvYs+A7m6j
d/nUIZ1e03adMZcl1RM7mMRkqojhvGBS6Ojbcsk2XEBEI5G7Um8331Al81Ju0U1eL2+N6bnpTF16
FTddZbqKn9A15HPmPenba8N5Dat+7U4BVNrRjNt8+tPUMuPvxkcuIm8VSO0ZiOgURq8400BFF4s5
LpDnoasgLRN4sywt3u7wMa0iMMp5sMBQjLWP2uqeUJbXEK0X30vpLaOz0ySYM7W/dzBbPYePSlEj
mCW0wfS2krwSMxfTIQouLZo+TlezJwKTsDcOYxjFCLG7TDTU+8rWqD6j3yOMkKpN8WDAx5/bvQ7R
L99DszUKe/XNcYtWVp1j045+Rz9qLKfHQCpiBnBHvI6W1D5ZYxnHo5e5BMCG7hH5IWRgvCzVFJYT
CXYhUjBHjRh8+pxwYFg0RrPGB5j5Hn+5oclGj0IQycu7u7tMz4RjSDB8l3z99H4UPGEw/d3Q309D
A53JCQkCAeYuFZNUt0DVLYr7q5+0FE6fR1YDf97j1OedrLCkCwrKgrRmF82UR2U5v2fsVQmIACKj
BbWH+4pmrbJO9GLC4cwzCSi/+oZCgMx9AyXFrpzwibE7jTGWWddcOgVQCnR7ByUeMg+6Iiw9UANA
OUnbv+urzk48sGXJ2nuW5JL0PiD1z05RKwbwg670ZLx2kXVF90lj4IXXMhSZmmTPdLf52kJhjAi5
0mb86OQzqCMkVYCpckSfhTaA5WmKpusEPHK3wNsnaFhiabvDczNTeADfCUhcsm4i/5W+V2ySSdfi
OfSunU9wFz+4UVdoXuiyrq4uqeS9cjuBfesKv7+jeIEB/IpiprBEW9w6HiB+sd8S+behNPZFxvk5
CKuJFDlZOka2jReg//o/7xY0nijR7Lu6kUkXGErIUzirYKYKIpY/XxCm7MVN+/JzZ1gkKEDcn9bk
YgTqej88W9QyVoWFpniLgsvdswzXd3yxFFF/hRIFfdp4pfQHZVfn0NM6A45F+O2I99oG75qkK1t9
LfiBBm+/Ib8leD6G1Meipj7SKocI+xOwSSNQfKSO53MHkEO1QTcNjC9TQwcwjyNa943dcLdCaDvx
U242FJkLZxPKFmIrasaukgjou3/ivIZCxjr9S0S/bCrr7II/rxF5asOO/UznnDnSty/cNgq2n0o8
2CiLlyw1PURV07pwSLzO+Ao4kQKXjrxIr1t188lqWbrdq63SLnrlPJ0C7jAcT2OwYavyry65xBYO
j/3UeDQ1Of7iX4qUJxIRo7/UdRVLIlh0HbkfH+GCvqV1AIyhglECNhcsbpAqOJe8jqtBaWemtXrW
WW3KIN+3Fdz5OF16f/E181lYt8uSLOuPTxLJaY337ARV8ckcUq4XVqvjlq9pGpawF6FInPQgfG9k
EGIv5bDeEL2u6ka4iiTS8+egagT2QUzurl+Wvac+ZISjDU42qiq0Mn7PRL5OnKC6mp0EuMGqxhVo
4+o8HarScRiNOlhC3fUBDifRM0eiB61sBqfa/evqDpCA6SJHOnDtwMxknBltKzO6EkSsmnK7c5s9
bt/SlOZBJPwmKp73zKb1V1Kb/KpM2CANmQcJYD3vFMEGEvBwBc5RfLYJnl1uJnmXuiXAaR3zPNwQ
9YBTeBmTh8F43kuRNGFLjnXqVA2ZCneWpyD3IzS3HZkde9sIz7IBYil1inDpZjtto0NvqnsBR7BV
qxoSnrLJzX21Ds1nDYTDyi160ue8tVku30YSZvLNayPxCXLOiEKoDJW3rRQKTh1DbtSSxdbg0rsc
1U1YwEvuDa0niDKoR/330XvNCOobPL/HhhYDe+Un1+yf0jfrWcdcxdvAnwWcING/3p/uzVMDeSAt
v+lU8WJ7ijlqvbGPEONt9GpIZzMt9Xu9ZiwJuN0KGPEduNSZQSiE6j2LBuq1CqdNjR06bOy+9N7y
tQZJT3HVRBV+sQZx/oMjS0qXjwPKLEr8aAZc1AP6A3qrq6StlVJMAkdoeTqxpkSdf92bq3e9lDyZ
6H/f+DlYfjHGw+B+EVAZBsxglIUsZxo1zGcAi34kOmvsyVzyzALQ30oPMceg9HYbl97RUTxB/40J
NgU2rtLvT96q4orz1RB5JCbItSNRjMc1/We0SsJJ4VGVvwpyqSGp/2YPMIsqz5yR0s6Z/RB/22Ge
pXRQje/IqoBZrA905UQ0IIQfhwEBtov78UmY5KE+NcPmHesanjASVZetn+4ZOloL5nl/GUd+FVvn
XH930IxiBLqG9Z5+gSQR5JsRoqfabc9WGfpXe07Nqg/kKW9fnY3Ihy5qev6qUMKwxAaa4zGGJxOR
vMyXvh5Har3hF68mh5NBjaxBD7TdRJ36uzZHF7sOZRelHYooM7aXoaa2bJTnMvZWcqY5Il46Zpfk
LEw1Pbr4HSxVhp6/jO8YNugn+K5L14i7o4gHgN/fAzObMn5UDkaKi2xL7soSgjieEMfUvT9Z70Yt
PYkEBX1tgOWjPcytSWshnwwHf0i+M7tyZCmvF8dVOBNFfUrBzN+fIh0CyBo/PaQqUvr+KMY6OLt3
+268AzxckZV6FBUyQH0UtIq8RM5BssD0bz6DZ/taOK64ZT0h/Ggxz6qjPLTED56Y0bdaMz9gbvYN
TaK4gdpXMVFe1cLU7hn+Qg2zhAZVWKsZwcbj6WyX8V1reJjqQq9TEe3EpfwPlPEUnx45Bei95tAj
gAfEZshAHbadbQ10Lmxn75AosIIzN09Qx8qqrwVLZAKpLIOGmqX8lw0kQILecYExKGPrPH8bVcdK
HiLl+cmAzZ//6Tg9kuW9MUyiWrW52N65GnBTn44n2WWsKEBOj6QpAD2/PkZMPr5NeFWwD3rBsvlo
bCO+MYimJX3IYujuMvJc/1pQLHGRL8/RgzNFlf6V5DxI7aEzX5+dD+W55VkcXoX9SU5jVcn8jZa6
jh+p7j5cFqKI/73D4SYDu8v/PgyJCTlRYRCH9NAghVFBx/+fpUtNC6afljQ/aSZ+jkrQPuWMDyvt
ekx5bEnyyGZXKgdmqj0ICXZJLLKAaFVuZYOpfM/lmeg7tXQzyv0mjgp26NPcjYJ3f5y6RX/wU6aI
YLUgrvrQeyDVXuMTWVzRXWVn3KYo4PKH430+kJ3/xq/ERlV0bO9INOjM7QtdgkMZhNFTbnZ6iCKp
rIRg35t2mh0QRGvKBdICwedDy3bpnQ6mAZU1h+wOTXJ7JXPs2tHJjHi/ag2CNqw+9x+d43RfImzk
seEwdqstkMTo7oaffC14Whu5qUu0ETzD3u+f+AUv7YyKuRbPrAkXMhX7sAC3xi6N9uISw/QK/XQl
KqV3CPqNCftV4sqOIWcwqzmB57rIUBqk/ojC31EfLGBA/MU3XvIklhZZMyTnhstb5h3EatVaiz0u
YTLRnRDn4A5wJ162m3sK+oz10TL/qMb7BD/D1H2CYtoy8WQO3rg8nz7Lo1k3EtRPN7PZvbp/6MTa
kChSWGRiWektKPG8M9Gj4h25NABbBLqg1VDA8CTL+gPKebfuTrZTotcdEM6WPbw4LwTlvOO2/Hjh
jwJhacQHyLWwZ98DZAGaeSvbeS12UmEGAXips5zq+eVEYisEkEkQyP+Qp0ayBQDLWskFw/pi5p1H
elG+z88ME2g9+8ZRfr/hcReFbMeG7ynIgAEm6nfi1bm+oY/fklIDCQUzC6X57MLn01J0lR3ZxvgN
Dz9IDWcG8qWb1wLW+H023d8oTe5v131+abBSPZrTqrE7on8qDC0FKOWzvChtUlup3XZ7zTBM8CJl
MqVi1YuTLLiOy//SINPoVMNE9oTusFhvS1iNlFOIRm8XbruYEmOCVvEZQCdYkePvGrdl1S1fyPb4
Kbf2sT+4VT0dAk7gbqILAJHANYCAgqA54AosdL6Y+CSf0g965PPhuXpJg6I6RcC4I46cCUFFlb/a
7RMFXNyY9oqURp2+XLCeN/Zgl6cATWM3Gi/c0nksLq4uuXjjw42uA7Mi2FTVvKcVPFyyFC0kUA4d
sDw8Z+oJ4A8EiU6mS0RabKTzDRsI9WCjwk8wTi17Ci7GeuChe96pdohMWwVO8TYMMFmGoZ8LCz45
3SI03kIZiOY4T/XKfh2EdDBrQQDFAyMgAFbibp/sNHj+MgN1+kyZztQjyEYoU8lJvn3eT6kFU2+B
tEZbZ/r0yKNVX0xPOYgBcUOxPkfTXjMbgSm0p7ec7/Oh0gxbpU+TFXQv6R7GfYKBcYKyF4BkBFWl
8EeOi25dzf7w9ug1H1QaRGQh6pbFHx8AEPagvnbUWj/ftmJTlWoFkXbPj4U0/f5GQReyj+2oVjrq
idAX8Dj+qjUk3Wn4c1gLt1z/XDrF9fGN4pnPQImXDV1dm8WgXvRRinGA736N/E6NY6sbSHg972AQ
35qFc+dsUl/lFcAx43157xdU2MsN9xpEGN4/AIC3TwFNi91AlrOc1iQ5rPR556Q3rfQwZDtOjcAi
W5MszlNFIChD9Q2jUqMv7n7vrwcZri1gGO6S13bfOQ3yrudPoj1MHBrC+8jWWQzA7FsfG9fV+Zr9
UKD2H9M0YnJhJmKPadLfK/XslM+pdABs5BLskedLV9cGlSJfRQlEMViNYM3kHp8axPlyL2o4HgkV
JnnqTiobzfKsEUuDS13l16fNs3LZBhYarmao41QXSLPDTzZoSX+ej5ZKzNYEpVd4+5FzMjfW9nlv
6SUca3n9jMok210FxWm6UCw+xz8kZ+GBXJMf1L2pGO9/ql/SzeNY6hRsGs8NYO2s8Mm3XAzt80s/
XHkdpuwpHZR/XINDh11AXAQOKv6C62O0vDHhwEXehFEXlFfKNRihu1ttcu10ZzSO1YE/+TJa6pJN
Glh2G5p/eAD91Dq1n8GVv922OH/3Z5tf9dQN7rbDu6r7WVo6Y6WfXuPw0yTZdfH3Ag36THyDnkAa
psBBmnjkkc9W1xeKKhYsWvYJ0jrVwpNnUlUPHlp6I4pdsqd4HMXOuVXmd4pFBjdvlF8Hbs6PHEiY
Jtpui53DXTP426Mw2bZUA2+P3JFAOf/j2XM037gJg4Mttb8veLhR3dOurKYUyO5ukWVHhA224PML
mpwY2ZReZekG5edEtOalvWW7BUD1AlI0O4Yq4zRJ9hpQWC7U55SDL59CtKDBen4KTnO/hahcR+kv
ASPChEvacRXypPY2hacxJCo5B/1akKdMYPe1egS37MJ0TPQ1u4fcW9ElSz2yOdYBFLKqLoMNBnVn
PTLrpqZXyl9KTkDP24THlTuOar5qdgPN8OubQ9SG+Wav+BlPYh/NSV0K1S2uzLGewDdnDzVbKTpy
18mYNbLXH5q0PdSLWsa5qEXMKwe2lvt3sGVH67M3ZEmI2lo04fQhiiccoE6qTBor+BivYqHiTchP
L45PG0CRK4xFmEdjtUEy1pNtIn0rXk6eqr2H5xxj0U0ahFqN5XxeeBceLZtxfRFF9dW1JZB8uBtO
0fGVcjZ3ob0caNKRBW/VyqLhbDf5EsnoCdEPeixc+Ba/tLUBGIpM4qUaYPjOGpqvRgE8wu1Jaivh
UjeG/Py3TLusriqQs5AVsXZYbDXSZM7CBNX00iQKEPKo1eO0XCakvRvXd9VkfPS3GSSAcUY3Fzxs
B1Ze5jVxRvgwmvwMQe+ulKW+ZkZwrtDzs+xQ23u9wgnJIVvwNxBrR9rfoi0v7wUEtuJr3t4Ik5Xk
Wi92bNchL/NbdwKXcw6lmFRj1aLZVdXeCuRqDEuNp+qkM5sgaZ6NTOTGt45D+qVTbv0emW0tcvAg
9mQYE958TpThzx87jzLP7yaaDVRWvFjZZajGU+yaKkb0pNRP4zr9h3oOCd5j8hPRdfdGuJ1n8eu5
/w1F9o0yRpp3WFFcnxJsOsJONrxgdaPz9j7tGbnFdShwcNl6HP5YBIutjD3jX4e7T4YHv7tqKhm0
5Q7PpF2hsl0S4Rk6mRFYBpLIq30/h1S25LFphjA+MK661+SD+vjo2ZewSSBoKzeglNBl5ZPvrFMJ
Bk5B3hns+3bXKQfKu144pI/C8lnp2zyG4pVFvD+nhiAMCyHxzlka3UN/ag1e7DDFXajI6Ovkg+K5
JqhbjgLZ+1ksXCRW5lZWsFBASsS86PvtaruKvOAl8hACjmesV80gdrgV9Rd/dKDEI0fAdQa/XufO
/7NF/dH42UvJtnbGZBBgk/Uh6LggDOMz62x7rU8CWieoymDAAMjPA+UHz5lM7ZpPsuibst/UHyYg
mZ5CqTWj9oJR6B6HQjbgz7WfX9JX7PIZYi38y0xkcAO7OrBfbX5g+rq4880QDagV96+Eoo262K/D
eo4BedlnuKocNpmeG+z6i4pjpnLv2o4hAfEfLkdB9X1TzKXRMCr8doBsCtGadU1sUUeAWCuC8XtI
+Dj20E3FbJyAikZruk97uCiolFJU0DGxc1FXZpF9ssgF9mVcK9EaM9qa6IxAF0RjWc52sPRH4z8B
yK8+8fixsXacZ9kY96MnuauMtylR5ix6TDFNDxEhfe87S3k3FumvTaGjey3d9hVt5jQk0r5in0P6
LDTpK+jvWP6vjxTH7NSamEZ45ZyXqzQAl+QJomj//FGsrrWtqVQzwhvvaC9RAKFgQEXDUG/gPnC7
UjjfAf9ub2goEg34aE2NDzzDprvIXBuTyuf8kCFWE9+lCHDNj8di7PI3O5zhrNCcyRA+WohnAtxx
o245DK4Ul33sEoQ0l59KVfCJ6sB3oX5mB1RoyERmM/fhMAlFuE1agE7VL0OKAQWz0eOLVzNZsuAv
x0OY9GpZmk0RDpyF20KZuLgAExyg6bUpz8G8Hbg63yVJgFCW2cwJtzv37Aj9HfC0aSXhn5tuwb8U
F1swE0kfs/H9ekk8TMy3Nyt+dhZqoHXY+a/mk6hCAf47gqOk67Inr9DmNxDu7sxMFlYWI+oIGZoy
avQizVYJlFD/JzEIRhEqdntxnqtdLIGhQ0qmeuiD+5KbnTJKzQN2LcROqxq47oeHZ0igzv1Z++/7
/+dEqUU3hCudED3OaQCrIZbQudvrPB1aYXov5MMcN2zm9Z8hCRK+YkSOlj9e9Ota9aJh5ESIkDbR
Fwl/w+ZWxt+bhiKQwVoz1/f8ilePeEYHAvqoFV8KWqGRVogDC20Om4TNcYjbjIND5UaYrmB8vJi2
gNP87xfSO3zO+6eu0wwItm5yxlPXoVkTxXwrgqx5plHRr89u/hJYXpJ+D5iuipSoyZRhsuh5rdxS
Fa7wiEYGuAdQyO6wmWyWMa2l8O7BeSiuQvVViGGVf4r9RKsKabgrQQFBXOsiXtE/TkZNtJdbHKsm
1SOLCfoC23XbUfBQ1EaRmB1RWsNCw6M+uCEeBgTc0vI8ttj2gpS8kdW6/SEkJtYAsVh9qtPJ4JBh
ztXyvt4lKz+qNu1jQwkGXM5iFl6owNgJ6bpr1jbq6zN+zSQOOLXT+DHYr2GJ2MWzhpPVOEZTnUlw
QQA55zgfO5a+bk+nMW3/aOsNIs5aAxJ9WwZ0APGEiS6C7W7ek11AtWlgMu2HZo8flzdcwulzTYaT
7Ce0U3L9MXWwbODnWcEdZumOZ8+c1ST2lJ0Or0ow6Q3Rcg9tE0eP1gaEnCwE9OwYzq8Vc47c3o46
I2b4eAG4+KIjcH0MlRkjRibdxSJotkHolJ7fbZ74miBG61JwyEmgLfTy7qEE3t8WxI+pXaBtB8/4
0yXlfJtBBP75RQzHybSDt9KNzI/b8Gcmu6DhIYlJV2P5zw9md+5mVKmI9+uV/c0RQB6kJpeLiEjn
ldNSieZXZKZqJtLX2PlVRMzB76aP8p/A90jfYhRVVQkslxh/G8vyeTr/WR4ReKz8rnddd7NQyIhT
aqZeAtMjBKakNSemmQKRv9KtQJUmTlDXa6wp4+///qKVrP7n8JFO8uLM45Xg592g/LIyYrXlodSO
q2DonAdGrcoyR78+epY5fupukElk8lZlhByhQMjucpteBmi0UYJUugWvjjTpeSdOitvvYXg2kCoP
VewHUDyisDO8fKwALMyM48YG82JXfDqRaDAG7Zg2ABkZPSsQlTHyQ2QN/luy+lQxl55sQFL6hOxh
3wDeE3MZ7iKSXTWkHSOLsaf3ZBLy+ae5pEFmyAZStEiabV6J+9NlDm3jmQKM4+usDHA8CkNUy5Fb
jfrw6YeMdZPHNcNz8tOOlW1J6uV86pYnYUwvYU2Q50TmNtzjCYLulxaALJE2wjlKKfZcWSiQach5
DCCy/V4E7LIB6TZGvTsXAOCfVpzGT3wfGao61qw2Pb3L/J1yCVrMNnDkRR7X/LD6HO+/PiNXX4m4
wBSqG0FvFLpPXHBHAY0/43OBRzrk8+9BIxdSLUaWMTlOI3QA3RYEhrwlj1t9e2mXSzFeN5tW25nl
eqTOB1iusxJDsnwjhVAz0c2o9wAK4RCG+ZNA1J6dApG9lbhs43CGlwG5HrNpKQ71xynIWKhf7ypt
AxLXsvLmAAPPtwpyBo+J7tks0OK5rYGS8wpggQ0bUcMNHdzwgwAek1wqdlBiEDU3ke8Qi1kRfz5c
9vGxULVIdc3IjAhuzsgD1K95ww99UiPHzOo+2B+XTHDl6WEyUN1FXXzkG/QZGwYhR8z6bVdSSHER
A5usaIsfMPbUW16tkeKB2C8N3gxFNdT/2nRFsCxCPA1buQeHbLCmZqYmQKVc6a2NbrH1MoWlewjm
6rqpqnutoqETX++ZWNsXKE2ugl8dCGIAtjKtVOjh6PuyOdGMh77UMt+gN4b7gdnZL7gZvoVK/BsI
jVgldAt69EUfYOUvLnFX5IoTt28/Ns+/aQsltGaT8UQ1mVA8hB1GuNPlyMtLaoaG4Xcsmn1YGB6p
eF22E2wf36MZHV1BrtW7FmCPdFjm5QLdUn+hvhCAfgrTrQN0LRuqwoiFVd68kQJA3g2ktKdH1ZzB
KXoBTY1nQmHv7AoamYGhxFQHbtfK7cHja7HBp77gz9zwi/9laWKTaOU8D1KKwaMVKv6lAhme+dqo
lDv5ZJQn379ukepVjOvzsMntfYPT5lFd0pIPqL3OX+OgZJAcjJ9vSHu3w/d/o1nWHNJllrV2fnd4
mCAq4hzrA5uNkBFgZIjGs2W3q0NBDuCkKXFA+yMf++DYi9ZWUZ31dwQYmRisuvGwUET8qnDfWW2F
3UlibnqbSnYTTxvG/gLpCntkbP0Qh+ToJ2LjLwBJuCZ32JV9xB7T4UKgmqua2R1qldtUrljJpNHf
TpIYzAFwR1fACMZR32hUc3KMsdfzRrv0f3lKAk6VboaOxV3XrZVvQCWfpZJApvNsV/Ocd0G8ulAT
I25uw3Q0xEAGh3nY4JG950sHs6vg6osHAvmtN5eLgK2qWSfwupuMH04HlGZKZ2aqe3XcmzA0H+JQ
f7yCujxGGUlMMSQtj+1bZkPmJgPD+llwtB0xPVv0cT0vcdNMw6D1ZYRQrMm7S0AjkcyjqKiPEk1a
BmFdAa2pgckRwRrWW41e8IhBTN++0p9ZEFk1RLxm+tNHgWxHt0w4xGwvfkjOFI2SfhF4zXutRWuh
/+zquwyAF/uwImMumd8PXeoomPGQXQxQFbKp3BVBm+3nm5U15xDa194GKQ9FXwSNve0vqP1sn8JW
yVi4ExLTrvHFn7TECum3HIbz+wHfl0r4I3KWIDPh6emEXQyNiWTjVf4GPzIi8OdYl3wVz03vYuzq
zmhWB0Hc4PGxaX6CPCRoKwWJOeOjHRzF+4OhtE8s+SvnUJzxRwmK0/BTo3vFFqaYSTtRXdSTB9MR
aMH/3IAGXb9pMxZZQ40/qGnnz9f13+D4/7ohBbE0pnI7oGZxLjkp8xjQfqIsIN4+boVHlEtXA71F
e0KQaRgVqvdYrLXO2EzobwoHoKK08FNtSaPQkjqlgD6sWWzA3x1PVjUOw8yWCUALK6PQ87FDV8u7
iM4/1KEw2dzEsicwXa7wR9CdNz+FJTKZjB0XJT4Bl3zVXGuQtnBgn8UpHi8FisJ4AZ4+SjnCIOfz
3rukaIIs9u4zLRLGQjcm8Ob7kfkBhqL6XF0lJNPN90ESQbJKaPje18ayGGTQgzENu1iC0GFV3lD6
r+2Z4nZR1LnrYNlVlxKCZD2mxrAljH2s89Z+bsNrMGZBCgJRwAh0zfCoDpqR1XLig0BUbtfEpmSY
FjFOahLDJPGGXm7QKCGW8cWWmSOF8nBD7bPgA9ULO57fAQyVHXoJd0+HuP4twuXc1CI2V5dVpTOV
PB9cw/ayJeDB0reFWnx3EPkkCDsyE3KJ+YVPGGjizConBj7smYmsUQpYsfS0UI4zlSz4QYzlQYvH
uVdF9LL64c6+XpXbuHlpBaa9UVORMjZ2FWHAibz5istEjMjCWEZ5Ryt22d12L0tb25ArKpLw6gU3
HDGAF2VY+9YV28SOnLnjopTMXJyUzVlLJwsm9p5JqxVYDRikn0x7W1pZpZIYrBjXNoAGHJyVN7Tv
Akhk+UM6a8QQuESpXl0XTNcqe20FbVuU4fTsBNu/L/Jz01YjP6K9w7M8/0YoTaUfmQc3OQgUl48+
p02OGCv7E2VLSEaQ8xD7CyEztUgyL8QRdsF+S3y8eImO7Ci6hysLW/hqJW6MSWxqptMst3zpOsjl
cvfai/+9CfiUL0Ew5NRl+TIHb8w30+t41/ZTcFX5JJzpmkj98Ygs7LoaxMoUhRemoKpstN4XG404
rs0idUonubq6n1aJKncN5kc+0vKKc4/ET1KhXnv8lxfQ5b67m1IDFpPwKmoBc7doE7zwRggRn6rl
lhRWWam2WCopZeaQ80K4dqQayjiikFyX/Wqf+7MJB71eLK4IaJXtGc3zeZuOJ816CtQlpt3FFgOW
FXhBW+mOyEcHk7xz7g/nwgXuq2IK2BbluJaJi/gpBJ93ziOoJPwE2rJUzCe+VgXZALXRaDR8/eQ9
zM70U/YJWmM/M62p/bHykiEV5BGtvuyprH5NXZm7dZIG4F6BU7UP/CbhN/qtLOpzVwaEpoOv6Pq7
fDFTNhUnRJ6xk+dFDIN1zhajO9hePwkondPGjt38v7Jc3OUqE3zALB2/kqka27UHIqjMwJ6N4I7M
I/pP8FYNMSWUQ+dHZHo9DlHzrbs6QEFaRyK6zgOhzCjQUz1RaA8VNzTx0972mfG5sPYQAUC2Ps/B
2f+PcS42Jh1QfKfIMN78S2/h9VmzjVI79H4cohsaExCaI8ZuuTuFZuvhky5D1Ags1XURZPymoG4z
93oq35g3Baz2crZVV/vOXkIXcwpA8QDZgdpuur3LyyVDW35Qx62Kjnz+piDjRTkR8HNNhrD8yl9q
q0qHuWLz8gvprLzcyrGfI+f+woqqaVO8xiEZ2qGjwsIE1cbEugfwuP84IYHRYkU25k9a6TyZCZ/A
A8whKIrcBNQvv+7rgi+3axRBJIFyaZT8E6fW4cT+J4sB+Yx2eDOGlHCz7xwUd4rT7OnfJFbnuUAY
ZzN2ZL42qhkNsFFxRIwJzQasJBAZhYZbO9NwpnO0/SJqtYnq7QHVLNFEKcVFv5RVE6Q4uLHvPRRO
ijD2ptP6WRN8M0o+u5DHeXg0dx+3B+fltlriJ0o3HigJQzuLe8yK+Mby1BfUJ2X49HoU8foUzryl
V3Mvbo37g2DYVzP+3Pgb19KIS6Pu0a4uZlD4QouWGREWNElfHw64OFWStUcAkczzuWK+KTaQdJpd
zZzuhvyEZAPnrWyvwqUMJXy79betToevxr5oQ71gY0nLn+/4Y6PGKWNEFtawoMon/TaYpE6GfucB
EqzC5hFMwpYEEOo4Xocxd4qJUQvtCBzrF3PeUIMEiWhOeBUo1hOvYfRqkFy4OzTPTKanqaWAsPET
p5gWhkJwYWUXzem5EZ7Akfeu8GNJGLcjYWIeyz/z1IG1CTgRslT4OUFejWvK8GHVBV9aTSt1r9fm
5OyMTuusQjviYM8fxyROofZzWq2UBqepSSu8usb5qB9x0XlRFZfAWgj8lEUMTl+QBA888QKtv+L8
SM2qRcD56XX7rdIbdS0Gfv2OSEjildLM29PKOJg1fTDFrqNlS5tvB8/BI5r/cOOrwEmMFC6ab0h/
ZDTo56cmjr/SRxQcX1yL3lX7WILrKAqkoVrq7qQZ4Bpda9rKH9DzXEo2MZGSPgBxBqu49yfOqI/b
jguakyj/uzvubhPSFqF4CAnB3prM2XX7ZsUSOcz+KUsxbuhFSh26P41Gc56xlLWfON9rPnQ1FU1j
cGybqC3y6Yg5fNX5v/8k8jhkne46b3PNNPp1Zl6f3/m7GlQTcQ5dTkwynLAnDvCafrhVK7y1Rfxn
bOJ04DS87omOJjEgRpjmhKSeka3/+XxKxWcuxGd6HvQbFLsK5/h27FAs7UspBrbfqzjCj1Fk2GMN
lAs+7v25Is3LI4P+103lYMuryL9ORKZXKr2yqG0wcgBkm91VK/IXwzSvaurtQUv34pgg0ks00nV/
CT0xqtOSotqV75lnQjrACPkiDPUWYPMPKAlzhYu3QjW42ElLxLFlvb7NxnrgWDKV2LJL6hHTptw3
1Q4JldymwbfSIdTm6yfFibxGfV0oyV63YehShWwyYSQYtY/8+1OgJhOtHFU7bRPDVspsEz22wRn/
k6U7Xq7eBWRfZL3939rGvV4shuENAoZ0teY/JzMwkDIfbMZUKKVbqR70BndcxHONKLhfCIGCEjP8
JDLnkjO+pTwSXCNHiCrddeUwYfWlIY0eClTIAhFRXM5jcD3Ok7BL3cTBDv8phlpyp64wMoif4EES
c2YwMAGCjfej6M3cXRHnEXNqIPepuQb2ehIuMCTa7jfrk9H6KY9FInqk7FgvEzAN+2k+I0Y+jcIS
rvFVAF7eDCPqLXutmDYckY9rq7SnqErD0c2pT2dDvfzSCrFdX7Z2pQpQZktTyN+WvRociITsHW5H
TiztSdHcvIJ3xMjYQiU/843v2RRv1Sj7eOuzE1V/Hr2qoBLUQVOr1Vj9XDVzLRJo1se+fQX8Eg3M
lcMUsuz/t5Oehz0GxCHdplPaaTA7hRrP6ulPsJI2YTbAASCCDPF3rufTn/nAu9+OVnTJ5U7ns9R0
zd675YmQZIrZCw/F72xcBSngrIKonbrm6DgNjCFzTj1P1ABpvfqy3acwzWls+pIvR0YISMjNZ1ze
75/AEW2HXvWGD/kwvW2Kgw0P4NL74AfqX0S8fhpYXwzkj8F+ne3IqXHe9yr0iDRJOnewMK2kmQLT
diha4yGa1uXhooMTEUSoFiXheyD5bvW/wPFSgksRGuwvlsNd/YdnQBBxTsj+/y1/KQp+4NHhgeQI
B4oDZCWVrnpvOPag+QrHz/RKq8X6EskX0Iwn9fNFpt+K1JwcAnZkBdM+aqgWE55dLVjDo1OVl6ot
2uGpn/lEi/AujLNhL1L1GHYeeGY2g4zZeVhLnPRK3iEwQas1QkXW/bwWxdlrpM0829is1Blme1LV
uVnbZqHTTyKnXUf7yVWakAez8D70Nof82oOgdW/j4M5t/NxK/I3xQ2WOeWHFdVc17Zi8SW7u9U7h
9EcifwPPOTSfPwzGuhIi3GKHXm69a1Taf4imvdGuNZXw9ndqCbGJ1fAjjNOjwNMTlrvwAzB7A18J
WaW4raPuMYGQ0wvLTsyxksCcMptkC1zyi3mbnEOCzQ1pSmkQtLSDoaAxBPagy9YTkHdnIIOOuvBa
d8a8t0qFPl4LMjW7Q0ETg0KU0iz0J4iivNfrw5yKp9jvA31i7mys3NKWJ/pgzvOcBI30sFKQZo3X
OWupzKt7E055YcrKmoxdW5OW5Vk22RwXgydeIWknrP2ko6kV0Xs7d6aAbvK52458OPSRn9GZ6w73
jfnQzrpwLpxqhNgA98fPH5Cad+wASYo/x9f5vQ/6Q1jVfZoQx0vV6goCrPvCwIcYvFAR0eq9ewdh
2ddMRDvRYPxvnTClJOxK42OEMOXLoH1FMrmebCU10XP64FeA8h4dyoyqdnor5sZ+JFFx+N78/eu5
r91nYUEov9fPV+Nn0KLoPlNIag3e0VPZM2sSsQJHIMG+tu4rT6c49w1Aa3Nm9D07IHgHiTylK/9d
6MyA4az5dRFNxTXHupYqKN0/jvTghqO2hYhUzWuhtjOp/fLEcC3969Aae+JrP2b0K5OUk/W/BRvU
ST6F7QqmjuxMigbbd1jNqbAUcT/Q+VsaJZRVTu14RC2Huyijrw/1Bw5itYr6AJmtfvucW9pEDAvy
9GPvbJ36MDi9PNkYXyn0ljAMECWPxib4dlfSA/tutdKlvJiYL6+8kh5YptIAXlGCJXPMhUjJt4VV
ZfgAnzKB27g4rtI8f4mhKGrgvbS+lpo0vezGEzKJsrIn84ifvNHersMzthwsPjdDipmdSjQbIBaM
MTkKqe66XC+vA8GNB443k35nJotY4CH/cWl+BkY5IPXz5KuAPn8xfh47TZUiiRpAequhRiLw6wbk
yPt+gCep49PoMUCnbOpCfwT7nAEgdgdqVLKkaebz0jBNTJhV4OJoPJ3slOiPCN7cxBqhBrm7ZrxQ
Bbgyi8avXSllj5CYzloveKOOneEGTQiMOtNKBtJEx7smg1wPjJhBvEG43+JvwFTvvIW3NOQWbYRV
/QQAvXKG8+/OXu30FNQGbfNxzpNwTkWN9cGJQK04ShkaDVhfqU0X2YbThi5WnN1UjhVAPv7yu6NI
pmqfZGUs4iIc3tvt/AN1sv7UxLkW9KOWSrXRTzkhTuamIlTYwyno+5yBUmpA7vDpsM0dpXBAdC5t
BLAefG0Y/QLVFVT811snr6OkIuu5Dil3kEnwGcrcYBtd0wM5GuNBlFx6qZprfwkM6NbGBkUxyC1E
gXa8/vt0ncFLxuTZ8+4HRn8LhttyFqUOQswUIFzrkgYgssLTOqpDief61Jg345ODF6USxFSlCJaS
W0ellgd+zI6rrdOhUsXQxx22X2JtxPkNf0gRcGC7lmU/B0OkGtD0OdmPccI2MfLR2PxlTKLFH/6W
t9mmPqAjlyzm1ZuAzgp5dQ0xaQh2/ZjMTyYH9ENHpfT41yNeNO5eKm55YbKzh/cPP/YV0I2NrQ16
Wo54KYfHOvUft9cUUtZSZP7IHzAzH8JCrPUexcaF6uIcQAGW0xh6H89hZB4fvt8ipGFvOr3fd7Pq
dbzgT23AByl2Gl/t0mXVgsVy1Fjub3YrXZkm1GeDrVu/wTCbE0T6HL0I7O2/H8mZUYwTca1FWoKV
1TgglHklM+B2CZ44ufABzhqhiPk4BhlO+At/tP+eRhoOXPPhjMXCgq99iBHnbQAnxpljlSFHzJl8
3zoqw5DrekymC00e3v6BHqaSX+xpSbxs0Jw4npMaxdjEzuINafp65wGnCZLVIld7ycwGDh1FyQGB
CVqzYcUKTXEPS6VI1c/6PchqJZl8lc8Oxy32mXARQuO30aIrI5O9TeAWlQwSleTP/fcpaEIK4xJZ
G+oW5sYM6FZDrlbf9D4Wkf1au4ceoaDDcc/QRV1xyotnmX0QYP2lwHwQDW6mMHziY6K0+e2EBK1J
cXWMhs9H6njb43X3KSp8bNXsfxUGQEbbGMa40Tekynb1L0Ss9OQV0C01PY9jGJMoGisSyz9WBxE0
3Ye9QP5LD+tymp08GxLMaViHoLKI//1O0Un58o3P9TfAm8F+3cMLhz3O2Qmoy/D9dHZyyU3Vm9l7
jLCehpHOutl8i/DjKK9DfSHTqenm77Wx81tx+eUB++ue8EHCxPr7R+3AjqiSyk/GjUfbDiPVjytB
6n86WSeK0YHouTaeOSEklx1Hnm18+3VHXf9GNI77qF0hk1+WHnhB/3PVNmUHEj+HpSMkjXaYXAR/
6nSttDuDLGuw2gc/QXjRvbyxMcth77uvf3gpT6C7/H2avBpgZ45Ecrwzs4aSRRl+PXxDBajhkzte
48hN5dT0y0lP9uU/zSK9325Dj8qdJAMY0htKZswOWFucvEjZXTJaVwFdISoEITLZttMldcSvV1F4
J2v6j4iUnqVVfYAVVMClNipoU6Rw6Ebqk1n2L5iz2r4bJBIvCFNQZRh/ZLOcwxY3dNxmrXnJiw2a
YxRVyWJomTllvnsoBqX5rwkQ7FDTAxqOc0oRS24SYNz8abvgB30bsanxdBNoOl7e4wCFJ3omZpUp
Cu6SarYHOA1qf5jlakyGMCamuoJ85IFe2LZll3wkVQUtJuUxtQRnYcvmfQQ6Vz9495YQ1IdOCGn/
qCJ/Pt3ZOudh9vYUe5+c5dbGLXUg59GRCKXCyhVFLlNz8qPBoqzhN5Ch6f01WKGWiYMPYgO1jSjX
z/naav6TA+5oKq6wZmgA8ukLDJ7ciiyYuq13NS/LdLz5U67iTyHz0Fx4LNxXtjeLdDfXBFApkL6m
D1Q9tg5KC2Ldv3tv+r+51JDYz3ARvlIOKB1l4qNcJGDtT33piZXve9x77YcwVfGMaKyMJvc2cbvB
kHbfzaneeT/FMvoPijxDTx5IqL8VtrGFUmFengkddecvty2HmA6tUZ2HLKvCOLUd/+xAi1zViXbp
PeBD5yXI1F8ODSMgW9NetrpdyBupnmw54hpui658YK/pedsmGdKPTVfvaSgpXF9r7WkFlKTuZMFf
C8iHVjrTqkFZORrbrJ2tDMytfV9ruTC8Hvzj6E1+yislddOett5jtfiaVh7FBNp5LZeKoCS39Qge
3dS8UGa+aqXl5l1eOu65a4FqIoWRsMbs2OXkG0VKtz/nhuJr2DFL6rqZcbaN8W5K0+hQdurCxif9
MwWi5ZUkg2N68nWkgcdoz26dKJXXYTHw42Si0Q/FCA+Rf4FRnXgimIAzjnbaXO0KmQzvT7SianF7
VWg4ViXrCZflanaWB81MHrt3xJh5izcFSEupuen8x6StKQRtr4i+qo55aPfw6POW0fJCA1capCVl
QJ1T9pDywNmFd14g1TskO+WGhiowg7PRNgcoeuQdjKT8tOnf5sEosmJHiD/V79EMhTWNE+ZbZYPB
5vjUPEYi9sjgwFt5YZ8T8te28Ad0GrNsptU1XUn8xo5sOzx5oZbaH7xKhDditR0vbJ4DuP2qcDfm
BaBJpPUePsBw8t3T+HEoJT2DrxfSTCbcPXwNisDHQzTvZWATNPNq6yjJM4c7PB/MgYZveU6YSoKz
Xi3VBneIQBzw82iVfpilV4EQ3a4qsMa3e6qPHDPTiXAn0ZWMdXIH5OxSxsddPnKBeu6mF+cOngwI
NJn8K9eYgxsDrKbn0du28F+Nkxo2H2goaUCZH91UCYTzm2CaIPBjoUsYEInwo3AikePbbHceAlfm
cxlItClJ+R98pjau2lUdhpFGGSuxrzQ08tYNfHiO1YJQ04dbVo/t5OyVx51EIETkqIBbnUkKOxRc
oMQmjyv66SIi0kt6bTwV00Zdjg0LVjLBFYF+fr/6LYlHFZWfuAqQl7Pr64/aAF2BqME9qYUpHP5m
lkI7hGFCZOuHR3LC8X5EFJgh8GRXYfQkCRemqd2O6YHwi2COS3SCJnr12rKhf+cGsBGF+lFNByXo
OootLkLNapxVePJV5rEBnNLGkL9ht5KGQgdnmZjCklD9mFACYsG+8eQ/Bxa9sAYj69ywm7pjGaOr
GmyJwq8RjCcn7uNF62dqZBJj+TXl959SulB66oy6zDlxlYSxHZ2l2gej66e4n3JEtP/9wnsgTEeU
3PgCPsHPMAsL/Nk5WQAV+UZLCPc6CVs8W+Wo8Vqkf1gPkbfKci2HYImYosjoa1SnjrvUjDGhwcko
fLttlnRuwKShD3I2+DTM5pijiJIug/+cgkHE8mhGqXccp04i3vXOu229BqlbKt9ttLz25H3kjvQ1
wai8BJdQ4kIrsH9Ou4D48ffcwUQD2nCDfDgKRCxBw21HH7qq/V9Jp5T+KuIoIOQw+v56IcJxgpiZ
wgzowvGYCPE1eWJmItwmVjyx2K8/zKGqauTg93/g11aUeN+F7f3UO8tYZC6DTmR8nlVHG7S9n3bV
Fjz0t2acRVDVqDkHHe5vgTTbjD1gkq29RKKrTFVg7OF4nrr/2ecymIuXZa68ahGZFj8ZHdfLf8XG
L6jkx5QyisjdiZW+yCpOiBKEyvk6FKCmm+bM9Z2T73PpEQn1CLpT8U+WJOuUOQN3mIt7w261cOwj
7ZEPvpFnSzSE6Bpa2VN6k4qPEN13EzeReQffLk7WQOBSi2dKOc9KdfvwZUO0Pr0sTmh/wsuxFty/
IKYWxGJImbP2lbeBdcJ1oV5vW5dssE48PrY4/lYK8GWA3gmGfOvPgsaiaEbP7dIR9UK3gV5sGUv+
X3NMch4m23k+jbgZ8mxg/XJFMmMbgp5Xeb7SeWEMwTIKxyKvTcy6Ib4HMutPS+oHZ8S3ZyCk7OoX
B/dgqj/39Ey+fDo35cEiGupi5huiNoWJ4WpXIQsVjbi/3+0hY/Mm7QkVzjwSCkU+GR9MVSn6+qar
vbjxkdXfv+Q0WoqirYpklKMvtV+twTszqRKwix3Gl4SsUhPi+TWOKJXtfEOTQxHTgPAuM81DjpDO
sWb+kDeajygVLP+2ChUjf31hcToOKuTNP5Gd+yAFYFp6iTrychtJyN4LJigk77Sc/Oq9VSCKmiRq
uP6lw7tGZTUaxC0Fk6ovZ6I04od2+vt3w6Ey+NjCGsm4SyhD+R80E839Q77031W9DqaollefFyk/
RjAE3xmuEQk8fKE6pD6CVRHhI4buu9MEaENNjXqxmIhg9WVIAn9+dIw5JgCgQB/7u8a82gO3aM1O
15YHgytw8VUcrjQLm7t3Yr2QZltWPVGQ/wkFv7aVRO5v8OMq6jZ0UM9geS+88zGg2GR2V9Qniyj0
2c3WrwLeE0aTxdecxht02azzynssnwcVWFRLh2qMUAYfWw9bdS/2tUNRGyLKXOEHiQD0zR/eVodX
GSaq4MFHJ8zBwNwEF5pcozki2f2np5G3aYfRL8/oWzwqOOZusn+DWG+B6rvY4flbmj9gMN/8KE61
KvLyVYq7nKAewugpKC0VmqRO6PeLH7lEkfMn2QCAqj0U1kPpdFT862UskmfD84VSR+f/0l1WI4c+
0cuLifpT0/dk8KEGK/J2rBR+JJEB0mgpRyF8jXD+kCQFd11jgiwmA4Cd9Ivt+0CJShkUH7FfFHGi
UaQSbGkUyUDOr0ol7Y47yxSkG0nUcHd2meymNkMViU1wX75But1lZ9hQjajyifJPeruat7i8lUyT
CXkw8kCcI0nMVgHMdIU9i6hxw7zZ9qwjmfqvZChT9IDilFu9xXGrSjhY+YFZj+CJtCeBDm80K/o4
nuVKrcOFlFzNNVt6tUZKDkkarPmQhsIkR6YFnSVneP3h+0z2W2qHlbFXEcbp62Gpb1zbD/DaEseH
5X3vkqVppernH3n2oM4bAgCU8wwB96I15OS3s/J28aRGgqcYSgrGqhMIrAPaXuMtGON1LkfCERkd
1IstQxHdkrKswww8lptzapFTnYfKDnB475uAiq0fzfskJegdjNiMttVzDloDPezwdsYKANsyfcBg
enyUuIHjX/ZgVy3qAOYJbWDWgjCeD0HuZJMrlECXsQE0GTWMaZHnB1YE43jdDLCjsJYd0oBGaPFP
EK9f8iNa66hL6ZzCnJet1jKSephnEzr9m2FkJ6DiS1ZkeGXxrCtE8e3Jj76Tt1V1Pkbjzx5czsRN
kw/Fe5ePf50x8kwFnxJVcmP18afx3aoixgYbejPasT5wyMiI+4E+qPmqXzsXnMmIivYM2MGLhcHs
tRfoVIvUkLZ1T08YBJ/Y7GokoU54gsWVWxO/mbPO9GymdmxGQ27qaIWabnUvjSw0Ri2sncZRS/pT
PeZMy4IXxuSZzOQzrWtG9ExkoxjZ0NuSafL4X4UIVa4SiU95fa4wTClThjrOo5qU/CTYx1t+Tp4y
sJSXlf0it8hlQmjfq/HlmkhMB8X8nY3I+tjOwwfjDRgdJPoqoGWXHEaMU4Pmx3xzMmngtpgFIBTa
DsWtHG/addVd1wGl5RAQKQdxEYLdBm6hYbBPHpz9tKx2hm69adm6m2RNEgKlan8VrKjCpbsAqjX5
KEkxr2bNIfOgJBd/0bYyjECbLlQsZMbStUB4ObCl967SOIvXTV8esnfcya/cSamZbagBD3l+R20J
H4DqIwrU9OVF8HsHT41QgaAEtJhaNBnYqRR43JckMM88YfN2w4gkTcWalKC1WH8vwIuXGwebSIaa
wPkGJm9oyjHv1u9TNGkJCsFHc413b75yg4MClDdKCrwuCXE72oMvagC5R9aEpkW1BcmUhNaNqAOs
vwYPgHWuMvZsYlxiLqZTDyyPqmfTDnOmSAoOavasjssNHQehnQT/Jxh3+LfGkppj8C0MSQrBbQLv
3NyE9drnpS9cpfVQ2KUuzv6QJ5SaLa9HaBF/rmKdOBXxcaTGyl4+um7IRt6JiIuk6/2bHXBC/EjB
gpijc6cvGlsEZh6qzNiyJbaNLgH5y0lrEtIACir4JkXYwbTAmDF2uaJ0BGNRr8x4UNW8MHCa5fNe
Jx89Ol+O+gwOyhlP4CtMc390Jpv08dvb5HVywkFr20ydgTBjHvbsLBdYZefYRVtP8UZ9LG2CDk1G
ogOyaFkGlK03k91wEOZJpSffZzLmPY5+i/uf+rXh2bozxG3e5NWCTTc5qaV3PqtKvdN9Ad4W6YPk
YBKHxYVVKHYe4nnRamoFk3zN1heMeF6ErRly0MT5sfM3Liup52PfhurB0ZXvwzUlQA0qWiBnOqqX
aZ1Mu/jV568amU7ampXs/UI4Rwq9RMbIV468wXVsnG8OpzDH2fRoVtbtM3zA6BeAiWKwqMVJAJSL
5hqNnuOX1OiiIEzI1eJGcJc2wktEVR4TjBPd9RJ0CFJbxwVeZfhUVqgYaWEXxNXwVuxINTm9wtv6
owa+7piNygNVW12mu+saSXw2Xvk4DHxkmFZHTLOFSO224SY+TpBWpED7b/ue17DtLpDnslaZC9Vj
ya9hUrcuZ1e3r/QwJRzbmR+G/VAXeHn5dqKlEKYSNF3QBOoU9de+J29YcsJNzpsYnXl3ZEdw5ph8
+FzbwVOu8rf7PJg757Li6OmfYJV0otBO0iZ5+mM3+v6dD/QmB69FpzJH22JqGNhnnpYRKUpWcPrr
nIvxk9B96YdCSRcpNlDrpHreuW4Jjn4bMPwigxDV+XdNMRjcTQgEq60+BKtZaemaDYh9z4p3CnUZ
mjLCV9lZAiGY1uvsURC5QP4dfebpbqqOSO/U0gDf7HE4MiA4S65RffUAb5w6R1jLdl8uKupojI8H
SRWk4zNQ+2W6Go/K3GTVyQWGo1H6KqfQSUCkf6ionPx+q/ER0VnjtWYi29l5vVXVOdtCWB7eh4ve
1lAesnhLuXwZNzaVU3VTmwjp/ErX7Sto7egIn19L5+QbkgJTeJ8Nlpl8s5sauNUmKP4PQaKFMt3k
3RYPQuJtDw6ZEIwyrmhVFhyNBxvms5bqsFCM2245SKtXgwjRweBvvXvNgtaHJhRwcxGx+UakD2Rt
7LPdrcg9srSWesCxbbowc8wnxB5rivzyZU5vWBzQBmP6lCBHfAvqXRxpMud6HSzfRO6jw6a3xHJp
FnHShaneyIRmec7+9K1+TRQmPL9hIK1ItuKrAZUNiNTEfS7+qhqMbIqCQWzoO94GIfuRMQoebT9+
x5bqg683u8SQB/j24Hu8Nd5KahX/MNjLw8l2rhn7Z6/+BDEEjZcFZmq7vwcD1lAeexORwJWWvpfm
zMPSsbpKOz6lEZ+rMoKI/WlkJ0en6Wquo0Xe9zEpY8WbnK+QjV20n3mJWCsDOzjOczszzlFuIlL6
1Ta2Qx/0RaJR2j/j0YOP9LKECFIFLUv2zSArXfuuUNvqkis89CkUO9X+ubGbfpn6zoWguWacshjK
JupgbxYLX1uWSert5+tmt1HBqAv4S7lzgl2T3jfNqcGOeZ99TOqUfUBwwR5gmP10kib8jf2Z6D5V
tJ2/1GPMbiV6VV7KvPA/yEDaorbVz5m5aFwm7vnrqudTryzsI5htf8FnjEjbsQEOVcp/xwn+e4x6
qcv22R591fpUbsfd13djRJwAWZrihdSWuXO7VIzOmMhOeaFR1LONIOlp12dJa1Dm1roboUQsaDh8
u+wV5FSBqMbOk/1M4L/L+GjuYVkqMGw0ownTY/TCRRwhIYGhm1xVCe+BzbBOVVYkEJWoANQ6s+GN
y+BIUiZR/6jOYeB9d6fCZd+YVNPdF2OHpaNCFxmaeRMIugPWx8dOMLo80uBSbriMZlIsGDUG7UwD
2ko5xBAs2gd7irRgoogCNiTmbbkg/EOnS6EILoLWWO9pJZ0wiTJSnTXp5MSG//qoIyctFLwrrayB
fEOLpNfQvKCGtMw4E2da9xzpgGk+Rr/Tf/AyBZ15cE/zaYBD7/B2kZ3VhE8s712pVBIITUhiveQg
z0u5Sh2IBfqrsfh1s9Vb0h2NG0lq9MEspZTcg6dnviv9O/4LMKe3rtMY8CqGSQh7WHtl8cw2WBk6
ra8kRjpdXj4jleZF6RmVa6A26ezOwYfymR26CrAJsHQq15Tibxp3S3ZfnRu6lXA6H8bx7mB5NB8T
P/25Q8VBJ/UKF+cNnP+ogWLOVXLrGPYtCetoXsVglW7CZlfYcDF6xxFNGlxgu+Br7ASBa3FK5Yv3
fmH3hqlv7JEsRsWCD44vXai7JdbsoydX7qBQPiinEptDAuEyVQJIBfzZOFWWR9/62ZpxmDh8LGok
bVutI4KZmJcnKZ9TWEnEZ3V9efbiIhQ+RQrl+B+u1T0iiikvT1PfQobcq/CZOS7JEpcKMlOBmVH6
6w0sXhDPYSULgnAY6nl3XrJ+s7MleqJ92onzDlouUsMA6Nyr1QccjZC5viyFZEJ9AavHoHD0q3oq
mY0nw6PDqts/OmNjnCT057Ylodu12aCrQv/HBewQLw5IBN4lZdeaPhvqf6J+p3Z8pt2c1tsI+SNd
aarosmJpA1ZVyGCv9jyNcaPMsWiFzmINcMbFP3JTgWKhfSh3qpNfYekb0GT5oQBFS9n8WMmrnmpD
5de52DBVDylUt4e4IvZKWp4aJW69ylMlqu2C41XrBLGz/Q+dOr9BYTSfQAos95F0ZwNXgD6A4P9Q
Dalny1lZUpCy+vzWGleYMcjlSZuNdQG8sEzKA5QxeFHRlRQ/MqH8j7vQ6YAFbv+qDyF0ouY0MJxc
0xYZ1pviXrCGD+7b4xX86TanOlbGVqlHbEGK2s6Z7oz+GrRcggMIlbynScgIZZccWPIoPYDPFpZ/
KHdkbQF0FuovsAppxVt5eXtSH1Vn0GgFmdm+6hNVVxsuPn2fe48BcV+8Lve+040eUYU6NHKBteqW
uo8nY3Xj2qjO0hVFrqSebGCH6Z/Nhm+jObsifGWgqTN7+nzln4/23N/Jlj4NJIvJiYSNizhrC/IJ
Cv1Xyz+qvq2iUm/IMsywaml4pf/AlxlCEWXrw0FZSES4kPVeQo4cg3jLVj7eng9eY0hqP515S70/
JiZQUU2Hj3vUuA59yLtDl7BTai/fDtg2bIr2O1PNTOsZhGtn3UtyBjPRD1wPgmTIHBhqbPbsxplg
/b9242UQF0LqK57MILWW7pKDcTuJy2wVMzugj8NkH/ql1HYXGUlyIh1ou1C14NsoZe2qCEl3fJhk
+4t7Nm/9QL61poPHJG1rQL7tdJKNVxRFpxUdBU4CoeGmLQC5fXrJHhX8wPfwKng9wBzVKlAgfem8
vZAHzYnnIFwB+GJ4+d40oK96XeC6iVV3LukUBIvBf7uurOk9MXFCu0GZ3bXKiBY6w2Uxe68uIKKa
m9KAe0OLsRNGw4FUnzaC1C+TrvxBgaJ/LOmuFnrbFt4Qiejecc8jFK/x2Uac0AuVQZgETyhl3AJY
C7MtcUFDF44pLYSyBKMvQzU7fkwJ6dKqkTQo2Mgy105ItLRTjSKYHO/NUxB10m4ujSMKBGJF631E
XVFOtPNgI7pP8qSGaW2ZussljsaGi18h9HcMilU2tRuQgTOuL0L7Ydo1Lsfk0IznN7pSaSAXqAK/
QZ/wzaRODR/ILj/xpNZPRIFta29cnTUGviNd+KvT2sPqDqFpxUakkbbmYHflkWMzbvSsubiGH14r
rsIgdZGHTEIBdWZeD5i5FxpyAxW/wWiVhioBJvFTO6f+y3fdvK/ZAFdnqp/JV6M9JSx3SQukMKCo
b/sbSTdXzhCmq6VvDCs6lrU4XvE0XlPQxnugIUWkr1K2jZoLWTo4FURUBS8clBBerpTptB8TX/Lu
TtxLrwwll2898rkv3x9Bc4oftwK+WeG/GhcSQ5T+3WtPzgfwhbVWEJwW2BR0Zu4FdH3iCHinmwm4
1b8Kacc/ooSvMJPEyuYi+7PuMJOhB/bJnzUP/fqVB5EmKP/5dPhn7yfI5vbjDz0OF2ZNblxyk6ux
UNt6wA8J+ltN//nxlRfl2kXKeguh3+Zp+gjfr1CjsnG9fNp1SHJpdKN7soaJsyZNGw3ah9qS8q2L
nAdiuuLS8VeimsUgAeZRlUk+J9ZJUgQ3CVx+ut8NZ6phyG7KM42w3TloaZFKu2m4K5fmRp+Adp7Y
niJcco5trxAWdaKPyFOB6LfCnVPcNOyWl+nGkNwtgN4kc+LJQQ7iV5PCMDabxm4uXWmpvFHS5QU3
zNDQZgDU6+hcqQ4kCeNXN8MqnnGyu/40OcFjMFvXyOFZktV6lMIRLdQFZRND6YvCRQZ+Dns7bvRS
EipsUITMCdN8DS4862aIjfgZM1ZJp0dgROc4QtLftU94nZoJhWLi/EwadQnZjMuim6KisdWKiKC1
RjPDuslX+jvFpLLyfpz6tlluT4V34GwpCFrSdkVV72tVgE9qVZzWhrtQ+O6+dzqCfQS62fGBYF4i
Sy4HRm8nPGBYh7zIqi4wxbw2kfs5z1U24xp8BYovgrPdStcfUwHCNaMZGdTHoR4tODQuzK/T5Tzk
GsPkUviOop9U72B/tPz/OWObVMJf1THF9pk85DYa+iPsxVPYJQKuJpXWM6kaGmmpPfIT48ghljX0
Sqg9v4pdq9BRaMh+ZJKaf3oBmI5JRCYZ0ltcIyfVYMYfV1xg6kAEFP/RlPtCxD+v+laVXBc26Lx0
K1uSPIf8kebZZNgRIqh7F/uZr0+QpZkUooEelFw+n82y8VX/RIi4Omb+YNelGF4ucFo7hVoZtMu3
667uq8xtBbdx2jeBDvr5u/p6wfUuczdNhPmLVX+0whDjgQ710s2L30GX4iswBJCuvrU2h9SLdTCQ
lagtVZvAEz15ARJGUhN2dl0us9214i1b1WgxNLYcdYo6yfPvtPcLYPuOvriPSjURHVDBrexY3sQl
6po80Ta8CgbTs5yCLwRu7GKj8ilERDJNWO6DyeiifkYv0Tcpj4vmkPO48qVFzIcfHf8k7ybTjRdW
ZhckBj8U9Ww0r8VCRT8Nim/oajebmWj/2I0ppO2i50PaEGxJJCD7Cgd1F7ZgjvO/AVQbPXXDFDQ+
GUoesRhYgXpZ+hmu28+vTAH6ez+SCfbmbOSE8LL+xo2jNTlKba6Ye18oN4HDinTIEzdWP7KxKXGN
2saGCjkjoXA93lBNTS+f94U93Ybq9FBjEUDDoTKeYgUaudCaxbvMYHaWCBNgc9OzK7770++DxDH8
oJMIcEuMK42rCcZmKosZv5pnt8QBNGWLhCDQo0fzf5xy50k1YPXtJC8k5BgqUTMgygBYafo8zuPc
ZVj7l8vGgM/uGfovc9vruKqRnMD0Kw27JpJDrt8Aexy/0G7duqzP/eur/gs4dSyQQcn7Z/i/gXdn
InB7KQSmlZmy4Dc0d2OGs7COIMoVB7Fb/w5tF5GKhBFtvdbt9ItrJzACRRIncWU/hQKIbrcBMevj
hA8/8Lj0KDSu8K56nDnC0vpX3a2pD9VjtHnkBNvouh9nXHBwq1JdQuKz5NNYOkOUMIZYI9rnNwUZ
fSzlCZLY7mvoH9axPDzCulVzFefSEM7sFc0HXMLdEJ5Sptx7/gHJMX4K+hoRMlJqihCWfguKXXR7
DK7pFPTNTMoBr/mVXsfMfjXenzY21CDFELk2AY4v6qKLdfICitfV3xJy9ETBjH4vLw+5Vj8IRV5E
FEgWPqrbaQI56Etd86zHe3uQkTI4k96sxww61gRKd/8NinLHG7FEy1MTeo2D3ro0cc49aoq5Nncs
a0GRey0GSzuRrjW/5ZnJ6e7Q1qgv/djT0E7mMVxUYxnDzE1WslYi2SLg6WVdDMMp8Ywpf89Kr5OT
JxZzWwDYr/tpd0FnepvyZutYBKhJjVYp2rl1Xe1grkzf7O9aTRj5blPTJLEAWtgrtoqpmus7Lden
Fv97P/jNEv4t+4dcmNdyoXyEGyq8xQTbtIVkBfywDGioH0X+G75CSbqzNj6Cr0/sOh0byfT4t9Jv
oan2pMP25sT+SWupc9ZhTZD7IR6h7LI4N+wqJoLigoTk2VugUi9FteSTRv0lk6GlcPZ6tq2bA8Ds
Zp1swVfj/OEffYg10cP40LH2VesJ8MVs/MEIC5qy5SyBYERPmDh3SLy0tYBxG6vIE7inEDhNcer6
F9yXas7oJwVxIEmAXIucr+TixRtjkd8wmEOJfJbOFcoEi/7aaZpaFcS0cnPZ+7ycUI2UKyfZQBVf
yus8hP4MbmcrmMW57ul2l3PP83p44C4J2TytqvvOF4+6Rvp09RcOWZWVSQ07qkiGbP6HRK8qv4vH
LYsdcXxTLikK0dpDdDzd+sYkHzv9fg7/o1Vn8TMibk4WS0vWFzGNcFnONOgoJKwDWs8CYb5F9Oy1
xIF7V7jbHfdi1P4HthZT8Q4YdSR9M3tu5B1f43mlY2MNPhIM9hr2vyQAm5Am7QLnO63iWih5WV6a
B8oE/ZViyw4Ll4mBRMNsf0HdVIC8EZSdHazmUzt4PYZgU9nCRRrBe4UGAE7vpC6gqtw9OZKJKp6w
4rAzc9BrruVgO7b/+upeUeXgvstu7KQSkqVaA8BqBhux5TFd2fYzmPDZnUAbbMGVpn5Xcnvia18K
yUeKNi8NpQLRBvP1If/vhf0TVR8j2EcFcDM73hEEzckIHYvAOO6UF7g6ncx1zjf5nDisj30iDGzp
owfnm5O0vvJwryfrhXGVMwm/AqyQOTwQhMsVCFBYV7dx5gkRPe/WJy/wOAi8dBqmngxg523PmU6l
dcFXWPIXrVeJMyUsJx2gQ0/EbzK7xyhAGENLeBHZpEZQmIwBdwKM0yTZe1KfblS2dJRc+KDqSeG1
f1ZuE6KtzmsVoecdlrh3axoC1uECNUxu4DGvbJR/GxDa+Vd73Vc+maLCa5naZpJqSihoLWVkePBU
khQE9Q8iE7Tdw4MFJUZbSPu5RlEzEL9PC8GFIhIbmV+6RRtCdKGeBOfh2luI83/7CDImTayjE8Do
V/0hyvJL5lhRyqCOcziIbDWAWoJatv7EM90Nzde8aPTLJPqAVIGBmqlsuXL+5qi1x2K9Zf5C459b
RTgiRMf54sg+7jcjbEKvE0P59JUr9MbXUqGE+6jGcnG5XzviaFneGOmwl7rb7UdWO+IE+9KgKqEA
0vku+iw94vtBlI6C0qENU4nuzaKHn2RaHijD1OzppaqAFBRLNi9l+KLCBjdJ5koWBuZQdHTgJgyv
rc/3E09UL0QAJtxJj+SlCX2m+wJF3QS8Sfz2WmDO3cwR3EauQqpANwMLoDFHSZdQo8EEUKRnRYbg
uDsmwHtzj4b8fNXi8ENiW/DR2hkp/+Y8ViQHUML95/hg7g9O0k5XbBOz4wVDgbckrzUVFZKRahAP
VTHxRZZo58GPqlksRlewWPixoOdIlbRGXgWu9drK1kxhMwx0OyZDsryRfcGRhdSsfgoEwcN1uvl7
pqHze+cMaZAONUYpC/YcSIMKeR6eoKs8kacNntDskF6tr5eDuj2mBND36wMj3cMRNH5EPWk8T87Q
ENhca9fSGu4Pq9SmLjjM7W1LepzCkeoSkfzL/0ezqN/3JYL4ZDqSRMMdpmrT1QoKq/IVCXWHnYFD
mp0pMwQaVyO+nCkUadPEYwo0Qlsb9nvYw3vBliPaVM62E3VOwAn6fS6+nJyZlMnKkWtUwdR/qcbq
sJ5nCbwTFg++i/hNCiO1QeENbZP+Gaj+Ryc8ilUOLGrpFA4Y/MjZQa4BuWb75zpbo/VOlEMe1vls
dAqOYiJNnTxdQ7CjrhtqmULy3M1RM6uyLyIVbctAH2Qh8p6mLRTJuo7mdKXs2h6XlWiXTNy0zAeC
CJf+2A3WtzgmhJypsY9HsCm7vWYqHFbrO8TSl0V/BBl0Qipcx/+gdweROlgjr5WzYrluIKq3agvN
DYnkTy9zVO6Um6fAFEdSAdMF+oGkTHsHX8tvUxhABIa3L1ZEyhitS7hZkQHKjiF18b3vrev9MRhC
nr10mhbn1Dz/55ex8/mBkgA47fDqUvuvS/RZTV023kIQXgVAKs2ulmj1kO0GeAzl7nKIGVAAamLi
qjnqCZvdy8oJHV9XQ+g37LM5X4E4Xs6D9lGr7XYx3MW4dv6AYJlPPY1zZHhWFNmn8EIhvQ9u9ROE
8clOSN479B59GNxLT14aiq/LDe24eqFCj36bNfSsKNCxhYWemdfPvLjA1wn4KDD9j1HJRZrSkZrv
GOuc6V6U6WpJdLsC3xktzE2Bhu6Vkr3ml/HYPcdrNc0YOfUlqsfLInuLPlBXeP9iRJIXwL7kwjNY
3RlI/XuCaHjDwjm7gPSolbeOHI+oXlJYUUYrA4370pMdeXbGXC5i49IPA4xdQ5lgU3aRUDlG50lh
cXpGngptMbukIqMVHZksCpOh2/NSQ8bM6qfk5u9EXkkiJS6aQucrIy2pFnjbPb74u7wFfyutjmaZ
TJaG48VuGFGRXLzJYARRHiJlTbADat3/vA/EPR8TV47paEAbn5+d5n3hkAcOW9iNAdQIWCWqCX3P
F8zeo6Tf0SbVfCkR6+Wou5KhvjV67w8e6izROdmfuDecXjQdGU4s5lLAuRnQvVzPkoqJox45Hqdf
xFDAHteMuTY4U51KgLYz1HLSLRjOkXBR2qONVnp1VBewpbrcSnY+KAnZXUhFTCuSpatdoYtdu6gL
Jfd7MEFKCEbHjVxtMoJEe60cioECZ5EnQKevJakukMRXatXd+UcPczy9XBug9Ueg7lq0MHgFoPay
+dV07DViAKIfAD+uq1t4JK4my6z8EKzB5ln19u2ClF8uNh1ZRJZY6UN5s2em7NYDtl9qsfCmxHC3
/9EeagNHwpotkUHqdqtatgKTVpviwVpHr4v+BaAABB37v5/l8cQrH/VSBtxl8LnHyLatXBj+inyM
sVYVeYu4qI0rlSGC5XIeSzGM0Ky6ilsUvIOyLd9+fxrdpK37lhlAzAGNjGzin2mjL1IaYwAe3NyG
buHROOyWp0fltGtJtOd31+mhbVHsVMYfOz7pwLxJSDRhNljmT4QeXBM5cVCAt9983geKkovPjzMp
+wmpCP4Ro+hg/m9n65wotVPmTG81fYrgVB7u3+M/LvnRtdju3up5XN5i8SK13JugNRaAiuySLrBY
MficRCStCGGXiRVGRzU3JaBQzgus/g9ruytH6vK+w9aRzUML3CvR0PYYmkBr2LUeatZZpBtj2Qqa
QrpENOhkwXV0GFpEeXUgyXYriaiYi8kVj4GEuJjDafSBikEVcuktUnlXNQKY3Iar3Z/+s0QsGMmC
nEVjzx7RhDFmo3zUSJ4bvPLx9MpjtftEshytgSCEmdGX21QIwXzhd0sxEfgr8t+ZR42toYddqHbX
UvW4JoxHjpbspTi+3ai/+dJvwMdCUSMx/5UdDUDLRkGlojAHDrhGgRb71d1IQ/QC7O9pYC8LRkCS
hw1DLPfwdiWS5XaCUa1sJcOMWID+9N/kr946ijx3ZkxWRc9gqwnmM/rmQ4k2+WhNFIueWquZC1r3
9G7tY/7Qpj2nDpUhpOuEVWLxqk2bIFze53chVsbIpDVQY2UAhYc0rf5ovpw70zuwWrpcuzE5J/QR
UEon0ssZ0KtMfFjG3vBOJkZtsTwOXRv2T+P3a01b8eDdeE1mq4Y3io0dxDGBxfbXK9WclZQ+yQOR
mtH4OnGps3UmtW7l8GwbLX8/eMKAw/ngrOSlAuV3jwazUIhevk9lfa29xjzAJrJjbSyKm/S1Eyhk
ntNmIaCY9VaUT4Qk9xid2HrIpjEWvmrhd8rnRlRinYG67TLjQlxjO0tZkHpGfQReXtpV833ph1OM
MDCGVVWFLY7lXsD5u1uczLVt9nWJHx0AcebF49APbPD7mpzU5PiY0J6M6UZgiVyPT/9KfjnvwOka
QceTrbqye3rx6Tf+3idmuY6i4q02i/QtUoGGSlvZhwpVgHnWsX9bnoU+fT+K56pUgPtlRZrdu8vH
QR1U51Scdh8foAqtFsBqZCpO7Fyg+eI9erXtiHYqtZrPtvXaFv/AOA8WpKmJ6dn9PJ+vJVUknOZs
Qp6ifpjJSXi31BUZo/BKY8Any3v3JPgkpTcA+X6ZTsFH3EIe9YUxzCmI1YDH883Nj9of9ouwYyB5
jWy/lLEi7L60Efvyr7MtGz8pnJoMD3gcEgF+mBH7LDlU6ZoXfj7vFy69MdhiVDlQjOhHZ8TXrFwW
Sx7363+tYXycpIfDUmiqVA03i8GXm1EDxVrwAopGbtdk0vHx1m77kq/YO3uLxq4IeVJMPpfmtnuL
HFseMIpx97XW4Hlr7aC6SW/gL9s9Dd9DxzUiEaSXTYugO6U57X2GH3fPwBmC/RZ3jdYARewz3Owf
k0Ds5t1zqRLe7nH8sfCQgctxNr4gfcPNPVQn9niNVsO7qczAqoN6MXx7dvJN9Ge8M2/ZyudTTGNe
3yYFu4m66VaozBo98Vp8aOv+bFxPCY/SUSxvIl1qs3y8758lh6RJ2pcjL0X9CPXAgVCYKkqWx8Xo
o/X9FMDb/BrEIo1pHEDdSZpQTVSRsSWAJ3JQ/LuEBPFvpadiXxUhQ2BFjqj04Q0o9POP7Yd8VC47
T+at9zWJuwGMMFxI1ok0b4mGQD8xPx8YfEmj31Ln8AgGNRnJxQeQgsqV+FDMv5dw/2HHT3a5UNd0
qOHnVWSHrmh7LS6+IlZzfXHOouHtn2QDQ0JC8a1MX+u8LiBVTHyIY5T3F8c7K3cT9ppQ1kr0o8xJ
2kNV3HCU52WHJwu7Nr+AwPNxcJLayEW7ZwsfpV9Q93xuBz/VHtpiuXHSE3FgDCD61JEkYfzXtFjR
cW2mR96Eeu6vQlzCoNm0aMDSzIQ4CtmB1HALQsrgceDYHbKb1uN3NXAUZnM09zjpwK6QrnwT60sC
SoR8rV7oSEN3zs1vGGu1asA3DEh80OmMNe6GnDPXokA4LYuuNgk+9yObwihrApAD28vGbU+rXcLP
HnF+oZaxzr/SarRXQtxCIxWsryNkTSpO7h1fUIThIkD9kYMJup9t69z0RD8KGWw9x1qnykY+BjU1
r59s7d+Fwb5GFUwmVHCSHzFOQdvoimFgbj41q0BsgCEpxbGC6quTd0bfUfOPzJk910JEqTI8/Ygm
sRyOlQD8mp2Tdcq4IuD+fSnBe+h/LlIUnFegRpgNMaNn8VE5MK61carIh4/Yd8GJpHrYzD2Zuf6p
3bF2J9iG3hRI5hGBFebvpV634AeleW1FHIIHX30LVD3M1/AKNcIfs2K0IweHFXq9fYWz4XVxFL/b
LqVLNYLSN65eSWwwS18iHTbjYQH4FGO9kalHgGA4oujc28aeWGKE3PyXvVBs+4MAYm1CqayAX942
o0PbldabCSPnxPSb9iW3VfsrUjecwIsfl8ztHY3A/jagFlOfcQMgg/XQwlghTCYQ7Idb+4sBzfF6
XwqY2bFLGNAZEcW9v4sCxcMfBuMhbMmvsQ/fDdbwzhNGWPbe0ibvPX2WDvWWmAyypvqCEzfsneRF
XqKfvOREqU/dSs4Cx26g48u+xUP8d7vwx8WK+tCEL0Pq02iJI0gl2v4Om2K7t3aCXmEeoh+CMzlJ
g64hj8mB6AtD31OCvIA00s2GJ287ZxgUO5v1rbahGm9x6nfg3dTCmHKLApUPTKYq8cnz0e7+U2Lg
eNQwwTc0O2I16pd1J/MBssXuqa79z8wyef0UckN1sr+uyKw4EsoIUAeH4cirlXOs8p9Xing3VU4d
YGekHBipW545yZLOeTOes3+BQG6qDE6M590qFjUOtXHBVrGYkzyQtlcgL32pRiQb0IbQdhkvkjWz
nyyak53p/sMpztynm1clOuc2c7JdEbg7cZwF+Uw3bHh8zKMTq7XHbIoLwcqgp9+EVpLVBD4gYQX5
jCulyliugqasT0KXPwJ6V6DZjoxXOMMGWq0Vluj2226jMMfSVSr3Nq+/IGbWAo6tjEzw09Kc90vC
dyLvL45f9NoJBZFbzMIP0e/UzS7xKBRW0I+5ioY5CfcGUltEt9oDjgxsp9ZXn6N+gQke0DWEaVhq
XAYWIkjBj0p8uSqgLgyQer8Z4IJ7HmEfF+1LjFa6j6i8U/5zverNkrAm9aZ9usdOaNiOjcWc8Jvm
a7h9CCs6hI2KB44TDEYUfImzqkwz1rzX4gY6hJpUwQH9gfvvgxhLCtRxc1lRnqBwLnVbjrv6GqGC
7ss6lGl0e95vhipYU0uIOS7nm63JMvDekMXPW9tmIvi4Jw2b5R9XIVeiwB08yjcu8H74uWPrY7rj
qXiLipaoh9nopVTA/RNkHG4Weu/lIaxH6qM+RSaVC5meqr5WtAw2atWfYKFjmgA64km0zaCVyNNZ
TPVtdGisRSdXu21J9llDNt23oSJLXOJ0E/2VmkQhbOk590hrrG9y5BxnkLcEDyBd6N2DEq8f09mM
yWlf/G2N5WCx+qIYhbPkInod5h1dD+YJhhnFM0bxzpVyw00rJ8NNx6CkDIw+jrYYSUDjyZ+DZq92
ihds2VhXBwNdYWrR1msKGfeNEQl3j733HQbGiI7AqIzOrfHD6Ze1t+yv0t1O0h3X6BYNwmUUG+zI
TdShHqh+Vski1UtqF/31MO7wyRqO3FEYaZZ3Q1U3L7WSh+ZN+vcwCwjOinvankbfQqqCI4W//INp
A5z6Qi+X7DYeuukL+mw4+5lwcEEo9t1wgy884xn1ByKfK+sCorpkcDFrbqQInbY8V/mjer+5ubBj
pFvOHZ3koVEmuqxvCGcFfSicPcHzj6aMH4n4+mITGxAo22HZgyXJx1qJSWzBSLwyf38yyd4qW2TD
dWm7F6LeUfxszoeo3iiQupty+ZM/d44rBBQLKetjzzPy3Om9Khu566JcqVLVJV6IV0gTpWfayDBp
4ChcKD1pYG/HjBqwzLik94SVph4QiEnWzNl2jpEqABG7km/F8IcUF4pxavx4oeXe3v1F5rfcytuV
1vGHgHbmxa56TUIr1jvhsfavZzlluZNVvP0TEFNy6IoF9HPRdOSls1CElYSfXWcKysNKK/TDQ7IA
4TFskuj5o/4lhOuIb2nNNmyhAH25DcIyufmY6lN7CY1v7bRH+VYReSa/Hm/Q0LnW2jy4KkGAqUT9
zZDFFKrfBLKttOb2mrPswo7EF0twJX/5T2rA9FwivN55TEiFXxip4aRUOWuBxMijfq7OMecqIZEL
OiDUaXRAXwQnQQ9HL+tnr/uAtFtk2uGulIBlk+DWN/nBUPwbDv5JudbVIvcLXR+ioVsInxj06tCD
UHmj7qjhTYODreuN9MtVRHzc6+aK+ZK5LkPfdJfFINyKjFqAOEpwaMrP3fG57qP+pjbZGkNuqDI/
BRjbPQj7iouIIt8cneCVdMWfcgyW2ygfP8VwGzqlCVxQv3TOjqBgQZJ90jHFhnatrx3C1fK3kmKl
tigmeOe3S0t/ngazn18RTghXwLIlRPd/vSjTnF5j/PQgG2Nc3bRxIJaVbJ9Au4hE8GiEuC6yktfp
uoRv7/ODBS8cMGex0Wq11NzCoo5COZqGHaYVVxwjIRwocOqbiSYYq1QDyr44zHkT7kHkumiFwHSO
6zVSxCYPWwOcxwkDUtd78PJ35U9jspXwXifkg4DiJe8A8rtfiwad3uHWTXE7YnMRxaCgjISY0VXk
h4i45OvYWTaufP3hlXrB2gwDXlONqLhylYcVOrKQmMI4UBsw6t4zqAG9HkkEk4xxjqkQ+phOEJQ4
lqTqWHWaJzXrltKlIp91Y6FjRZQcb1zqshQpoyBA2AZsTXJXhpeG+kza7I+wXo2UTv8q4in9FuS5
4dHZH7cYFsJP5K0zxpf31V7mT8bMj05NkaPoQOQRo1kXyhvWoQnYngtXUz/m0NrTwJX1Wdw166ao
oVf3WE46fHqzsxK3qt0GBiLP4KySEbSadrKIPr/4MpI0qVw9evxhA0UbPIjRYx/G6ZHi5ethDjOa
ynBVsDIToG/Ypz5bjFzjV6PkLTDauz75AfrH7sEf5H5qON12Jjsr7dbqOFYe6lac4vO/R/TYu9sp
CuHI8UduvQHhWOOFXoMkl2CxDw0RH4aEvab/0TXa6/aEkbIqtWknMXdg/4zQYutvTZHgBn2b9L27
xleTo6P6A8g86vEcHmWAiDbVNqSkq3b1789WNtL0NNOQWtRGkRmfEGJhcCetHlAHLoslOvMHpqI2
QSlSJjZLA8hHidgNs4Ijl8pCWYpq+c3ErTZUcI8XLv5xXUy0S8Ny/WVFqqON2QpGd5std4K6R0Gy
r6JbrUK65hchUH0xkcVZEmzTsGSPcRJdCBPDlsa/cC1VLDhnCV/ih99m8cN4XWxgUbe7BzACDXxG
PHYQDvs8a/XPlMLfaHbBDsVCELJNj5sAJiyZhnApjrli9yJDQZ16tg66a10TYoM9ZWE+iMLYcnRs
Sted8w9YcOe22+KKAMNSDRor6E5WgpRp1hkG4VR3zsb409mDjjZdSRLncNOcOPoFHB+YoZCVAzgJ
7KL4FGFVGcZJMCv2MEHQqJvmqEEK6vWFY7xkQrPjNKnI2R+QAjqyExbECugt/oxEIPaOuHO/QQEg
SYiPD6T+tHvYRR1qg0VpTMLOs+InImCjDhJa3zq7hlAWcD3DgnvtDnQdTiGt13KnjQZ0d9/7aa2e
qycR0aDf22vxytoI2vHi+shUNb+Av5HXUbm6DobHPxsYoYICCqXScx/yP8+CdjL9HFiNLHMesoO3
/a8SxYFaxzUn8mkgJ3dw9cUp4pVZcuPFHIA1zBFrpv8/1fO3b6RMteXroj/HOr+m/jdlrSOHHubS
2gjnvFSzyROkxSP1xkgkMYY7dLUYqsyBSpMKg0vKlBEWoTXTCKdYNpMdN2l011Hs7ikNvAagRZlr
qaOQ2xS9upMjMmrM5lFrDf6VsfH7+Wh4cfKiwiB65jDbiz8qOMt+tWbQfAbmMMQTmdyHjFDl/3vX
XEXLXAK+WVbYEhDLVdpeELmbWC09A0dtQZdMa1HddRJemznsrbmTCRgwW/vKjSTLbxjNdPARuvTV
Iq/80+riTf2yLHLeh3L04R/VHalb6LL5yN7v3afpMH96aXGqQF7stA8N3B55mUXqKn5L/Li061Gg
S8U03XWnQX29KnDh7P7u78siTdFSCSghqw2jpfWfvmYCJnFdhwMW7Nm8qABqPKKRZJqdM7S3B5PB
eaYFat0RelFW+BmORbPJhtq5QxD6LPuJVCf/AYWVahAupw6TFx0nxoCMh5a9+ylKoZHK5Y96CBx1
ZScAuHoOKuwOsatAGBYBsviq+5wQA+Ls/JWVl6Ah963Qy/h6GAlJGrkCybpP7fegyGuOaEg5FPpj
ciPdS1uoc2HV6P+lV8i9a5/GKXOTMp4uhCaENq3s1C8TFIEOBa+1AdAYdkbFFFC740Q/h6xebjLI
Q7dWzQheeroDK5gEvG0c1sfPdw716hFlc++d7Vhhd1qra8TGX6yG2usUmgaqA5YIJGfJ56YSowOC
QLmN0rVlgHh/GtKYVVe6U+jjdtjI+UsWbMv0Xv+p0nNeX3zt5XJTR+ktWmHl1K95boPvB2RbE3ZT
uyEguiufsdLF01vib4vqVtV+/wkfCbu9Ryee3BJfh7xW1OQ63RPPTHAzqyRBma6AX+ltjheEjAMZ
Xlt+FYejhdlGjHDxbA85H0EgraV1gNjoctPOcubwmEng8O/62Xaa0KgtygwcSUNdbj5qU58TtDHP
YL9SES4vg540iOG0VA3p+OgnFf4uL4bhaogWsepxTtFKqMZOcWei4KWdvEP984v4fbhBCcNqAi0y
fborjhY3Dpb7GFp1Caaf4UMNd6QW1BAggdE90XPqFkH9WmMBeA3uObrvZjYfeHFfr6gJ7U8W+RQ/
74Nmb1oJluE8nhqoL46EzBd7A29mQAsup+E0oU79vCf+fguTcd3pBfJGjIil0+oFsmxWl8Wl5VaH
nJ/qwg3aFHFc3cV1I/BM1hPw4IlU+M1VYqMixbkWKRVqRWDn0gkPfCWXK2bgj+W0VHj2sxGxBDCh
UeaMeQhYRlTOJPfxxH7qZ/xCMO/X82EwEQkkWBKIna4Cv9HdOgK0+cFx6VxVliQavrGNYI00LO1Y
HlGpfC1qZHHXEi0j4FMhqnU8KW/qRPv5gtrCjRH2Sdmf4ceIz7PqDyvCqoBBZvXjyKMzK8Y459qo
EMbqP9wgxtV2GypDZ4o3IUb5IQymOvnINFC7mdGhz+1xAY2LjNZ9D3aY1qPj8tXQO6J1oJzmAY2c
+/7JDiSy0TOIrS2zvy1SwV/4t5RtyFRe8uclKN1SPL+vs49gUvMQWqo1vjuRi6nZDCUgoLTLr7yO
h7GB/SDVGPKkBQ4Ghx3DUMopD6tgQWQ8oio2+7rVb5roCfMBlblgVOIsRUctnOxSQkpXAflkqDwM
OTQZFmAYJqdZrK1odhTVN5LSJY8eCPVwMT0lE7woAvGoc62mZekR2HgTmUcrRe8b90HAQWj6SEEd
1PUvc3HvW+mPXpqW3mL4ff1EiP6d3KuvivDFOHXiXFJ9S8uEhcKYTy4i85SUVdzv1fRF9Yv9vlUI
iGrxdhrcN+s0o0BZxlBv+/O/maqAAud4aNAN83GtmEYdOoaMVOWNdPIfeUG2HazgpHk4sfBm2ivf
vVaKDrF01pAXEWbDjPAqVgj1Lx4NsvYr8VSFDeN5Ox2KS9cUATy+emPqRPfpkhexHXwUrwvY2vro
9jC11+DEvyI+tQCtpY3ojoR5fZFM7PpcjnAg2gw/bfWj9qRLjEeRsDpY4j/iyIKj++KfvtLh+KJd
VceS9+aJsxk6Sbifxbps/tEtIM1DrE8AvQYGrR68Keae3Rxho3a72X6fK9OWbVOccar9zlEb8Utw
gmFYo41IxtuNYCfRvtn9Q/fji88p2Oj4NIvvjrWmVoiEd/2LH9LMejdPE9IBmqqKoP/fdOHTpdki
edsvYKdOntC9TXzl75sMkl5ANunWOcRA6KW54T6ciTCpwrY8eOs1iM7V//4w2pQfzr0R+MImgsjD
LJgh9o3WNkCZhg0Z1+uiWw1xXzvgaDwrLwi2vItTjKyRnt1Xrs5ozv3DaujfbCpTCyHVUscZnMB5
S0fItXMkvWKmR9SyyN5+685KxbIkfZ0ahWCq2w3SkZKTebE/xJOEwjTmtJsDAxXCOkUQh2LgtQmt
HSt156Jhd4VtTlCCnFVEfxtXtQZTDSAQzUYSkfg8DEGZFqBfaw4d0YpW+J3gqrfwL8soRcQ1apbH
J75I1JquOVziKnH1TowpHBcXpFoDnYl8UBqKLQSgEjOSwi6Peh9bdlxG/1qGwDlWuPJEo8L8DVQR
iVQw8Mki1LMZXpQekd8HIBxg+bIksw0FCAhA660tZBCHcOeWCWA5eR9PqGhXbV9HppULGIeK61nk
fJtp8K3LpzZS37zPdN+uOTVNR5QRkpVVQLcV2u/PD5U3Ne2UA5q4tcHAAQOXZx1smDyZamL8mnUx
oN9MMC0pF/UkP1Wd8bUvaa/oyG1ryctScf0vK3oPRC7TmsbQSKgedWRAl2Yx2zDwPZ56KdqG0oFV
fDV48usZxMWRnJ3iBbtS60imHO0HfZ/q27/TAwNR4s2R0PH8vhMIforYAgeRSH371UcJYneDOqsz
Dinn8dNvow7AiqRQ8Bpv+hZ7HURzUWlkO2jwgbluCP+fiLV+feQvhwdk8vS+WT8A8LfUOZ1V+3Mt
zIJ36Tco/75zGXoXEv45sPVi1HIMlUHl7snsUkXQucvfqrIL0+xWYSSVd/Ij/F3+GifNtfGqod2A
5197ubJFhPjBe85IKUrUvWP3jXbx4rLyJlseI8/jfLrjfU8fhXdcgzXW3WOgqQNvHtAauMcOrQmb
Yfxq1+4/tV2WUtiLMLSvRVV2NP6F2PleSaIna1v5MKgMv9CublAcV5UlDoQYmFM/jYn4Oz8554c/
QdqgWJtZynTvUUVRAsDqHcTuJhUyBKQIUYp2nxgbu7frAu73FBCf3sylsiIyCz3dYC7tCYWH8qZv
iWGl18aSM0xkqJVVtqxpSGnBTbwwLq6PRj5AcnjB/1Ytl8DDobg+O0YjLUjwj1TRgt7x8BEr9cPM
r6l1HMPpu433AdLEuGX1ru0OVv3lUf0sIHtHjRWu2pWmkUeR09qwvvejdAewE+Pel8wEkzY4Myeu
Kn7cDOCkPUZBymjwaPlzD1kAD/OrXtwND4vdscwWtiBGboZ3qHmv0N4z1/DXC+zRaqbZQw6BF3Nj
JILdieay9SWSiss7BJagwuAJ6D1bM25CyZKhlRvn1xCBd1VlrB8uHrcMe2FjPAabND6C9o8SSl1N
bjX1fknq7Ssc2BcjEF5i63GTU9gcZakQnnnheoDAWgK1ijfV3CA2GknaI9IQTcjAxmEh8wfTMOoa
7NzE2kKwKP+rHKM8R9ri8G94O3ZprqEhs4FuXDyTBFzrMM5nHtZ60ycNKLkOkdlEHDHFLeyj2kvU
qOoZiTUNHuoDWbIFvMopd2cerUmOVSxkonLQ8Wvc0IjyxxGfKqPRDX9eQMJv1aqGx+dYkFVrRkDH
jBu84R9QK5wgS0hQJnGZ4iNGmMwENA8MUkThsWoKetEjY4N5rS31Kts6Aalg5U0qJIFhRiLsT+ed
azlb709eA2/vquM8eB2z2VQm3cBO6jljc0+Rsaf9D8yI2bappOwhtWYxo1sRS4QSmwTVAtD4nVJ0
7hO1h1nLne2s4+YA/fwV8kEeaiwifVkXEScYKEDLM4VenQmqssJC3ve7lxPSedWIj0/P9NM2xOhO
y04GRgUxxDvMAFxoCP690A+8Er01VIULBpGjiF2YeB9cR6SqpM1Vwew29cs6sOj4+jHMVjciEL4P
maZsQFRTmBuNibs8KD+gAWCRnd0bl3O3C44SdjPk3XOl6wyB7F8l2+AsuGFt52Xb4FUQ7JoTrWrf
5M3Y4Nj9Dar+RDtqxpF7LIUlGiRa3yJ+X9r95ged3f/3EWfuSE0n+kbRBhPbqSqXEAhIsb8euDGY
wmoMYc4uPsZ4jeQfO3eZt5dO+X7Ktw0/pv/JrW5SLjf7bVSPq/QNHFP0bS/KasxJ8qAXi0q+3UIj
R5uGDStJAc2ncsR+b+zPR8dfqpI79BJnoAL5F5Gz+07A+mun52cGVlMxD/2+loNcO/k/OtyK57j7
vKVEl/dERwWiRF6qA4HwnnkwBTWn2qbbXGzjmls2qbz2yopdQ64NHqpwAhCzwM9+k9hwuii/GNk+
QcdxFbWABqfZeXy9BI7QWC2Gebub/LT8/SG3tvDp9zaC9rC4u0znQ7yeAf2JiWa4Ll+mo4l5vNjS
egHCmSKAmvcorhOwMvdOibGmqwXx3MH3wm8U2mV4DK+r0zEpSABljjdxSLXdqe+0VVSDh1ThvbOQ
qZCPPy2IOKihdIsy+/3eG/x4Lin1KiRpXbdr7GUJIka5nxL20zlVrYnPCuSUpjNHdo1oqp4ZbVCx
AGesc9Mm7gDufcupE0iP+gJOQSQNBfgE7tHSm1Utzs9RMx0tJJSoS9mProG5alGhtK/VfQXgx/sN
05O+BJ91wCHn+j7mXVnkYkH41YUbIrge6M2GbG1zivzqCjTk+QkY+RIaiMOKp4cBs40Np9vqTP98
2fY3Gh0aKUEB1jl+HcxVn8zk0e7PcVinGCylwCoh0tWClu4XRoVQ6xBNtBgKiijm7nByoXfYSYEA
82KZ1JcL/C32yNozXNBXrz8WwuqbA1KgeDQ9ka2taFfH1JEqMdsCELR7ddqludydw6gckkTxdCqI
P0ELmEO5KCi4H+Rzx43M2U4rAzSNHb04T+bYQhlFg4wh6Y3pxfO8klztVY3G23GDQUZR/UXDUCcb
pI1iPLOarfQVjrLLX+ZnVxJSfbj3mC7ILwttvLGv2pH8I+napeGqSIX9RGJkzOTVKyYELMPZndcN
/+bc7t84RndH5KbiaHTqyEbgCPBjIGL84paXg+Ee7mBQmzyoUVxH7BK7+Q4L5x54+8vUqwcYbgdx
ssrR3tHdvVbHbdjQd/bwfI8gFTQv626ZW857N9I2wO+uX6lJMNrD7gNYPMbvX9Gyi7OXj46baoOw
f64wNyZDVKnHj3JcflBOt1vysdi0D5xZelEMvNCvIsazPbhPNKJ7Lf+fTKgf18Iis81cDvG+f5Un
M1sR7RmfP9ur7QK2V/2k9iVwlx1S5HzgzAU5lh0xq9Tp5sabidUd1qMc3BdmlbhxeCh8cE9wju0i
+c9Z/ejFGse+K7L+Gi4rB1JmMPYfXImiBVJsgKuojOh4a0nvqdVw+CsuUhOzd2qlj9Ml8ZyhC0Rl
F5GfdfTvnFzhb2ooBL2Dbdsw+poz7wVJGk5vNLrmwVnQ0IT4UE+/FqFkPYQqANS1B+wV8mXa/rg0
U0uFcGRochHpyOzb8gO8YZS14MIv1XswbsXywFzYyExuH+/cxmjQ7dj3drVuaCVUWtQ5VFtGhlsa
h9TCH6r2c11MVaTU4t+dlcBL0asTnoTokHR9s3BdjdVGFY0CGtd+47cYQVHaQNUf+C5BXkQhcrMx
/iWcPZdL3koH5gN7VAPCTC5TS53ZxBJd28XpBUuQkRBZ6/UGLEgxlmqGPXmqd/WO0bc+h3m2J7nv
kWrQpj7mtBjrbQVobfgRpR2yLrgUteXvufJgqPQTiDLWFP1qT5sWVAWLFWjC4U7pU4rxZlHCS8+6
Uuin47HUYSElmKzaT9Vgnnoydz4fio5lxjhE6IKa6+SXGYTbNThThOYQL71j5OmQ6c+NDLv5axPi
3ETp0+QSp9xcFl9X6HRg9yyNMy6MtlMjWS1/c3UD63yQ9qtkiQzReEw4abm/MZK6ysVqoi4TqWH+
CDDFCeSXrv0c2oujzw5ELKZsoLrzSumWRzLy1C6/XJ16F8jbI4bVslxAltgI71OFV3TZUa4Vw2UF
FM/qwGgGDKFqr3upy9UB6yneTbtFnq7vuyIHOiuNPQmTDRq3pXCHDCmiwF+4RLzORsS9FKyWVEb6
WPsGjtnwK9p9gSLQb5z7Jug0x/BGc82YIQNFDlb0P9V0hdGBS+9cekDYKODHcqdUN01iw6O8aVDE
BXGYrJT4BFCiPqQ/rD4lnCg8MkKHYukXwwVxqE6S32r6agO+eVYSVkY0Hbsd76FZjZaN8eMKxkA8
F1DfiPWIjlFVL1Az2SGhCY/jcJXqjUm8h9XcJxmJEP6tbm4/Wufh9RTjy/wT9NHjLM1R7BVdSvKQ
qpFpt2MA/hocxdHkRMI5VC5wvBclpbAwkMeU2Xfftv4l+fWeslNlR+WvjsdE0j5FQLhEKAHk7old
ix1F5wpccVIxlfo5xZGy1Ax8/hnPnIxkMLG1mcvqRNFY6SiXFI2BJar9jrTmhFHezm6H78ym7BUO
7OH6+cUNi3EwxgdZrh3ZwBxgtEKAuAIK299kQw/bLs83go6xEDyUFxyv859fYMUMTyhkaqNuP9DL
NCMFKQHJnia/Kcwz9eMie+fAngN2lloMR6AdcBIJltc0uOnBZziiD4L3V/QlFwa6GAkSdYBPdNiZ
Fa/Yt5EgQfRguGAz6sTR9E0MHw+G/VBe3tDGswSg0Ufu8ekTNPV7OoLta8buggBTP1bZWP0l/MiO
FtfiShwr4NR/NoATwtuJ/2C6847CmVd6Y/8mEJ7fWCfEZ9Gt3J54Q2673zhWBdzHcwbgly4p+H1s
BE/uDrvxZWByH3S6X6Xk9L05xb+FlfAAAqQtoQN4zKmtatrK2MKRcwF5gVZjPlpcDQKEGZP7qyLL
woWfqhAqArmLkCWdROC1nec6fKarb9/vQ33Y44mKtCO76ip2tCFiJKa5aG7xFX6qPEJwboj6wsNM
j/LfkHxpIlzehoWtL38bog1akMQ+zrQs6SHR1iAAK+T1ujVpaQJv+zYNLNpWoM/1CdD4AZCN0OLS
29FB8QWF7yU2NCPDQtgH1033Tw6zfoBg78Sqco52vUqO6KaGz3a2SXrCLKShjpngwq84qZ74iu0S
dU/czEBmnCTNFEUCsb92cI71vhagnNIcdzTW9XgN2q0L1nZ5HZ6CiFjB6pXxgGOV5hp6aZfyjFq8
IVEFB7/dnd9doRiLh8DBlWAg02p5Scre7CRzyyevFgvu8WfBMm3wEtui1tmJC0vr2hsIkgarVr+E
fEOpunMBqmkWE2VUxUAsqF0vnvWCl52aE/4e4V90pN0ZTZbiFUTiZ6D67R0q85u/ziEg/LINbHb/
NtFE58OarHd7wDmZ9RYU02+cfSl0R4TIQy9vX4eZDYAYc0R3na7oMPVp8kw6uWxaGnfaASXNMcoF
5JwEhYFXx1LHMmkEyNalJPmqwTTWnT9g65c1ZxB2vL2xBHJV+iznteqLwzxJSRYvLi4Qk4+uUZVk
1qrA1zyoc7KPXUKXL629VHNrTgLiGSu6x24kPt9oV4zaOxYdlwvHiiS5Vj7xt9AKiO8DakoEcxbL
qBSMHqvVTRRR7Tdv9pdZhWvxN4s7zQzvz0dhkv5co+DnQO+gfgTw3zSYi8ZiEfe71U2rqfNPGT53
tMUabyQmUDDwv+sqqxoSphqoiVviK83EQnV2XXgA8TkhPzezjMItRYWzUFapzuT8tFf/AEiVqabK
mE88IHa6cJBX27zitoq+MgWuWLwx1DT9AWzJduUExt4CT1fwJ02RJUC7hAzFARKR8t8hkDOdTMTh
DFz0tMkMA3i6ALmFJcnfGNziICC3GIAHfl0QUy6FAejUHpvkusHMKoVHHT/h6r2chifcLQCPalrO
XfPmfx2dlPMuWO03skuVjDgXV2MzNN0XD+c09pqItU5JbtNzFnhGzVK5k++G+tKRYjHGwzcRq1v/
4dsUJzkQWWgavonNuM3nbP8uUnpdCBx7V4kP5E6q9dBhPW2csqXZy1C16++Sh19/uBAbG22oDJRf
eJD6wlTjlH+InPdmLmFmL3f4jWD8CNo6VATjWNjEaQdJsP6cYFlqagwBlkiTDieEuGTEsI2L2s8K
G+35z8lnWJBgzsPw7G+b81e1iCBiP/Qnb/F1vZqI/Xq2CF4vEmkRaqKTap/e55TqQgAVJWaPaKtY
RTN0Rcv0HPWZ5vp6kVLg8EfdRQVZNDDHpl0E0JkhhZXYbrjTmixR4OFy4XaCeXiUdcSVBVGSsy/D
xZnpCgiYtaRNlrVLchm0D9WqqpKMSjrr8pLLPl9JDkDuqjDb3qIj25BkCgmCwNckinsaCFTtuU0P
Cl03nopE22Seyfe0QUupdGduf2Pi+g8d0sVY9gJq9Om/b47DRrtuQWlgLuiUGEO/QHr5L0pfqcsI
bbqLlKh9EA+5SUgNkaWS6WsJTnD5E/7dA3fn8hulhCwBcsphNZTQTxz5Fo3D66YuLGdhReayiyOv
MVf0WUzJpn7U5IUF3MaZMCQ+kXC9vO3hTr9mUhvxUy8awpTyMn5HrZJLgkbDsrDZGESPfaGmGWyv
R4B+Ey/PC4f5M+6LyWfiVM0Hu8kI4diMI+YnXDF2HszviUj5zJMwzWnT2ZLuXwEf0V4p/elejJQv
xA61E0413TROCkryy6rSa6DkHKk13k55wbtG5cwOdGyawtRmfrEMmH/NY5kSnuvxuLcou31RF+qt
OBScM7mmWRXGBwyc3fAgGjV1jkeVa6A4mq1ZJ3L+ncz8nwgDIA7DuII3NyE71HqoU41JInh4hj5B
G0FqX1tQH7bxaAWoRnxiCjpwuYxvpQ79m7ALQm38H+OPh9q9X78jnjIwWXnRlKZPV7CHgOz+WnAK
yDMgF4bTUcSsmRGMknY8l3MaRifp39dDl8MvvmlRqSaPy+ztK8XC9SZ1JjH43XmJ2CdMOsZtZ3gL
Ga8ms9C8Cna8GE1a5VkmBsh7pgR7iwfC3Lkw14X+lLfafFukPpejXXApTWOmTIXNtt11PUTc6myy
ygO7eYtnxpkCLclbr5sahelY9VTs6qA/aXc4ZqrPc2gF9bfvOqQ+ICAGD+r+tNnIY9R+s0sr0r7d
gS4qjCDAktHDvxTPPji+iMPd1K9GiWFyMQSVCeaEQqmHJZflo/Jw0uzdBN6v6g/o9ILyhpwdPV36
+WrQIBsXvhqqolw7zRMYBUiaGA+j8/Fq34RKxy/P/94v66cqgBVYxodkY+i2xs703ZlP8wHm/zVO
6coizznJUWcq6MbZOX5/tu6AHzhe2JhfQfOJL4c1TXkNhmd9dSS6v6X1LcowJIRpJRAQfMvEG+1o
i9Kqp/6rQchxYnxafQkqWIZwQwpBxVETJXpGXhC44xEetX5mlmfjFcOkDrWa/w6U9+pfzCANQZ3w
1sUYE1Yy+Nd5PHN2kwkyLUtnJdWrFxzXpqWai3L1bZaZrKoQsFrkOKDM4loE5rrqXf+KVJa6nppo
x7RL8NEUnhIy9qnNKc+JuXbbtEUJwnOnsLGxskZ+9MSm302E6dW76idp6s5K3gwysJGXROpTyV8p
Vuzy1xVwY3DmrbJpz24ivofVLtqsbgpsPrsGwR1vnB8W4BL4DDMzKFfjRszlHorTyJIcnkAHqlO9
DQiFc74rkmIcHTtX++NQ/PBxFEmMeqb323PSYjNe/8/bd4Z9lGNlHLWWPgu8vjU74o3XUehdIVsL
r2hbB9QYCTJJJLegPkxbbpklcKhF5iruahtWaigrk/aetKgyYFfsrG8HcPOBbwr0BFIfZE7/q9R/
Fd+110I5nvX1ZbjVAdp1JSzZJ+s1wY0QZ4wJE1EDP2opimOU2BDRFh9afBB/ttpX6M1QlzzQUMMT
/wd366c8bc7TtdOTuZzN3f4a6euoLBU32DfYZ9/F04pu83yBWGnPHQsEjyh57Z13G6A1RjJR6/Jw
iwcvuhDfZJKUMbiAKCthG/jrEg5E0H1Kf1nddivfxdgCBVGPboDPAML/ukPSE1tfHJyWe7r9QpFT
snHnV5SiYPgFckytAlsBtKK2I7QuHsarpySiJiLlrfZEd6xoTOoM00pS45CJdBSy30M5PjEXC/3k
KxclXbNqYKPwWYPDkDbJbsCla6ykSmPVd432nISxH9DqKtWTlTT2VHhcZ49bCwtSNCzKv4di1Ngv
8HY7K875pR4Rekau63sQXVhGhpM4sN+/jeaOyZUfblbIBZLQjuRBXa2GBgzsYFrANQHY+gaj0Lpp
Av2bPd5pFLZ7XCp5iP5qvH+6Q6gnQyi5CUiR03Zg6lLgcPEZZLoGO09E7iP1KMJYWcVszsTP/qVI
hUbbdsn60wnFDrc9tqwpruT/D6l0G0E90rR74nko9QmUblcBfXWi2rbo9v9svS8UOsPlpwP8+aEe
COAqstqTtuW4sRZZSUZfSURmlnE5COVew9xsbtbbMkEb2vHdjbpHeLm0GXjAhjiotgsYMFkH2qyA
ULUOh4StNk1BdQAopu/zNubrzPa7hpMUmocVzFsF+2FAv+IrQzJEioLZYADx/0Zi8GhDTn8QXMBE
N0IugCea9GbFWtt81yilTqx4RghpEkyAsuTmZoz55KlsNun4Kirm/lVs2qDu97Kwz7YzP8IzCBl3
F6srH8/YhiNL8xBOTvs07L0ytXlTQLclH2aFfEsuWOhY3QRD3dtzJQH2miS99SGEUxXE7pirA9Jj
8euBKbc8nV5ZaCtUFRqZdt9lzY1w0lGOElm4sxs6whjt+YyQcZvqmeNtFg6dIEu5h8J9pSlRd8R2
DIU7UhhVl5pTvtzK80cE59W95wlk0qPhRJGvTN0qRLzFGz6UJUD2VvqbbygmEfxnd0nqlPhiWLTC
cxtd0a/64P5+mDpFbNB1sNij+ZVuFptJmB7dfjvHNmgxwqlDaKuIK/AQ3pAg45qbGkkzzt3rsrWA
zhjURZH/ycBGV2Txb17BxGsZynzkNH9rr8tJSwktzI/mH3ymxXUrZSs+SCVVhSncDbxIbsdHBOAA
kCEtAJyW1vk5mUST5irSRVcEhv8oOJpf/O+FFn9XiCu5u7BaS1s1e8e7wyry9LeY72+D6qh3Ry3M
D3gREZOARswo3zMasAqW+InMqkrO2xyR0U9u6ziEPhSuThQgPG1aBEszwk4Sd67gDX+jGOTBVLjU
yz1eeI/1cq+9vtZF2e9tNTtRK8CjXpsG2VfdrYYGZFGB4gEk5V3Dxremm9Tg1Ekd5afkCT0PVM2Q
XfasHNLuHOJL/6E/MYPWrhMUy+arb69Bz32wxAjeeLd4MVpCrpTF74L9z0E5lweggfYQcn2m8WGP
WsTyTuxbEX487LLBSo5tuA4nXF1ZihMbSMWzHlZxlsnYRQAoWNyUo6kvNSnVJLQhicV/i4SOQ9Lx
cOMfebhC8tKSizGl7e4YWuzB3C7sJzjkB95VvwzlaPia05yBwk9F06vbDxWj8KkkpaNr+2exqN/8
LWTLCbJqAIyuw+KbhGJjQy6/mi9MSHnk1IVLR1mQNK/76HtebwXBaPljqhD71QgxxuIghdSDmf6T
VTHKv18ZhOM3RgQP8NXJxp+7KfEHA7SOIGRWNf5w+rDaRtAoK4RrLb7DLHmGasJpF4NgCb7AAKfx
QNcI9zmh+34T9hmvLbPwPYdNsXbPW5jjNYF9RrJP5zgiuuTFvISybpWorpaE5EU668I1qgMj81g7
BpuZbmxWuzX01oD8hMtv9hqmgw4e6qpB12eKVMRTr5qKbxp/ZgpKsZsR7XtHDPn4mfztyhFcE+XX
xz53urj4AsD5cFWBcBk2f96lCOJ3tUxFBxJfDtfhJ1nF6MiLs3iUhauDi124dTk6PHz2HKalO39S
EozjDZnANdMhll2e909XfnHGC4D6K1ETzppA9GxwS1PVefMH5Zw02an2r39mcG5QnA89j6WtHD8y
NHNVY1S+RZMR2Dxy0/2xiXmmSm738fgWZJdb7p8FYTzLrTl4C8yV0y3JF9RSdfjdzbFt30jj7GIF
jPQAOgS/BPnx9mV/1gI2VTsoFFBRVTy6cE3LwKeLVed21jjuMxb6HooUM8qXmNtq5l7cL910fYbL
PGYZAhynIMWr5oXvWDokHADDRjebTeiCu+l15b/h5pUmBCLYte8IVM0wOr+TiVzV14KwUyaAMGJM
yYTiqR169Ee4nuawN5R5CqLSwL2mB24CKw1U9eUimdVdnvC6GNSBEmlSGQNCcieC+Uq0ziV9hnMl
FWBVJX0Oecp8BBXmK7noC6G+HOa7FJ65OLfcrWwpLNJ1kxQyDDl/hk5MyQOL58A9mMMdbKnVbbpu
X4i38INqdIj1HuKwl2HznSTEA+YlGukvWVuVPinnzbRyax/2gBGOGyM+I9oYXxLCp88/YlWSJMkd
yS0WhecoMFUAGEK1USE5CZDnXDOrVluf11O8c9EtktwWCiE7eGvdx1aVcE+R36e1hwU5kOn80x8G
fDB3JojukQ2V8dx56GcAGN//F/ZBYIXHK/enOHC+ZYw6ZzvMiyZfW+0F9JS10sDSh/y/SOTL7LNS
eXN41JRDkidpiJh4PeZK+L8lV1D/O/AKTjNijAZ0o9yeW0OOoNoZCXiVKfEX+iGLTS795Rk9w8zf
0+1yDOLph8mBIaWBgfPOylvq5t93VEgK1tqGt1pvBuFxr8M6blczy+Qds3ktj/yxnEfd9OT4fayg
IyLOFb8GdwLQPzzCWqpEXhj4sXmlQhhIHXZnPkFPZVouYbtBhUOwrmluj8pTSuS7Xx+aJwV7XGSZ
TicBYMB1JgWFOXVMm8ZY2OL8voBfoqJ+fieIjtiANl9EfGvqmlqR7nI9Q2kaBcMiy93o8X41sjiT
/XT5eYbxk4M0ZlTxeSa6wTPuO8MBnk25EA4mx5ZTwAL3Idpe8M0//1WFmRKXmwWxED8BTJUYFLm5
3dR2uxhGf0Chm42pxA8RFs/vMIBqmOmvYKPYKeO/vLwb1/O2yKUuW002tJ4yE+lzCbbmB7nRhy0S
tJucf/hfesdH4lajzYRKhFSjRuK6gxnY0X7iHyND7XgCxnKxRPMuS/1qDAnWpR3rJLDI9xPqC+vj
gfVexSgKLofip7QOGiOzQUskE288XXKczP5mW7FamTucqEQVC7+x+OnqN7++Z+jj8L3m0TP7NWhj
r78Ys/Nyaq0TlTmTBzpsfZty5cuCk9XkjsAWbJFu7qYh96j85wtbjNI8Ka+KfZnbo8JIeQWOJQnq
oUpzbj7VyUAjXCT/l0LQ61syY07/J2v2F1wySPP5Qqj3p+7/pHIN1t5sxj7hmo8fp6faVjhp9jar
uqesVS/BM87P35hdNQRlT21pI1kQIRbSQKCg5M1EmRiSZYh3ydcqp0NxeAPTbtTKUGv9vcWcjbRg
gIw5o4JDbgRe1weGBy+Se/fF8ILygZqekyZYwFVdZr5CBnTSgEnjHQZXXJkylDVXzvDkugTNWT3/
iiQharnXs0g6tC7KDFtYUSD7LkW+D31sj5CnXaLLTwm7SNp6GIGmlmuS4JLxtB+BrM0XpabqDLcX
uz0/Fdd+dutsM+R4hnyLDMHCBqP3WrjForrpADRHi8Laf6LoUi1mJ/VT9z9MOcBefWtw/EYeM5Mm
7x7D8zLZnmVgwfEiJ89oPclhiAHDomc74n1rZcGGvP4APL7pdTe3PMwQcYAe1qWN2AEdPLgZD6rL
eGMZDRR5Dx7ZwVjEd1uxTuunp1cloCc5LvXIqWcB0lEQnqKxYHG1CYV0c6+Gaf1KNroUlV9kdBz+
JKXL7gZo4vGoos+Lv4JpEFfOmD6gO3rnxagx9QBQ6ZRrO5cdVepi2k5+ia2EOEii2r1Wgg6BhvQM
/DfUO3cZa0iyofuKJFh9Opkbs900AB5qhiDNp1gwwhoGjLBGEvXbvRptUrNBC9MKk828VjbMjG2e
XeOEKd9KFL7xt1DntV6SrOjlq6ykQSnLKpn/lZjuzqx0fUVaBbpce/0BQPOWkTINUBLapFC6mIfX
+gQKhSJi/myYmrMFuoC2p96gB/Dp6E73g/w06pApMW7ILBbreZb8CWtPflQssQwMvSL6YqHp8lDZ
k2JXJs8YkqdaxwNG8DbsXCzY8QpYozq4hWILle9khmIFCzHAoBAJ1pcAAkFzPUfEbpqfY8x9+F+5
1MWSDYnLFCxq0hOdGspPy4eEs8+m/4/uYDHlW4CEaEZ2I0OPJnZfg4bk9lSmCbg6jYznZcPA3DYE
FbX7+ssD0hGbukADNMCLmR5ZwaVWKdUWuEok3/uE+K3tr8YZFCh+ZltlrAeYInAnVw5ixhQ/qnaV
hClwpswskbV0OlANaDNlzueddwhuGjBHXNTMO1uKsssvHG7wit81neMdQF9FNBvxjb86kGXd9j4e
nABz0w8e8pnBeidv1AXRDHtRWtq2lp7Kgh5tqcIQ8k0T3cmL0kRXxnd3v6tKX2cRoxljvgg08hN7
PNo3qxRy3pF90uNkbYZk8/7rjnJJQd1JScDm/Bza08YFOKtWg5Kwpk63/kM0E7q3Z56iqQo+pJL3
E+TVIlQ71CPaIRsdqKOK2h4zE+4ombv9tg2FJ6TDBliCOME9M6k/HlDY1zdH9zRtmtf31zZPNG5/
eS0OQN+UfdqHRf1TVaFf4gNimttzRFAM/YXxqd8Ms6ANhGR3Oqa5nyHUXhNIEMteL88cy0ql68v7
1jPw4bUwtOnTKTyIx7lYh4v/NN3Zg+3DFGtILUMOt4HcjhJ3CUky2nogvwXhGPB10u7Rfvcwg0CA
oVnNwym2wk1JLAtdLLLB9cwTtO2E7GQ1OmyhpccIbnnoJnDUoaS5m7lMTmQJR4YGc+ohW0e9Clsb
GxfbK4BLGzr8JeOcBZ6PzBnF7WyMZiGLEFC+X9LbUcX3uy05Pds5l/9iVTmFG9qOOB5eknM3SvvR
3l/cQoxpkt/S/X8sYB/LcfHbBTRasUaTfC/qJtS9bEiYfycu+I3tjdz2c4qTmXntbn0+LANx/9tx
5x1KOn2BqrabAUfI5Dv6Zu+FeaTfaN0du/Nj0JzMIMA/T2yL3mYEAoMQYD7Fka5//6GZawvH14D1
GbVF5I/NxPpLkIwrrI7PqbMjRAR+YiZqYgyRBgFlpF+wboGB49O7JyQ3DXFvbefI3vtmy0b1zLKE
JPQ8ak0876uwjRL+Sjxuqt6dxWQ1jD/PVW1wC1ZJfchXhL7e9Y1Z7+fuq0SeYzEy5v69tKHNy7Cy
YYmf8PYZPjMO6hJEnvL+J1OOov1LN6j480/HVxtwiZTm7Lsr7WXqSZ/unnuNeINpX00D8lr+mXpr
CFomF5xq2bnYSgmVTS/cce//MW2mZI4tJT6Bdp3LGljqhlOAH1L0KXbA4XCSsRTwKmdS9HjE2BO7
FQbJxgCphDojcMA907uracSR9BSpzH317RS7oI+16eh8w9GUnvXOoZj45PiAIcM5GxrgriW48tpM
8z+ifwFzpWzngHOarq9WhDK+0tyyAcbtYHl/qmjigCfsUfXSU/aiJnG+VRGHXV0zMjMh3REh/wch
Jg0smRuhNqGK0Pd5BVjJRXXyoqzBooh6at0fYVEWjBzJG0GGpmTYi7UVZktv2hjKzAVKSlpnx/0R
LWW3qGNDs1E/xuTntBF2YdJlL51uf+3ttYCeaV/cDYF9v2W3A+jaXOpGocNiVe76Vb5w/ypwlkGG
c1YR0/lPLyaN7PSl2N234IHz7qTAZ3j0H53iEJRiueNBTKg1ui4+WGj6LdR9g4aPxxS3Z2WQyVqy
WMdbaBeSWsa72mPL4t0QGkdtr8JzIC4QS816nYtQyegT5PRDRCcidOreNSoZSV/NNaqroKMTCIK6
Pcd7+JIxA8yKx/HCFivizMS81zsMOxnzKnFbu1kKtV4sKkK2AY5t3GwQmQAfU3hJW+kxQf65DN1r
z8hz0qLp7okYgdOf2qoliFvcP/WCcFVs+WadRcfo4Xx2GEyV+tmSVb3wTmQNACL4xK+BvLIFgTrY
vGK2VKj6KKtvHiS1W55zIUYAqvbhc6Of1lIKC6n02Rjrq/aWUj9B+61iI3Y0bI0bU4nVZbvYroWQ
2RuaadtQhU2yCbMweyuhpjWC1b7+ncLdU5UoK09wj7tb7aGFjGBg3op9x7LSDxyxRCU/CQUEfBGl
2/idxOyY3QUOws7R2OuXvpSVnaHjqiWuJC+9T27JRaWs8oyhGD8pbIJQz/UDObEDiXxvxWPfz2YX
5AN89pj3Ho1QFwKsXGauYPNIE0m7NMn3D0YBG8fgBkKEmzckHv53JiM6zo7JW/YmdrJnnRl56aYC
BNVAbZF3rB/h05bz12dJuw2vVj3fTXOo/IP9l50Il8cX+cgclWZS4mq/3WsYaiespEiLrXp6KAl4
D6e8w1H3cg+WvGjj0MmX1INtKxpzBXgnn+ulCrv5DkaG99kM5/p7h241B6Ti0H7mqs5cbYTqgOCQ
gk1rHwisL0Ik6C2bNf2/VUaG6RRvZn5hG1/Ua/tqUgxzOlWttYSV0cHc+wPl+bBkpWJ61rqyJVZn
okm1QUeqsrBYR3+PYozOsDZqSJbJSMX7ZCpFr3wsc6O5UC313GBiBI2eYS76ck47NlfpuGGENmUc
E6M9D+0EdpLmiAT7t3hnA1vWMkx2XfvX1w4aviQxwBLoTebN89LVMpamAcRhUy1PwsEVDqG5gPql
qEUg4vWaN0Qg6WJFnmgqpb/NGDxDfPt/yVQdoWa7yzrjS9zbx90Kpd9/U4C5aJ+7xbNLLmOiHXCV
Rhg+8lhK0pGyOM62lYvVikj6mZ08+CNX4glmCKi4DnuftFaK3YoSpReEI49AUztvQWGPQGAubIaj
xqaWGImTUEBNt5MLg0yYQCedFlnQlY4Ud7YaiB2Ez0gnhUXNuCxkEXu7SPG8PQ+0RUvP62V9S1Jt
hE0m4aAOjyZI8PFIhZ4/+z5lY/Vb8AQx3DsCqbS1GKedO/jmxPB9ZUdBNwJUB5mZCdZBCFFewOya
0jmM3d+8ROUaIx+5TckfPh30tZGwebrA6nXGk9MsPaGjzx7PaSab08/Ho70zjhIpnSbBQtO6ggzr
b7lOXueeR/waN84Rwidwr7HnE5LjCLXV/VmtlELhnuXU51B8vHhdBUt1xPLO20PngxvEFSbvmrgw
ut92ekIc/a4tx+HqJ+pjcfxkzqJI8rNntYfh8FBE9SrIuoEO4HXrN/en6UqlLALXtaL2bskldLcq
ag2lcPwm6Q/51KqIC6YVcMcHT474H1tiuvCfHBC53sUnyL14oUtl+HAiom61SMfW+vm/joUqKk67
alKvYeOwKSf3V75ekjN+zbLRR5ccwOIIZkPiFK/yQvZDwnb/lw3CTEQCETxjerdYOLtiGrnJ3Ys4
Rwh4Mt+uqUgy9wr+EW5y5817y3nbncCLWKkQEtBvpWbbRkq7FLaGSonLnFNtHGqfod4tXBHo6lDO
sPIuK3HOc754ExDLubXzr2SkC7U1VPVaQwwGehzmerLlJ6vh/DNbsVm0R23NfZONo70w29w/2LSP
2Zeh7Y8vSLGjl1hMm53PhZzeKKEqqLPNRzInpQ9SC4eDEMtw1cs23SekLsqVYsJJQAR7xfZJNJg2
fdcoorOFRkHVV8SApze32Tjeq5Lm2iQXQm1mvx87ys7iBKnViH5je3ozggBtVEY2+BjT39Bca6Xk
9tXz5ln5GRhF5TPdxlhUCl8gAz3tpbNkY8oP3pxLm+Gt5HkrWkvROPUYvCbGAeKAyo6Rfhzq4A1h
vLGI2g8TVtW4JnYp79vof6yoVsuquBTo8KAsTGy9syPEC+6AO5XOtQFxCPtAa2kHiOTAyiW73gWS
v04+Yf7VviIqwNnZOsBJb3PoOo1D9wuJ0a5moJhGvZF1R6ArnpyQgdvxImuXYhB0W+zuVm1EXMqD
RoPqVIXXlhn+LmVMN9xzmgQ6aQCSXp8Uw/QNHJRytyyl5obW9oHJ+/gVo3UyS2h5pQUMtQ9hQV+l
2fw5KG4KWQY+4C41mVeO91KpaWw9ZRTMpUZBKaI3HGWaXFbgLADy3G/NEGKIHfN8xQ57CoMHwfUf
Qzj15Ctwyje0EdF4FKD1zmXXKIKwF5oqLnL8ND/v4xDDJk/K8EJsBc26iz4dXsII0euCyT1eRO/1
R+pylSIVG+y+aEEHU99SHDkAqk77RWNdmLGy3/12Y41O++qv6gune/okcjx/OE5nQBA9CKsPZnm8
uMAbDmMxTUSXFtLhYwmLY81RP2bZWEZ/q3F8LuOQCY3xRp3g0CIl2Fg0mWUbBY3OwyOyAMeX65cB
e0VUwdgzu0Yp6jgC2pu4E7N2oV2ILMyYppnNiGbuQWNeRrB7qp17uvL8Dn1imErt746WcmkN0Vwq
+Aj230ziwVclaEByDstR6ikQVPJKBGcapKgDJE812/rtLGSQp3IzAM2bElw67MZHNp+z7iUbahCN
Y52FWtCzIoS8l+EM26MhHQYYF0IqMSdXgjRqxzEcZJNB2qVrudB/lgv3S6c/HUGdDeSjSbRf3dgm
g7npbdVYiFoxSn5EwjGnqTIidRcjBI/eqNvopXzwMpWOIoAeGdeFFAtpru5k6WzH9bPo9LjresU/
xDQzODIfEyLSe0VEgB6WSn0MTjFvyH6L4DDQH3VjZ/HmKK7o/rDNbfdM8R3DtaeaFo6dCl/XCzh+
2qBMZOR0xP6cRWUFlYoDlM6seE2HsTWBoOA5BwjrVH+XAqdX4LHWORu07ATFbSMuhPElRv8c0MC3
CB4QNA8PYCjvPqR688vArj+7CgzzCVwM8kTx2D2Hd+f0STv20GNa2XT9Oyo4eY6+ECfgD0pxVlGJ
iK7Yu2tuzIzLDz0DyRk0i/1hKB44sy3LGIo9SY7egG6XU9KJ2t3Uo7IgAQw5TUkeerIQebqw2luP
dZF//BS7wfMXjfgtrGkOD7bgK7br0kU3PUHUpoydmPw+1ssTPZUlHfiZikyO+yebj8ITMN5BeiF6
CUVC6pGOsFKbtWwChkU6ThHAmbe8dTHAdG/FddZw0NVLJIpfWiEHA6OKe+W10Xn+exiA/YFVq7eQ
Cu4iLJXrWLhrixab51pIGZ+EA6nfCZj9VznxnsOJLWsytJB3XqWbELlB7Ecu5qJzkkAlTQxOtpy1
uX+zlZsX6VynEbnm9MuDLEw6St5u/4YdP0j6G1T0fw3flEudVw9gIfJYBhOHlulp43Uucp4OJgss
jF5RdO74DiyOK/1SoQkStjDqUTK0PqV4Vid7uIu/sz8mvnNXAkVFkLjhxtcYo6DejrmzsYZ2Joms
gFv0I3F+IESxF31d4ObOtIb1txuG16ZH+YFwoaVAtDlhamNCZcxB/LWHYbdqDvZWRKChtOpN1XUE
BuJjJtqcSm2/O1uTuqslWeTCOCEpNk5LLcIh08TnPZm4TTqC8V0zEg91jzWqt4fpVnWPRxuBsprk
pmYKVUIOPjOMLYtEyWGtkmw+3JufCF4KX37gvWgXpW4b++Weja3h8AlOTj66pyEurXCusGxjm94N
bkOzT09jAUXTp6Ztrgv5dPPkyu1un6/mxA+fXnNg4nwI8K/eYHHsd4Wm131wApsslgwecRje8thI
GoW7D8dPAmTMEd8Q8Q8LymRzUOnLd8LvBPHNCyxdGF/jGbI5WWaH5OTa9aPoyfEYlQM4JzRQmJ5O
b7bGAZc06u14X75N3g4yeaJEELSBQz2f77D2s+GgybwDH4RXup/KTWVT8iiVhjbNdxk22dbt3HQE
isp5EDSq3R9+rE6f7eYxQU0kSnfqsRK4NADCxClA1LI6qpmmQSTCrX8a7NwRUQqN30ysYkjso/Xh
NOgfFEgTo8YB5h534HuxgUU3bj5SIvD1WEtXR15hKAZzXp7zkF88eUln5UeovIqM63haGssXEzyU
HUrjmqAWjAMO3npX/cWeFasSVU4kN8164CRUhLzpWdY1g9gsuyoiLhW2ol7Lbxo0Q+/FzfFM4cQ2
wl1vJ79MuZeYA37HwigVwUsvrjqZYXVX3nB+GixPuk6APLpPi6zsnvsoCKtudw9L1ami4fxR7odr
+wFwIKzoQTamJ7dnGStlNAT15+Y2QmqYPTTRZBCMgIjDSWO3IqFCrlIFFRFRPZ0hfwNNafrkkl1+
i9aZ3PcPdstd3A4KqhOXQhvRXUIrHwXiIytyfOrdFfij7uhO0ZEtT5eiaLNCsuVkEZAcELEs13Gy
MIUF+OOMJOQKyV0Ozk+H4MqBRZ5wjb+6wDAgj4U77UOGbJijw86OjfToC+n9ibGJfOVqlOnG/iTv
nuRbOeDpgLkrwQokE/xuRL4qjwGp21Q7H0jJ3PR4Hgu6hi2ocoU/SXygzBEom+rTnfW/t/p+QNei
TdHZsgZHddVDeu6Dsal6hDisIf1soQn8M3khKCnQOkNPIgbauKzaXmbwYTBl/zwIghFR1sP5x4Jy
jxgfd3uEYrIolf62l3Q3AMcirBSHgPJT8BlVc+307fPRWAYvCMcrPg3AUK4IPUiSrbj2CDZsH8qw
1LmHn/L22HY0FlrwqEJICAHmbwCTR3722hCVimTCgN8Juh2IqKjlfFEWiOUJL4c+SaPCwhVcCoCt
uVdhIW7+pxkC4kVIz0KcjtxmBOlnRgI4ZwWCpUao1IEgNq8mn/6KvURLVrYWa5oFdiQVaD7Y7IPX
FJ4rmPuml+c6aYLAV/yVRz+236HdVs3K7HFKZ/tHfhEzUz3HFIyzZmiDwKlsZeqQSXJUUHr9fTmD
cK3x/+psbuLgr5GW9OUOYDQhB7ZC1f8xIGoET7Jv55WRdnjrzkceJA/35czslMQqlL0q3BeJ5WT7
As5iQbunNnb4W7Jl1gatbRYz9S9W0Vi0CIa7TxtAMCXccaUZ2o3X6t4nWvKV2p5POtHpSOU12fWE
wdSRSCnYro+iLSO7X2MTICkuHMOzcDYHoBB6dWCTUesFDET/+NGxPE9OWI07VVqBskZfeUjqpsCw
bgjdNQ6S6klqGZzYc4/tofsDuNQRvED2y1bTzVqIaXL5dX4XyHC7PoU6iTCnIDGgTj1hJ391ah0p
jSURzfcf4WUrWvWIJ0DTp9qK88OeBo0eGJ933JgU3cRos+w2dWMlDwM5R2m4Kg9RYOXoUXOYyVCE
LCA3ZlzeiAc/enebJeVeCa2SNXYpbU5X547cY39eDQmBALSYYoOviSgwxqNmbGBadkgXntez/JYG
pw7t59Xv6fZCaz5ncXS4yDRx3g5eBX/M4F7I2a4vYqAQ/WG5uqr9Sz86bCC+UejejrsgCFInnMls
27KFX/Q+ko7E7F9VFXb7qxz2dsW1awmQzh+MOFTFK+aKSn2scT/Wt1uKh01/Anr4XZxZ+MNoaxDV
S5Zpf77nMNukzGUykAw2tB2lMKuDLocHMB4ksQu2LTZwpIbW9yZNIClVMW3g520HweLI8RzLvZ5L
NaltMwN4sioooZBWH6nZu2FjNlY4X2ACfh+Ypg3Cp0BBTfavLlMYRd0/sM0ohFCw0Gid1xX4m4/0
HZEbmZ1Z+q/01GYTt/U2l9CuApvKk2BG9czH/51JoC7t0geIQzWLIqyQpNwifzvSD0jpxDKqqkKp
mCZSO7ocf6mOMkx0q8wpl86Vb3kGCiD8IG0FUPSRaoz4cnVZWXGjTOwlUzuR+MIGwsEaPErlcttX
OSczxQ4DQD0SBfaqSNTsK9Yc76zUOHrgWfXT+GK9tum5srzXD3GPFT4KjRdcbZaTk6k5DuvEv6+v
7Vth2erzHjI+HdUjqS/UikEg/1BmbF/OGkp8SxbKvemH/ZyyIJoUcvBKrDVQ8U8NNH3dsIHGUVP0
ZqxNawpQKHAaOoNY58ChUTRAY2dG3aZOedwen2qBEvGidso0tsITXQ6ltGY5mvYDrWJwQyJXEdCy
CTx5Tng/tUmzFunkIjnAc8ccQvz5y9oiNwssAAHGRXDh4E2JdSTYW6iOUmT0wqWqceYXPBdVx5HE
aSyv8VGyEGZiCtP+bF/3U9cwBxZYnDq06aqE0i0Y0vuacsCrIpzTaLAJtai8RVHxNWcv8G/cpJc1
rTK/UNR2HAXGzPAGMX7QD0obdTrcJ2bG06u0fXYEKyuscEFXg7eNGpVjeg4eXH57NHygyB0su5p6
v1uFh4dyqcEGGtHrVPozBmEdcp8SaFGgJ+oQ86vMyaCkvrUktQEqdb57ZutRLX0+YVEdftFmZiGs
I5cvSLYhGe3K1ied8207Rqq8uAhPNyH99y+OU9l0JJ5PCAhPcVT89hc/pZ4ibLuj6/OxIpXOVhuU
dslInc7jE6KAa7cE8s2mqtMpNn5fTxid2hD0dvG3JzLLfcIAZK+UJxNjN+84EU0xcyK/iRrkjetp
DOVOOZmClmD4e9tuwCGJmFZhHuJ357ViY5oO2d+lu9VdLPhh6hHAzsqMtj0LF7iPXQEjJTVx2cfg
72ksAkr5Sqbx/H8pRrMkinsG8mi7FdBZMkIMwjJ5LR7QAUFBUcS8qbrmcPVeU7rd/lxa60LJjoT1
Jeu+5uS4CeM0ygpE3HDOeXmiWCWYHyBZhjpEAlznjOiKTWIs6HbSm7e6AIBDeRpWkLfHuWXIZNf2
N5aOrAB/XJvzdVRgwlrA2n0V+k6WZAqUDewBiG0rjamRxR3HmTZkw6OOpJRVHZH99DXDl8aYbOc9
ChxHIDCvjnnKyZflYuBRJWODPwpSbR2qNNxK/8VoDWI47ULHgu0ZVGOWwO2Hnb5hOE8tj1NGBLxy
/zSbugnEgbyd95X5thOmVpe0rY5rBMgVzuhrqyTxKbkXdlaaGrCbC2R/jccacqC3WKcq9rmmMjT3
qXihUVnC5abpZi4zhTWdrVVozWO6U9/3lmECUFTIH7GTrKmYeaIWSzO/yJnCEXXFUPW4YBY1RSaP
yF3smLjfMlSjVo2T1zKMejUgYmsIHBnq0NSshG2Yhd03YLyKcxnetnwWP9iaOz8cMHjKSQLyF3M2
sipYnuVwm/HbA19yuIkvoDwLo0J7CXzxVbHy56FKrIbjnaXZrTUUQQydpHOow51Z6f8e1KjtE4N3
48r/GXdIecYWuo3bdn4iiREnsnU6uoxBPF8Bl2EWxWXKcLWSWzto1HMxe1yrFzXwmWQB8qJeLu4l
KGg2rbpQYyJJ2bC3lWY4KNPkWL8dE+1IMkXwJNklo1hoaG8lv5HABpFgTZYov7x+ZXL+k0jf9PlR
h3D80/+vlNymt04RQhm+531cFq/k9351plHlBtEmHOs4AuHOniA7zX6SSygLHRjP1BKmj19oISHJ
OqwcXWKlVPfs39MRfd5FGyvOv5pHXe+AU0hzNwcT546O8XGQo3CYsM1pgnFqCsTeS1gmiLREkruD
SQJobS6Vv6OVRjIS9rX2/vqjUUs65XBsT8BUhSLTdZfLLC7jI1uTLrj9+mdlDkFdKT8API3H1eEe
GjFCCGM9sfEMkE5RUYsxvjBpikHQwj5OZR+0a4VQN87lzGnD3dYr5EAb0hj7OLNgUcS8gRjDlyMY
qgY6/Tyw7UvcDkCI66AH4HxdqTU1DKWH8PKjHkKdOyhWz6IyhE1PEFAousQU/hqFwkR1FmCwQZZZ
/iHDbyAq9LsYxo1N2WUUVALVwkW8O6Dbp/+7smpP6UlYxFaMmrAo//n9aA3zQRWW5WPmsFiQtPux
/6RKwZuC7L87fXCToLJgNXy533VgI5MnLnCbZF8sFQQRDQnin+KOWRL5HZtAcJq7XOib/P/4zRy7
3VNWTT8COX0iBzk4kyavb2dXnkx/ROXs+mopRFnP/tlyltxWaJoc9BvA3RQipZLs2anTFHGnuO0I
jI5UoA78o4VE/k32W1OxmxdvnwNaDe0fgFaOLeokmKCDueLpX8gkSGwkILSJGWw032Exw6i1vep3
zWK4C75AbVmILtfrsF7ie+Le149N3/Wpe0mf/e9HGRv03DC4uJqnHt/bLq0ykJ8f44THB597lCyV
lsKoZAe2loAEC0QH/vUZhoAmev61cglO/nQ+p0IdfCz3hDWGHXschJHz3TBf0dRMUyQHQ/5dzfWa
gGtTeNGVThLgwiKj8adiBxdiOvwh0fbFaoExnUGgB39w9F/sYnsBXV579EpsZ7WWEgzA3F+MvR4J
c2PK/2NA2duxAELEISHzu+AAGqZQxPJnHkBiv4TeMB+cErBJSn6qld1g0SR+MULi+zgPkGBD+yMk
h3WiVsz7oEjyFlvF9qHN7rfEeto6e4+Mh08wAPFSR7j0wax+N3CU+7YY1/+eMey1rzMO4oWnOOKm
pmGRrJHGkn68mfefoaanLs6EBa84I5M8G1dJL0k7bhDc95CSJWGQ18jH7HJa2fzhOCnRBtJGTXpY
gUocvQ1qAQKwDEIj7igXPDfgOHBASMCpoMDx8SNI72ZMuw1+r2O3s92GhDYK6pQAlRjkthXG55V+
5xJ/L7yAxezps+EfZDIzHKkHEirzn/+gwb8aGp8sguJMO53wBYGA39YLB2DIAmvRoCaJ7+xGTBOM
lwOt8kwsi55jBz8QPWGhN/1QDV9WCPZhhHaF7Gd9gfX03DXxdkjlD+dtQQ6cSmfx1rDyjP0Tiq7E
sKdD0tH9fYPSfRbwnaWG5TbC52s6ONeDfndLDelcBTFZc8bSLSpZV8ARYWSAH/fLSODHjEItNHjz
3N0hpa4LtPgThtp8NbsDrqsUg02dIADn2fznT2O1arPgwymNvO6TBfTbIR5tkxsSHe+DUkPxA9cF
mcw3CWvE1v9sdS+Me+/DAZHXxFyHZUOz9q61blZiDG4Ao2OlyE1rnFi1udooMvu3v6kGimLFnAuU
+jPDxq8pouwItXxPI/SqHnQNT5b1A8aPjyO1GreCLc4bca8ol4Mfu/+H9NcRFjPl9AQB0rw2Bsb3
x9YMzpoJSpb29I7sDKi5kH21D5ESYwGJEwenFrqzHSj/yxk0zdRP/QI+3Ec8cqX+BcZrb8Hy4ogc
9E69C64Vb8tx9N70Eb0e/86AaTaWmmFE2FyGIhQHNxvNu143Y1rn2UW/TgnpkgD2ef0lmgik/g+n
Vq5GuTf2EJFRacYp/PxBy3RVlS3I02q3TPd7Bsmu5PSVSVl+jHaVCig2LDbSVT3mOE3hs+Cip93+
4/YYPHxwarv+Xba8lTjuvTjohR0ZRViQdJ86kYFi4r+hnidNd6WxbLmuqBcbPX9rImzUTvtnBsRP
XnHX3A+zb7XCtKXTjinC0whIxcaJUxpWNyujTRJ+b3mKyaLD6XQT4Zo3SV3/DvjXo/CZLNz89cy2
Gsc1m15C4Idcm1B06M8M0uDWgF2pTd7gLZBftDpjacoOlUSN1UyYeYGkF1/ks7ELclII7dINhLlH
3o0BoMXpyPS7DsFaK7o5x3DxbWAhEP0u1CK7DHopBUek+roIfXENCrDKkgd7vuqcXW7zgQ56ovLi
PvxJYf6I+u5ckzB1RAFbcgP3LmcXjdX/iXVMCGLfw1Tp/ngRg1JCPC1en+/1IaitA8thPqzIvJ3a
wNhQx1JYEWAFcl6RwkFjC+LyvkJzPbzJNn1G+EKU4RBHJ91VRVcjNgqgu6YYeTc3qqI0YoJQi+xH
jNFNkunYplAKD2CFImAK0/mngCdPC696pf+JZuGXkwfPOYVQB2tp/tanAxegTi3PVI2qu6bAYBjp
mgxHtokwj+9uq3oSoYrKEq7Xj7+i99eGxTD2XRB0erUoh8kDkq70NMZP9xA3w3NXk0grSq4KkzYm
OpGocEmkSV/cAus3Dp/AeJLvjt3OTSfmXxMi+mctwtSFtrbEnQOoy9jJR0A48BAUs2BG/J4uKJjz
4TxdbVfo+I/wQV0NWTSRzUVKAsx16mUg84HJKqBvkfGP/+zGBzrEauU0Yvzsu6fLSZ5fFy8zZMd0
59QqPJDAMUi+GZkNepHdJveLbE3kjc4x5nsEJSsjKNZMwkyanYXWJ/uLJwJu14qyFKxrKqYK/ooi
EM4dd3mNkVBdquBmUw49GZphWmRT7VKOsFnJvi9PJGtQ/XU16cB0PGy7M7j7uNdgWEF3vLBcfc1y
oWCyNRy/o8KzmITAJCKNtUmkvUk/NZ9Z2C+7OxhecFF5duwGFr6m2SgqKnqHFGO0d17empDm7SaV
E3Y5eDr5QqFijwxAUyeDvYawHLjovOAPNqbKrxDDZ/ojjBVzsTU8t2HkB7G/X/Vu+SHfBX4B/DvY
cRCHAof/RmBWs3BAf9U7jMNZ8UVMD4Y+C5O7doONhsCQ1/KWa19X9NMloJ0G26mbBwvhQiY03/45
0mpvzJ3ZA4zDG3YEqhr6rg81DWSEo2TYJnWN2WFUYhJJ4Xr0L1AtkVHnASZVxjLEEYqLW7CwdIRy
lNh5NgBdO6Kt+e9LoIHdH3ZN8Vp1gyshoqzrsebu3Ip19CFFQjtdpc/FTqaQbIiwPQJ1bp6NPoI3
xB18K2TzEFDRpx3Q867ronrKQ0TZCZISLT2y4GR/iTadRLO4uRSAm4bWkdJLvf06Aer4yV4qdsci
YL1UIsv6RenRx1yC7SZUHfvpx7q0S+hQwMIEgQgvv5daCE+o4pclg9WQbJ/ukrcSaTAoDt47OfGh
sOqEtIX4ox16e1uDEbERXsl4b+wbo2VuwiJYf7TksDjJJdYrm6NSDbPL4R1wGcrD1PHnk4kyKrxb
GSJjG5izcobxCziI/7x5v7jX9JJEIpktWK30lwq12i/eMWMA2G6T00Xs1oWrdVe7yuutFCuGAJ1u
ys1S9PuP2OdP9wn61cd7KJ4X4zos93DGHrzo83UsCJWso7jrdoO+9zEzetlAnLIHlx00fIm/wt8i
Ub9O8SYG70AXvSYZq8YdNSJq3LWzyqN1c0i07+KGzeA5FSRxWMITNpfPKXyw7L3HcqefuhDPz/Fi
CQ3aT3/IdfLsqErHpVwbuHABiiRU8PVinOBhAZTMsz5PvCAkEOHfciSCnP1kxRxvOShif3F2UXn6
eHnWll3LaXe1DeWlRv769HGfkEdXregXB/K2JbKRWnmestqUAN2ZEH1hbjseCK/6ZLj8khdq3NqU
fLehWkIc3Z2EkH2mwhtfjP2erz68PwsJGO0RnXuOlmGOxmizjEzXMMr2+nWVL7AE5/34PSbm017c
0ZUtENjmMSJxrvAbM9KYRa/FWT+jlIHG9t8wpv1yjk/l8oDGQF+qdjx/cmcsM8S8CKO2Wq4Dxyjn
Ifu69VktxvLn7gc+s5vdJqj2GcCEoI3wtQD7n1ZARhiBjjMUGLuG36zz9nuSLuzwerK4bd8ggYRe
1Asvut3zEXKlpqweH7QLNLl0ou5GLNhPt40AvHhpf8oGhxyuJpb7NNESGir6YV7aMDZQ3HeJ3Bgj
+b+X2sARrAWbsRl1eNpPvyWJ2AmgX3uog6wLr8Wbn9QuhpPS8U0s0NG4a0Tsj2e4+YqMaeRuK0eA
lMR9SGU7YMaBDcrsmCxaditNHJBmSzD99ZIfFWmYMWWTiDDUln5Y+ejPZPY/LDvKvoiyONNuCsEX
RiS3oZrFhxzPyzApi2+mV0JcMqY/a4RA9xUw0XZp3begvnZKIhqAjBVIi/ZAZkP4seGb0Hgs2Eac
ac0D+GMx32bgaejOJpo/URtHKWv3Klw0vj3XqpMiciwHMnIXlpp5xnFkBEC/cbUYbT7qZmkdz7hO
y1XHFu3xSSI7rg93v6FsdQ8eAhhMf7SW5Pc2zK9BmlJNZP9f7fAIuEd5xXjJ7wEEJEYxtJSmY+QD
xpRYbq0uSmuzdyZy8AGouiqoFZaunHfcVIIOom8k1CXABijBxn34w9adVwxlfi9jpibHXHgZ/zzX
9tToT5rcYGiQKlHSv9QMVeTxvbp7bRPpY5dWyKLIFoI2pXTNeChoG3w/4x6wBDo3Ow2qYNVt72pi
hGDpVdxrut6rEx4wS52Lv5DAvnEancmi3Prg7ByptaF1+8Kydtt+CmmM1lTNA18zAXfwoTe1Zf8E
JsbQ2f6t5pxOvwQFIuSNV+beICEH2GWilSXP+PhWLSBrvI/GC6pIKQkJWEBkb5eWdPs9azhzPSvH
+pkQ5ZFCM0N55Ri3hjl4x0vIrzlN8TTjAVOhGDyghA/uXCIyIiUmcbcink7q9lL/pSy+Hf3mjPaA
1IUjRtcnVUENQy+wfB3glyX0KC/onpWdWY2U+0NAex0oqzORo034/O8am/UKInJLN2dFwwDghUjL
88Xph4niyzgkfYO/3WGNTTHkIeh1XtkMi4S1MKwRuQo13JA723hgHl8mCjJmHT2wXVAm3hcdBTq1
nScJkSOuNrKBFY+3fotP+QJEvqKp5Jaycz9U8JuZCpk9HYgYPpozagIqMtl0gHHXkQymg5sIXHZW
/nSER6UKuIx1zS3e6/B1FqR5V3tCzU+ihJ7o/EdC2yj2yrxeDKDtEl0jaThAjAebBsDpGuRkEQhv
wlN2txeq5JMHenCcEIZE8wEfgdura79pG5jzLBRrU/nYeb9qaiqUQj14soMxzO3gRlyXs/bepcLG
VUEqWtx1JUmY3xl2or5FoNujzDjlrPjylDOpyB95qdMssEMogBfpnNgQelECHELwAQg2nGEgbzxW
VdF5L1KCgLmWIAGfhQcG/BYvWthacwZ472yK6gTFBsTyBEt79IompOWsiS6o4cCFMd1x0HzE0kTS
c33mpWrX+4evxnxbdDPlz2AYbKveftf94kYHmgJWvJPn9VcyGohdmGXlWTlpjBLJKWhVJE0jVEa4
AakR9Q0k2LjsWAIV17CP6C609FHZtSFcV35dv4I8Djfk4mX6V7M3tcYkkv0EZ1HN9QwCiLLY6hGB
y4/WQLKFuQraqnsetzf8vqw0tfcnV0p7yAOao6LG5oFWc3VFcMTf/5rjVpza/lpr3ld0azzviLwD
4PoUEFvwEql13tqdeqEmY333vxyVZLDwRvO/O8Wr9BqKDziIP+23dxXm22rhmLtX59s2igsHQslr
1U9JeAtQq3+KR/NuofamsP31KiBM0PCfSs4QGQnRWyn2BW7GFBVyVZCKOO2f4MWTH5wrebz/36Id
c5F8Os4DiTcE0P1BDlLrYA8jWYcc5Cfl/7cZxG0hlMqE0rKiGnMgw5Ff0XV4zgHMJMbmGZMmM13/
cWdKnvjq8gBXnAhxQe44pqkEMsQS0R5+wfZLO0CowcOwOpSJuS1jWKa92PkHlHDGbYbF5FL3hTDW
3Fn4Ti4zc9d1ZCzlKuu3QJYz+hOtYtOX6WcisywEzf0aChBtppf/wZ3LpnfTFvhPBwEnxYVgNxPT
bW7TuyzbWaWqVdFPUboygORN5cMinEsZMMsYBgDXQw147ONoeOOowy5iCQq5q+ZqgyVRUoPhjicB
RIqVuOG8Ko4SNWbwWBp10j1wNHBv20/D9QAak5Yc2DTrDzjGPm7TsJFWTY1uRWGcWiMh5D7lPF5Z
KxGIn3L7Z19vErz2qBjxSMrF9HksPKJzhCwx+pzCasqM3LoSa8QitIy6SiCsSoyrL4ydUrfbwGRb
hbekgmp6fmVK4imU+QxTcQEEeajnLPBlpqsUb4CRlbfXxL39wFm5HGCZPasfpZBL1btLGH4gMah4
70Bel0U4E1JXr3cODY6AiBvnoUoDg4IGJtSsMKRHmwRSJdShtGN3R8sqzbYU0OmOQWCM6mNCxcye
HC1hZkI2j172Sr+dI/0PYnSgBwxGEQDY7+AB5q5WKz92LZsQxQLakEKBCH1SCJHyD64AmuKX5Xmb
zfhR2oYfHG/IWTa2punjnGrLC0JBN9rADFhfuLFyIiwmSPkOLyoOlnD1EHfZh27OExucPj5Vc6bH
c1H6/WNY6oCrBM+xI4YqbAmguhESU4aRSLSxoB0FRsl5hPcHG2K+4kK0S2Z8S+8JpKOBcQjvfa1U
ddDyT8pxrkxnWdAWBDZ0iKASlTJ/KSmM2Qxr4GO1k7nyyMDQpygoakimgIERmCrZ4Ezm/mKmQGLm
opUgWG8NLMMYj15JtBntfJ2chV1l9T2t3D3loRntWQQ0D/d8o4wWuVIUTX+EVz2kBNNm1J6Q7y0g
qZLeWbWo8twYoJtmMTGYcWbE0JR+All4S8+WDnNRu8h6xN+IuBhViz5lQw29R4PXYnqkkxquQaRX
rorp+wyY/bQ59U2BcbmtPxqC2BI2xjwCoefPoG2+D8lm+AH+2a6tQg6xgaTyV3ZLsdNJD3QS/uYV
cfYx08BWAVHDRTA0b8pOpkG9eHwDaLZ0H8B1vO1jMnpUgjsnj4zNVeQ9b/6aZUa8OtiIdERwqSWh
PusQ2gG9WKl9qZRNqweBw2XSawFVnHXS6x+/p1tOu1xHu2VVELKBUG6Zfron817mdZGXGO+yVnLw
hAcV6eD8FP/C5NTrAY5p0g6zJOVEUXk+BoYuiY4pg0RaA3ogj8qf2Rgr392b2J6opfBs6Z2IGWkh
8xUmMob/O7E6Mu/cVgfTz8iEVnGxuYRZNvHyq8gvqNtXme70cSC0oxZ7M7rocD0RR/ROGSQqTooJ
O1OYJ360wLKo5rsoQfziOHP4/ClTeqQ8digZKEioz9d94tdiCh0N9jgqdIxFlPrMvdZJbFHLPfhz
IB2gfZJTSM0jMmL2Idm1iKiO173VNsQmbf6pB/pb4IQcM46vlw+hsoNG6pwbnDQwuaxE3qeDS3/B
OCRmMou8bIFAOCWdHBEb61eqps798ShJl090N9p1B89Dvs+IOAa/YLQ2T2HCEysC+mGEX0+xYdxN
VG5SGE07m7GlBOD/J99CZBiJesOiFs0QbIQhoTVl74w67FkqtUXIzQUIvX5hBASo8fJvMMKkcVmB
j+9BeuToqb4D2bKbvNfL29clPmVyhZnOt4Wv7XU8lx49tg95xqpFw4SliVAqeuZvMoCeN4TVGbDq
SElicezWMw+1U/aFVQapAd6vqGxvMMhn1SengSz2YSs+z9X7R2Mj/EfcYZDmioXdzobKFUWG0Xcu
Yev8ODbgtS9aezK/3WFFXnj+qHjxsBm+BwfjfGgpnEwZVTtumJyCZ9cy6Fy+9U4EOlODjFQGAI9/
Bhlez3dSzEbNaFsNXAaPu5OOIviO2Xdn2mdFkt9/m2pR9NgCeVFuIPjvZFfYcoL3haVZEZ/+Mckw
u6lUoc1dwzC81BkMk6xADJcsGvo5T3RTndEDGnqqbEtwviSNFcD2273fSqk9rMSXWW4R8roj/+RU
NVVDGn6U6OVMekc52ixoSfEHtCDrU2xBwl5zR9c8ed1zRRMQwM2n0EYtfeLh5SMc/TYImCVf158l
KeowwD5WYJ0WdThKZvnNed4AA9b42JyLxlDr+ecvYEPQBPoF3qE8pEA6asYKfE2uG8H1+cWSx+BF
Vc7wQKxJW4pJkM0vli9k8KQsrLMzFzlp22ScnwvZ2AMqVJyjqDj6SwwDkxV4lc8nM+LmTeUxulGT
Gghj0nQnFJsNfJeM+mbWvUdIN1MsPezF72ubSXM8CHTBKbO+BVlbgO2xUtKDUVieuPupOTPXflDP
uP7fyNF/Qw6Enc0ti8ik8QmUUk4Up6uAzbS5232SOcpy1JCE+46W2GepawaK4sWK9KQtu4X14E5j
H4XSPtRd8bCEv3o8NtoKSYpno+0nO2aWNQQr6y7nhFjOQBYolnQ7GscKvDlwKOULostqemJjw+dl
ScBC5TKceyNPX5Qdwic5HWp7C2Wv5RykUHKw5ABbCM9Ik/ivAzyjnxdeZAw+o8gzetGna4L4kjnU
87WVmgYSK8BTe1crw04sXI9Ue02yFTJ4EGNvAwplHYwUjv+X9QCl9t9zHBBFux5YCgMPZLgO4fh+
Ae0OtqRpUTz0GmBJemH2q1bRiYX3HvklB1rd86KZXApr8oJI+dJFbUABmZ0wW9MmbbWBuDs7X4xK
iEdJuexKK9fZzeVYW9/OO19EekWJ3u713+2elTif/CkMX6wFKHoRq8B42ZOD/u2P0KCvOVqCwXOS
lOQGRcTN38xgiR7l5sgo/CcEmplAOo+N5Xm8puCW7Qaphboym89S9dtoOJ2A2m1LjcvJ3au0R8Xs
M756jJcJOVU0kSqA84LUxnLwaKZuppGGcMDC3hNXNmeSzXNS7N4+fNicQky/wa4ih+u0GLKNLZp+
qFI5bdvOQbRXrj3srcMHjD7C20t/dVMr63ntFagQg7JNlZRjvv8AF9tPHTWXWgUudhvSGIBTzHKZ
oYw3diMzyXqXw2YtKQi6cs26WfW5wvt/XLwHh0zO08sEqE1Ee3TApAeJuNyk7v5trWxpDmOYWLs6
OtcTUKKFqyUeuRzechMeTpFlgz5UBh26rh8bEhx0D7xh1DI9ItQ0oeCaPoTf+3FJ4+CfdUJqOvH+
RxUBFf4XZyogoa1lnWD8KpxeOBlPH5IWImkHW4qxB2VKUiDw1NZybUOdXhdeeYSPiVJahN+NViLJ
EqgdM+Ol1BzlGL1yMc/f5KjyDJLLYL6cFUwmMFlXfou4W5JcuoSMx8IyC1jKxLPp/zj5FGnXrOcU
UgLv9sPIQlg/8EirqCFWXZzBYbnICDsV/1kJav3EJKC3+avjRC4eLU7iHJ7IUIeitKmx6gkE/gs4
DyCMy2+7uhJumXWF/jLvGjsMt0Omzn4Ib3+jK/FpVjY0E+xWlO1KwMp1tUwXibd1GDGfsMmW6ilt
hGVpnd2XV6fj7vUF/sYNWYWzhnoResZkhLmuemFssV6QXWx2RVIhqU/WJTfhK/WhZ1OFK+Ny0dM7
+BopJmPUrdydqegJ/G2yqqd3dSUANLAia/7zMRq+fvdCOYLLEoOLSgf04Hg+TU2AWfhts5fREdaz
aGfFlRVGzPYb0KtcPZw9ySIdhdTkiWEWDCHaHz2byZH+lKCqC0arSLxwsl8vLmcQfCka73jreFhR
C6JxqrclSi97CcUswL3CSZ/UxDPITsUhcOnj/hrn4Z5x7KNGr5M3DEUmxRHu/KiKMPd0IgZ+KeX7
DB68UP0OzYE87kubAH7nAHZ19xgw5u/hoeSdooB2GoUGWdNuoeZ3mjbxn0zNlhzqFPhz7dvdJYEI
L5uBza5/B621CciuYZDLiKreueOo5nXlSaqsMcaRWUrzOTbpgfZeQ0CEwEOMF4EGiXN2NGtCDXfM
vSBP8vKANs1iYv5oO7Egsx7XiRyMIgsgKgaicrluydJszwrwqrHcM7Jd72HFlBkV5DR8DCQZzfWG
Uki/c5vS8AnyzlmLrRIYXApyTH6AJOZNbO0OZD36lV2znPixPlxUzKIJdmJJjLIiIB2jC6JzDCd5
nALMIJg8z7V0oxsn6PLMqsaqD2yb2DGc6PD0FeahnymlX5v2Je/dGtlB5zZIy/jdLdFabvfWKD8o
AJL8W+gNq5xM3CLyKANu4gfYElJ+BNX73tTu5nMFVNih7XT5BBndyRjqquSFbQrXORwXOQAMx2/a
SWf51OeduWsmC+DydvpgscLwpZrRLt5GCpNp9zR12meEcoNxKkUvoN5lDwyY0n2gdbfDb7XQWi0+
7+HoGKCSFFljlKyRPa1hqKCrZsK0lnol5ggSKBskTkoaO+FJESLNRb8++LJV+aqSfFrXBkFuInUJ
Rgw3KOT0jMke/xQvv0BNmGxt3B39f2/83/wkj6UU5rGAKCU/D0ggbAWlnhI+pBvkEvdM/gvwaslD
Q+H4pqvjrfZt1UXOocxEJTAB+AIh6sWDQZQ2lw9gmZexZxUQqJ08gqNtw9v9jl4P5EA+Cvm9qt2I
UWqa6XKl850pqOfmgy3AMvDf/J40fJN8q4n5kwjTjlQEZCVBv5eEpS57Zc3H+PkIyfk7yEuFWeS2
ZzEiBmg/tCYoOOiLcHqZ34FfMoA3C7iUJfOQG+MliW5YL/2O6PVCFfPAyFC1p56X6nKajVq7lv8f
7JaWdNAE25cRun1ke2MA3BzHbQ9TV/oUDLezwUb/8Ufl5JMBEdhQtEVSv82xcqngIdh91Ph7uzys
fcJhzetL9OZUlFYtn59S1wLwuHY7iUoNnzE36CjdvKW5z2XD1YGNKZ1XMld9dIDZti7x/2e7d2cc
VvfJ77ShxnzG5ZsWXechYaVDtac1lZG05CsMEvRtB3N2wBIFjl6XMBx0XhCyIq0kpCnuo3PmLiYl
Gd/T/u4LI6s2o/OUfaGLphSmLYwM3rbTzo2Q3h3SpdCTFML4WbH4nPtXHMigCe1SlWP1hMuNU1n4
5UVV6FGn1b4sng92ncQRK0Gmc0t8c6BZtYnueFwi37K3l7XQddIm6sWU/3cv0x6+P/NL9sm221ko
TRyQAQD/9EAZWe81sBo8A/T5x5nIap0F/A/rX5CWkSyG6u9lmOri/Dripj0yPH4GJ860K957ClRu
b4ptVnhg+R2Ypp3DoicwTg4kMbe1saAcPQPS6dA9XFKD26zAyEvvkG8MeOK0b4OZrgu8RT8rK3/7
JLs3TmjD3H3nDxSfmQyiybl2A8pZYGTnH1RgztpjE8zxNDAQ4bUd/OXqo2VpMaLchRMF3aPDxKeY
4tmL3LMkxqRasODhL3Yy9iPw40YkrcqnYc94TnHbJ/rA/+e/khsbq6lj07cDjVm+6mCgQI10br7o
r9r8X3zD1CvCS+au9cL2U5aHprLn2nTwtxsKXDQikoJoVvTEVS6T7/GEssoU8bqdc/WEKVGflV86
+TCicZx55EhySpijZz5/wzoRSaN+lgBWbbfF6qYh1gRkYoHEw+7shGBFcBaCe8AB5S7UD6Dh51Ag
o/UHPDmdvKE/1cCE9MnRHPj37TLXylofW6QF2RPCQXkCpsPG/ycEyEUCndlCpTDNoz2UQdAdJSEd
FmohOqRrdqrpztgws65Wq305PSxqVRFHfmErZRY4Y4AMTTxpM1gPdchUXOuUKMNofJ5jLxcSUJPk
mgnX1u7GItrzr4s/QIZOKQurUkUIyDILctOAUR25FKnkQmU7Q5Fn4iHbC/D7qQVDi+AbBTxLyeM+
i9L95sphBcrWZ1zvjxYn+OgA+0+7LKHGkSvNceRxKjhRo7xCTdw2ED/7Aj4MI82zEmawtHI5QpTB
5Rhor43CG6qn2T7Gcz2TRZvHkIHUVy6Ajfut/ShRtVOiagR7hUqKhrjJUlrZ28j85qtQLYCLqBX+
tKKznttCKMmAn9lKnP6sz3tz2t4gYl+tCgzinbAIRhKCPLcdvScRClJekymzeNwcKgbUG10BRXVw
Tu98GWZ+C0sIDfPY565y1l+ogMShJ/gi8E7xeBgsfVmzz7nZJU7PgJVAuT/MXegfsjxEL8gIYbCd
ABMVYP4oBbSMTEROPr7jSHw61ACQv5i8gq5FMavgH2nj1Zw9FFo16qOPb8yoXxW/jZF6fmO9TmD7
MsZT772LMbFT9WTkqv1LkVDVIbs+QQjI4OIpyObVApgGAgHXTW+JBhKP37B03sz5QJI2Ln5msBZ0
L/D+82FxmCuU3SukZvbQtXuZEfFUGWPSiLu1VCDlFTSXMbM/Bp+8C6MTl1gm4JoYjl2yyh/QGtAc
eQGDSi6ciq13qaO0gGSAZrdHY0QPn7D0Mp2GywFs4acyiYHLcjY0Xab4E9G/6q69FTvR85ZPpDyb
kRKKrg9k0/hOu5PpvNAjGJQ5ksZrdxaZmjEv+p25vkI/nKMeg3upOoPHFDtAbRfMfqEvq2u8TjD+
kuW6XwdeXHGEE7BWsOVtbmP6A6wnWO6BH7nsJXsP1MuxfMXyCAbiToS92cKKoMUhKwst4eflpfGy
z7C9mvrsDY1dHwZ2COXTZr6aqdWx0g5lJMqFre36ZQpBhuCULn/UEN9o3GAhThlhvJYQ+eEt/ub4
I2PXlwgGWBSZTc5bsZNRzuAaSj7ZPECQcvdCQBv9kZG0Sf4PVzHo6jFU2Gtyre1O8k7S0dUIiSs9
cGQVUR1Djw8MX8Fz+E9ohW+Sb1eLWzvjCuQsleL+eTkMxt7afMU5Df3O4FHtMShEmTmJ5wzJkHeg
aYG+Z21Gv8OXmR1Ie0sPgc+ppIvbSQvAsiO+4E2F3ygFuWsRhWfuKCgmPizuYasNJYVUU3+BTDyt
rEcrgUPHu424t9D8SmG6svdjQAAcihmPjGzZFY0JeVVw8B5njcLH1LFdcYtSPkvps1Z2bsrTy04o
nokPc5pccdqmb64eKeEZwJzhDxo8CpBvW45mB7ZPRvLqeokqFm8bToD2yEPPXgmNviKIwM/rSsVr
ArX+YJpI2W8zMIsfaFIaJ7gaE+Dm8m7Ph9VEDfFddO8aftaOmsJHgX+lDG/ETlPZ9rE/RTsuuRBz
XOjwOLO84yTKiE4h7xOSusWWh/daBF5jzxY4E5586lhs+9asD1aE7tNPp3S7Gxw6qK1WNg/lAZ8z
y+Jli9nxVyCZ2YVkHXuRlB+JAk4c99Fw0I7HbDU5RfhxkaxUV9+kmRzQSC4KwkdsRK9QVKedgYCd
fun3TRC9dbIi8aptSPHmpsK3KTWN6Tk7NxQLbITTGioJafvblhBmU3Lx/T6/Gj9oD95NGGxZXeku
eiX+3NkCmrRNPfxLmMY//iX5vQ+rh01EImXlooYwx3AmmBwl7clCvmhCte5ZsitDiwTV5JD9zax3
eg/Vdvs7u8h+8SNBBTIGjhb7eApFsCU9LZfBKz5pg//X5Y12wbDU3LKiM5Z2/Mr59hO+HKVOYVGV
ZSVFGGJ71dFEWe9/7WssS3acA/8XzbUf4cmc4UrD9I/1ZF8Nz6Aqgfz6Yi25i+9hZ9VPsem+0LNZ
jblQNgybiez75P6jCFCrFQTY/oVsfA6ihoGJkJPITwIiQUCxee+phCEdoHL1UM6WWynETHO9fKjp
Oz1oTZxCAciicQEkm0t43lCGwnPvJq/RdlkohVr1zjjd0XifAfFhIT+sfg78hiR4I181QORlRoWL
Xrt6eULRgySnCWrFoarVGJgUMd2/adLKFixrmX8i7gQSLUP6AI9NTQWpkLFAVqH0DggM+XZeX6cB
GCA9rJeZTc4W7nZBzL0wGkLolOForXgwtP9bogwriEDanvFbnAxUvSRqx1rIZnasAsOfBPaJGqE5
GVXj92zBTFxuSi3YhfCwzrZYedo5IEaD/1vc3iTEXaC8e0+qKK3o+izX8gmRLm2037PRqjloDusR
peLFucAFF5TVBd/HfSIyVUgmaO1M4B+le1AOSJjHckY5vC0dTQlCuXx2ZU8aSpwNiFnvgujCKZU4
9eAS1GmqzeLRrZcA+SkrbSzH9esJn4f2JYXWR10uCgJpiWgCRk0qPMXqj1KSz2UISBhhl/wBkIst
8zNzVaFADInLuBL95JYKfGKqUWkYv7tWGXYEk2Py1+fVbt7Iy1gQnC5t4ggs8ZrUokvYpc6o0VBv
Xg0oxW0Eq0+mbyr07loq1jNhshhpN3WQqQigvPZBIEjHcIGZqZoZzNAeWJ4IpGX09U4JttAoBxPy
UvO5KIA+qEW4F6iMxkoQAf0EcWhoO0nNWCBW+K/sPunMGUKwhxbQZuUxzUAK+Slmr8ltKOpNjVdb
Hdb612mgO5chjZbTNoipb6pA+3/w3Yr1ynDUBpIPmMv6UaAcfDi6NM4OShtq9k2DiBsNtg3EY3nl
00oimZYH+yz/hZfAP7DLccXVl7JHRsARuhJE3F2jzgY8+M04sEFrkPfKWEScNppx8iLbgK4fc640
ns/gEnDKhgOFhOegTHqAxeRamR4df1mlKmPW3l0/T8t8Df2c/RDfA0gzw8lDIYyYrqfIYEn46f/3
vQg2J/xRGm7li+gqjG2hFvKBdxMPhCJTLdSqo9Xn20bvkeCLJ9p36F8zQDAhTiLki0Y6UI6fyQ8Q
NOV2a42sgzyJ3PrVB1XA6xr81Ey7BF991FnFwCCVveLwn8shcBEObRsWWGsmxHROzzplgFl251BK
Ys7JnXLKNXekbQC0uPydIrX4dnzopmtzOdb2K5xs/kbfC+kSkC4JQlDjij5Hj995Tl+02yS1osz8
F43X06awVlKyJNH8YZtWS/Wwe4RdW26F6fUxlEteX2X5K2nzQPSFL8KYp1pHwbkOYLSL/YTJ4mEO
G5GZphNwb5ThnQh/HAv/QK1Hm1E7tFBQjnmTC4VX6tAuGLUgREyK1wJ4Hj57LruQ5WypbKnhISyt
eqNI8ZdnWkeUIMvdwY0KzSjtMnWzLXcsP8NsZOTcl53P7Ghh932rgJc0MzcXkEAwzqWbV2msy9zW
MK9ElVhUZBJ0V/N8/x0Z1WMhI1hWNGmwIi4XqKJ7OwWiZDfLIIp4jsYIoqvjl/mr5r4sWdx3lGl7
ilXyXwelQUCgGd0Rn/5NpJSUQRS4+tH8b1kwcUi2NxaoIjbLAOIpUCbOTnKJeZaTEh1h4u9mDOjy
M7yxf1d5ODySQFDA+oSTqFX1QCEzena/Wm/vUZHC2IHWnLwae4/EBULg+VR3YWxkNfpBOLnCv/HG
6d/BcgYuPvPW1GQ8S+mG2CaWZZpwCntEFjtzXDacXHNRawV7nURkY/nQAwzmoCGL658MCoGxKCZY
DwJEN+JpSZ0u3NeBQFBWa/lkPthiwnvqJnIB2gRQ/r54iyO2u75FK4K65kpxnF39bK7N8pIDzWMs
E4sHXZiBxXmrnIorpaNuISfu9jF7KSikqXd9MrhOTBth92n54n7mM3vSo4mzq1kOvfV2rNrbXw7c
I1n98yhI/H4kfBALSnpYFe1i9QAZ9YsaZ886BMTfrcQSIa39qE9Z6nThVMCkrZMNuQTIh7jR9iDJ
bGy5wodmKAvC1TfTEs9IuhSFkaFBvwFu5IWuXdfN3Af2uzrQmXLFmw5mM+wvY0Zsvq1HEznH//uT
HRV8f52VEkLjRGIiMBfYxw1k4rqLiA9k/JkcKj1Yys2UA0mW3BLwVUYFWtccrpE7a4Cy22twBLYC
EmoZhi8H+emE2KovVsek8GJADW/iXrbuE43hdn2zW/iwROch+ZsdYPCwIfv0jbwrYl1pJcjuN7QR
QF61B4eFaOk7HAJyIb8Po0H4aGHVkfg+pIK3zkjod3B1p8SLqD0vkPiNKQ578Fv0rz24L4M3e3J4
GBHbgVdRDjeT+TROIYH/hgiB1zovC53+iio5Wp7VkSzOFLhMZeXO4QrT/He5kh6hk9XyKdTMntcD
Z/qa4Ra284cZEBkvnZ0omQT62s2qxdS1uLr7HFGfceUTOhqOHZWaXqwXKrZHHjNDLdessfzdzYfO
/EhpxrxTxkmfUZfAZdnSztwJsu1M6aHHx0fASP+TiBasAxS48FH3+VljLkr0uYrPq+Es7yADqP+8
ICLrGsmlFiWUIqVdkW9fGXbUjdDeyhpMCXIUrIoDZVUMZpIFuQEYamTgNSz7AO8MVXx989GNxoC8
NC1WtgdqxXmZ/+vG6PSQo7PBC/khB1zMxPHJZ5+zKsIosyAmBVPXo0kLY2nsoN3aALukkLWCqWc+
MlTZOzJeU/Wif7k0idpzMZdyHKXNKZOdI+1ZmZmzzOp2imsa0nETDcqkVo5DOurAo7Nk3PVMJzbU
Ngv+aPRD6aQtobigs++ZXloW5Lz02SVx8bfZ7JNUWWAAnJ1doWLyEgo2LiPd85YjP99tUbif3naE
DdlWst8ID9sqocuEvYjm27k4KnB8g0i7SZjG+6UsJu2UM/idxWw2jbKrkOMvpViy998IjWvif14T
W26C9/IE5cJNXoRqzDLhz9ztWqR/YS3Qz43zacRyOA3DnVBifMK+R0q8Xbu4wJiJ8GPoJ4rlO/kj
F6h2qeSdIQEK0CuBIP6vzDjJJYB3F/FGIY1of9rLBs1Ex3SMJcNMUkgl9b5GyGLArBtiLu3UNLoo
7oEuWv8kWl/SH4MxWVGRt1Mfp85KPqij8qPx9WSvQtfV8d5SldIiivzLuGq8aBF1cTT0+C7bdPHZ
1oTi5N/fvdthAVVj2evX1Qe2sKSP/hbxPxZyt/a2nNkeR78zi9HMl6L8iINRua9+HF3pNED/NgoS
LiQy61ayxQ0e4YgwwFBBRnbt2E3WHpAragugISBMi7MrV3u860OEZEtyMLdDLWgqnGAvJazDdIfi
b/a+L6ENM3YZfNKrbYqkLUgyUhe3dWutbew3bJIu8qmMORvgGzV5rxnmFQXEWWwi4S64+obnWlyL
ieq9Q8kAYZjNCAk81k4xFoiDTUs/BPABdXVR7FTK+S4By0bAQfw7eBb0NCH8o+fXZuQMvnPRLOQg
oJEBcNMdWE3unTYPxbQLrznWKKzC1kDtudDif5RL/k/Z6WSAVwdX7StClkwb0CI4BiGao/iPNzZa
wfKyDIuK3asM048swPUXZPIJdXPbPvM3xAG0vGCLJgqyCtkiuMovqI/Toa7jDeYXTFOjPhxOY5A/
DVfcUw5MTZkwNonh6v5LVq+JlvGaKrpU789lAPRpUMDeEchsNfUEGNb+Yk9mjS1l0s1WKFCh7a6F
OQRf1s1i2MFNLbfWWNpa3tRm0bM9HmuQG2OjfocqqojVC+kwQDszoXZZ4DMd5NNxh3oDkyiRCRoP
t4ug7+OiEEP4VS4zdl+HadHGRLUYVkGk+dDZoyHrrPndEDNaKXZ5cMKHYuoQJiC+sMjn256i4aUv
POf/68ovk3/3fkaePEvZrteeIAr0lKLx5e53F6kb4yPbd2YHX01cnzfN/4w0gdKYg87/cSw5z69J
KsE9ynCVnYJd2gis+I0mrbAyamY5BwFR0wjpFZa8iRos9o3dhJ9LYkZ4ra2YEkbPwbLWaHoeSgK6
lxcRE1Sr8F5oKTZR9ir3l7ZEPl748qEEsDQ3rXA8rQ/xx5oIP7x43Y5Zngs2g3bWDAI4F7sn+miz
+xRMKthTLXp41daiscAOtWPHUZpvSGB0NmQoSIN5E1F9DGwk+KJxB1GJfqidokcqQIv5d13DjRFF
ecS7JssGME7a/ATclek9uOdztxHVUPMdKAmb2NKU2lJ101Bsl3ZzS5Q1XtTcMsvfMJvM3TpL7o9O
6BxsqPuLIb0DsYgUqDN85e5uazn1MdfeOanUdsgyFh1tmeqSTOw/r0dz7o5F1cCgcFJs5v1fiYzr
/IjT+IjF5p6gQCqlzja4N3U7DQw2qQC1ZmUXbZJmF646+yh+/E9ie4uHMwjulGf3vi1BQmU5mh3B
O/Jv6bhFCoExXwYdcnECdKm6gO8xtzwnogLoX1PjdVYC31k01hvXV/r0DzRu0WJGd8QGCBu8vxV5
6OKpY9hX4vUtwKRAYPCE/DWAkOa7wuowFNfOGE6d0omnh/TY59rf/tmmTrAaVuiZ4DCLFXPdC8/3
vaglIrewhYnLXUl+ulFhXSuoTlyRrjwLulMMyLWxq7wbtP2KFIbeoihFCOL9LtSLaSp6GXvoKV2t
Qx39i+QjT277x+y6BcNtG5RV25S/BB7jCWVav3P3Q1MY7i+BV1vRpKB5tq78IJdeuK9CS/5BbRSG
2dKfArNNIM82qQt9BumkTAAMjXLGasfg4hEQFZZ8rzFeSmi08rahphE6AV0Vp6C+UiNqEDxiMwux
DkHvTuPOjP46nLnxOmzjWvY8IHEtlQFyt6+fKVCYH2x+4ogyHey48r7Tv0V3mIrgYk73zcqdy2Jg
ETizee9LfJJVxymNwoBuNvRfDm8TcHsIoqBL6+OArCD4h3PVrfO3Lo38nGiN3fNcGpyjFiKRrkLQ
4M2kNlVyhlgf4CoKDmXZ3PZaOi62Y/iiOQPgAEEVLryTOireWBd5WXxN4S1OJDIpIR4gHd0qxEVP
Md2eVFkYHhPd9EGr1zGnfm8tI5EmnIW08id4qaAlIqvwwlmM2I2/o9MXhU14cKDIXaiWR36xQ0Pb
N8VcRzA11a8mMYGJPYrl9WnSwnCOllvu2tapZJ+6WRg5lUMqyANvlbGOYbmteynrtQ2QlNqKzju7
PwHlVkHHBrhaLit0uGpcQch/AQkyUgwZ9S5g0dVr2Sk1dgmtZnxVcumL9kk3L568R8ZIxr2fE+xB
LZtVAbdfE8JuBlHjz1k2cX7XtEhKiY2vHYGp3gc3OpN8KuhRUQMZtIp/AOWZOSzK9vaIC2vMMvFf
IdR+vfNc+aTEDIO9m2kOVp8/iUyEhk5Sa1IlGUTgJGJo8Pzm1c4DRZaI5L7kFoiTDM6ylEJtRuuy
F2Xi2pZFX1ugpkmya1siPdwCrgJUUyh18lywYaKHa4hMAbOa+9vOJGi16k5qX8qx6qfZgi6iCsqv
qS0eOIPsG6LfFftnMaUvL6bnUQIu8twffSnWUD0C3v0MuF857NbDnaFNQDng9PI7ibyJWONdnbkl
1ySeMeI3QHxdVjgLBCeVSxu16zWg6EhygxSMyll54oBBxWnwrCS9rL8ko7z4M/hNePs7f+DlqNv7
EotLs8NRt39OMGaZyEZZMw2Lhp6BZGPofS3GOPnSYeGygo5f7NRmVM5qa9XTNEtsRaQAcHDNBkVc
3U+Kdp3SmijnDooMoMFr09VSCz2yl0F59sx9+drVYEEHkJTZjZYiGf5BYBd4yzldYHmIbZg7VQma
1s87VEt6N1eiVKlP03oE6ifYcTgYRKOGre3E7bktHPoU+doeNjDJ2SlmY6Kjjhr4lWKSZgCFISqI
7ZiP0fELLQukNnIiAnwI9Pf1gUDxnrbEA3HYlQh6X/rBtlvXjrOV4uhUAd9AM1eXmSyVAoTfpC5h
ueF9AehwLVputx3PZ3u07oOr8e75wpsMUZa0EDHbDGwamByqLa/vgqfu/wOG0B17v+lLCDhV86s6
J+ketr4zhCvSh1xp5dufYTPw7PQxaM/wabazky+eB9vXu4sHi4s3jKQsrhwt5KBcrFHt7owzuwlU
9xnJdOVfpyGB3Y/MCjYxxb3qCxrbN9flW4D+kJVbYwMVuFs73Y5hB6Jy6ndGR9HXhbYT/rehtRXq
1I3mq9iIIh5U77FjAmcQB/N2faXGQ9PG8V/IrNCFuSc3s22ZOdqGWQNg0Xv7iV58sFx3oO5eedMd
SDqejFOl64HsG29MEcIL+p1WgL0NaUayfqPGpk1kr972/5XrRKGfg5Z7RaCBHQhNfhRiU+JMr9T2
4Sc0TNBnNAkq8VoknuMvHDM/VGTzReo1ExfkJzzWIt6PrmTUdYicC1Jo0bzcvsM/TNDrF/uKv7e1
h5akGPLAZv98/gHQGrnqATaS/YGTo+pZD5bkeE6GAtU7Umpq0D/PUEns88tYEawpRyQhP/uYwA8f
HCxEnfhAE9cl697gfESAV/16guXYtr/M1MkMxoTlvyNV7qEWK5YlKkogIyOk4/QYBhMqn9JjK7xJ
WQj1NT4PgESkDp266pVYZ248hPL8YYB1K+BqofxOdntL9vhuMouxi45z0al5rYNFK9knCV2ydOlP
KVOmkB+kHiQJ17HVE+IgN1iKYRTAgRmmfwa7s05icK3/7tu+NY6+XRCJac8Bl5O3wGsGEHbB1F01
T72Jt0k2D5q9OxzrjimbFcQy5+XLFmAB6j4nIXPk8qqzfv00QASwWmQoBnh3Ts77/96lXApWgv8c
mHtFGzKcErYOe81yw3bv1c1cQ58zfeKh5NX++lhQ9mBzrWGjNqEeoR5vhDNSlsCcV68CgQureQKr
s5neblz45YRpLwhFT5BY38hLgbGX08DyZgrrCCVAa6e3LzT5TIz5CRby2++DcsNRqrdOblXLwLBp
15ZQU0q+Mb+cCyZaI9qHLBQdkwTfigkIBXmfyNjwZAZFDNj4C+VPMoZk8clA72X1GODB0y5N5mnQ
5mW9sCxLv0N8y8PubPTgRmmR/vPGivSBmEt4xqJZU0YGH6Spq4f/9r/tSDNuRu22QPCQROdxN0go
HudXgOr9teweX+FmnP8Zxim7uSGb5eTaYOjfpveFJmLY5RHFg4nBpgp2PUpB4yJRkqBk4xyDvpjF
Uzr2m3rJcYfRhLUlOH6S62NgQByM3fd9rtYuT1GuRbS46jeNhpNn40b88fCQmIhE6Cy5Femtoich
1Mg+iXCSjEQix1RS4TURkn4sAHETeMoryPyCMJkMHlVe0JBnn/9028OiN/QDmJ7DjN25xS8PE3RR
3IFLFhuX/YT2gKjkU0oDW6p8/BgYlM4aUmjnu4yaz99wf/8g6WuF4jNw4xDWxdDh7eXO41MsGBBl
1YwLqSPRHU46JWIHvz4Hwwkk2OyIAs7tNNRCfgWN7V6IRWJPpblm95IxgWB3KAVOneXX6znMRFIE
R2D2QzwOmoy4xbAcJAiiOq5cE/KXZmE3oEj0OXe5aF9A1ucclYRPdMuA5ylT09XLRKdMoy5g8o7m
E3kXKRRnWGEOccHOlUzYy4nYydVz4k7ofTyg5qnJsc93o2sJEaPOpx4Dr6+OPlzl5T5XPpBKIWK+
u07yKGxrQ7gEttfZM4vEHHRfq6p/gWr1LpOl/iQZd+AOhO1JeJ9n6wqO5BSPmvaAumtqmmkT3Xgw
GM1YN8TTs/RlrWsuSBnoC3a9LNR3D/3vggbsxyWeE5X2JwVFHMSQyXhIL2figlp6v2ybEXw6VCGi
QeqZHkzyJHFsuXBmPqLucpmYak4kq3nQjmj21wHdH/6WP7c88XkTnQXnyEiv7KPaQv/cS3fKTFE3
1imADYyzevqUIPW+XCh7VMCpd1Syi88Q0TZF5rGEzp1qVJAp2QDOB1EISwgdGrQiPT7yf1SS6ugq
Ly5yajhgYWeBV1Uj/umgbtoDsknf95c35lab7zQl+UlvNqS3IfDpixRotwQMmEaLKTyM0vy+j0lT
H4MsiFAUzfUygjXnNdFS+5A4uQT+ATwXvol9UotgJ4jzfkh9Qaxsr+RoVG2lWEkhJuFSdXKk+Xf8
unPTeDSyUstYBMcoGUBmT+yaBECV2WP8AbX+mfNP0rsAtyV4g7bmwI8wqDlW3w9uU2GMLXuEbL65
p1SqsRNy/URm9o3D37sli4Tx7NEh3WrXzdovEsQ2v6uvPbJ/wji75PvVWv5KhfyKi7+eTSQfFwMz
AYdLyrDY6iMQnhGVN4pL2XgSfwEO7A502ViLmn6j47hOVZPUDhZYgspuK+Cj77kpWS/W2IADRhW8
h8DvctbcFO6Yq8ID0NpCw/w5n+ckXFHAKm+j0urtU/CJQiOQQH7h4myR3Mft0eEnfVlLsXYzlNLb
7UbfvD0x43O9O5fBZ9a1OXUSKPVEJ9qNHiR8EF0sF+uFVXGhW+6Sjwn8UEB90ucOXR4yB6kLykvr
lObxZRkeZBteijoml0XSDOvrhwzzw8UZtg9u/2U0ZtVTjlREvAcRk6qt1/24ZDuVoTs7bl1/I+TN
lkdEzqV9r0nAqlQ0PFNZP8LYNdlhbmfo9ghs5LqaBA3wTWwSiFlZQRrZxXKhrmNP2R3iX2stLYo2
m1M2xKuxK98yKXP6jGdN1n7NIItoU1vYuYg9L8ZW4tUG5PsaN20KhiQYLQ45tJCSpIYvh4suYOXT
YkAnEAS3TpzUiwn7NAvK7h5WbjOpNKBvPqhvDTecJ2rZTE+15sJB5JG8H652OuwSDUvvvU10EX05
PM2T3Exz3VBoHKPoQCYe/inkZIOsBMqwynn9CGV7TLfA+ZrNuoLsxiIA//RXLN0K1kIbRYPrlw/d
YsThV/DRSMVujQmgTrYMj4QVulOwmg6I3kB7r6SUTpJY3W1zsuyD7remRyWZPr2d6LsGaTK1fIkF
sQGIb7d/GAg6VClmNaxJwif0MbM3pKu7b2ZUE5/pZZ97tviNeoOg8CMJN6pBYq8tEGR1eXpxaGYz
4FTDdv4wHmXLuxN7lPlhErlW3yBr2gjOVBhDfdoxa1+sYS0gPJ5aQ8MTgKlkKhc+OGt3nFfZ8pj4
NULRrhG+9JxjTgv49T5XBHCWnsCvgN2CB8qIaouNaA1X/9g6VD8ONFbMqH11QuqPUWfUvsjkWtve
4u4i4G7f42nb/AtOWsQLqo71r+XFRN5AKny4Q3kJaNGXxbwUaXPn6G8deA4uoehU6Jmny4Q46KcT
Ljy3mRIWmj5PqAuVf58z7n/pnl4dUlNzus+84usjOJwnsP0m6TDYDzOTHLvHtKzqCxy78XgZJrZs
2aGjtsOVNGD6hqfBJi+Pq1pLhUdQ83SH87x9GJG4xg975VAcexVe7Buh3LS7ypgqlh5zrICvIJKy
x87bxyGF3usQSIHr8YPmK+x7n92CKF5XyCqLzXlkCl88Isl/TFW1S8vzi2A6buvXKcJHAGDJYYLh
AfK1w0htBkgtKC/YyLh3JdMMhi8TlTtgBkwj5Tq04uhC10Y6CwbdDc7GqZiTNz0lOdShl2KOrZa1
ACWTyPUR+/S1uu0iMUiUWxtzkjXwoofRLmJJpCGVHrs7bFwo/saSOYPTTqzzwsnGHaqwQ1vKGfIg
YiIfsTFs839bwcnO1K1a4rwqSApGsERV2pK06sWkViyU5PibdeNpRsPjYw5s7USljj6DTFpY9S3O
0TpcrZZuOWXYTsuiuLeNYtMRNs2swekxx7RMvfxuAO+OVbLT+H+rPI1Jzxq5X8drTVA41BjXYM9M
QsrCWuvhMkCmhp118RJi4woJdpm4u2wkjKxSvn/s8aOzf3QLMt21/RTKxqOe2Zk09GxO+f3zmPEF
JBTUnjlM6W/zeR7DywiPA0428lcyPAV25mppepjQXjrkZwo7c8B/LDo08bLSU/TkRKk1QcKBZ9iF
w3QFh7ygeidLZeUuvcR4WzbdQfsT410EiAUz5QxdAUuVlkwqEgufZ86VeNIItRC4wtAXNWz8sGUN
IeBNqXCJ4yh4LfbL3k+0AwrZE29Z2GtJnfR1b52ACK49heSKBDlB0lmCYwyh4NCbYndCSxilBwIJ
he9pGlEwDI8BQC7cofB3GcQ1okcfjlfkaScIzjuy/5g2QJWsmgDTybUGoD3sMNtV3Y1dMY+XkLxw
hNc4A1seMiJxYhV44uMYeFyHjqsNNefmMfSPxcDrTr3GOApveAnYTMvTBh1pgqZBRMoi4YimaQpI
KDQi5WisOfsXyIWQEK8GACM9IYo6TR5DIzsIjKa/vxMxr1oqSj4bP0QQ/br6QpgbCEJjP3a7Uf57
5jEGlVTfrqVm28pQWXppKzcF4cj//o8ChWHdUT+6mkQhAoGPH9B5HNopkacH10182Ke3GcmvTm5v
kzDgDfugQs/FAJvLJSMvoKdgfddqLbjxLrGAdQvTFMU5iGGVciIxqLXNHzxoZxLawlPsplx2RV2d
zOldHoIZA2LHFf5TrFHe0Rxgk96lH8HsWS2gQ6kleyOE6oyFpE5AoGdfoNLEWFX/zYjg0uY+Ex5w
HKpJ2zmD6Qzd8V8cZ5PUUj/riRBM1McxHf/sf1cH2y5qandC0j+UwGpQp+EEJVByaT56+BYgGQdX
b+AP9ubog266O5XLDhcZoGWaDUnYo2W0zzMrczxdSYqLGOvv4lVj2PCvo57PLWyKbC/i4QuY8qXp
QVhY1+Cz7wNXiyqZp9FtfYYgKW/qPOd8mjsuT+JDytovD7p0y2Juv9KWCCzbH/YTEhAmaR+1lh0E
4wWIY6gyz4OP3JgT6Zwt+LVKMcjg8BxecH6Unva7rjlOPZSDE50QRNwGJuCicwcfHOiTiFJyF747
txfFvUODYVfCPabwnMrPWr939vu+bQcBKPP1OjKE9cibGgHflNMY3uw+GdfE1n6evC/2GfxyxLBv
6qdeocGrKMBB8SC8DBfsN9FvioS2GRjpip+YbcnCy8+qjL4tODTpEc4VAqG1FY/K2fLBj3FmCpGZ
jE0BEKV3mTUVlYQ0rNuMoG5BlKI55TIT6Pk5RQnXDMPhg7UxeH5hASmEQepI9QKVovIDOouJo4ES
pYX4ul4oHrZpGoKVHq+fweMJrPqiX2IyASBurBS4THYv1YAOE/DGB+yXSrmjR0w6RbwcRjSkazW3
3GQaBeGjudc0Uc2zNmVf6w3MlSVh/ms4y58eN9yWg1Zncu2uq/xNQUsLOybchDUkmlmrn7oPFcEy
ANG0vsTBeIwQGKTklzVLRVmcnSv9BRPwMrLylwznX0VxElszLZ2FcOEcIP5tOi0PY7xonkYYGzpU
6k+O1eGLclebwEJTJhAqGt268hgggWr6u8LVs1ana2i1VKOEc4d+1IoerP6+ygU0d80epCxwobc6
8YXZ82TypvC6xzHcS9pk2rdnGddHHyginlPNu3t3A8L5zsLcdodZbzpx4DJ9nEQjn0gxMmacsw7p
1tlA4rxr1buZzTlu0G7kdNqE8hD//Kto1nQJnraxQ9z88XIEUhGkTZk7pgOU2SIqpWpWI5SA9+EL
HFlC/MCLp3hU0DhZ4dvg9TmP50ImPbuh+A9NaiEYjYthZiveDFoxi9IhogNk2UpF6UUyJcsWc291
GPfRt3wk0hVvE6FUEDt6ecuAUlQBVF0rZ+AyBVlYrgeXfemQUi/NzHIFC9oojDbydQvvQZ3m36aQ
E6odhiFkQEoyDmxKUEWEr7qCnHQ6hVCUOaX4n9VbBTpUoKgfSgBRaSZ2DztYK5uVhfWIYVaRyjg1
05BJHmH8G1yaeQ7Ukzkauw9yqVJjY9OoesmAd9lGYDCdw2f5SeW3mD2Lar7apFJq3GobSx0ZcSxM
YDCTeMswl3xGdXXh2/ZMUdxNxuVWuy1hftzked3z7KU5ni+WzhWaMuMb8bW1BxtVy/HPxkUYa8Wf
lM0iyk3xy+nME0sgqooUmtFCIcOnx/RJCOyjMXFONNBp848iACL2KhPBz0j2UsJxnhBp/v5pVlIo
q93O09jciqxZKYB/5cUIxiFkVQfs8LXQsB2ntSvzS3upwMTFSDr8BtLG1D59FEE/8DV/R7fkprwi
bGEUM/CwOcMOFbuczr5G6tGf9/wsCkuQleePCyqI363PAvxCl2kxtNn4Q2nTcIEgrUJFE+3EWd2b
YK3fWoKpj6/CpIsmpHWCnxCoSaLKsvF3xB8/6UeNruJUdvuZ1Js5QmK2WUC4lkmF0kCQr+jaDAhz
hu1n3Pudy/B82ZT9deidQfw2P+7OBAt1c3XbgbJPpGHT81yF4uY1M6Cg50dSxXgH8g+n4NEZlbib
Shz5mRY8z3KUvQMDoORn2XqalE6CCM9FGIhK0h1uYmf/JAcCcQ+Ejag+RxQm0MO3Ni+aCbbeZPVc
1iHTOiu9WheBUVO+0A8MpqWQGVmdL2oaX1oEn8HvkukR9faDeVwpcOkxGWuXmTxRFvkPBAP10Cf3
bltfF095AQlJNhY+dlPrj7j5zYEJ5Sz1TRbVnuHjxDJ9pv6VlOcGa8DclgoRRGRlm/DwSv4dUMEG
HsGcmJj2wIgRQRjpwoXVvP0IjnAQx3gEFMAFj5IaLze3UKXvETzen/5y6W9U6kVdVZdUAcaMwHSd
jM8r7I/X0JpV6H91DUDCJktyLEFdPQwqJTpDsbrdlDEzKelGqGGl/PY2M6kq9eidIhb9r9OGMIth
fNHMzOpdKgZU/DdpMwu60qnICQWPkCMPGPYlss5YX6+96qnMmbOGxxTE8wvpunlyLdIo9gTl67yN
caXuvQjoJNP/b4ZCUN3bk+KroUNdPjg+dTkDY3nY8hDWL9NgNPgF5PvqHdaelNJUCvaHv3525Hr+
HrBj4B7YecFTXLoUCEKHtK+sjei2huFMo+e9L9RJ2/NhN0erIp0rvNAKV41Cm6BLbkGyQ3kaHIPP
VdNz5ThScShFTM7UXysldlewpqrraO4rvQL+tnoWiSWQ4YG0FC+uPleVwCzWgM0258Pzt0Siynnl
HgCw6peuhjao7u84FgkRYtZMzivw4sr2c2iRd9qPdOz5+Wws/566BEc3XPnyRWv1RJzLBCaIjhJF
lvo01VIGkoI9DHqvKntUVwPhMgxUHx/CHnRLD96OwsVQblaZABy7fjbTiyzJbxfIm5e61DffipJK
6XNf1Hzvpyw2uFQ25xCFVizzkKOQ9TzxKQsMbwJZCfojjjHlwHm0LaYqCh5xNNUebYgwi4OUzT1O
mii2WvezLGqnnCrI1XjH6XhL/khYibrhOffwlBe0XZEt6iV/oISTQxv19rfFBYW0HLl5s/Hjnf/Y
DQ2PCIFkkAFfof59uG1jsH5bVTI1kzlD+LolKdm6FBwykmklF0qXTP+6hn2bao+1lMgsP0XlojyN
Pl/a+nCckEv5HsggXlk68Fx7mbWf9pZ22zrQd3gJnaBBJSrcvpVpAGCbL2Uq5PisGV2hEr6vOleW
9sIOcJixsbvI8aI9Oy2cM0o9cuuPgX1ajeYw9yb+7MRo5hnE38WRZ0pVzpi3vKEqPG+E0NCtZw38
yiTlSikmwX1DgqO7r1CEDJri8qK9eKDqZGBxuKYvhCSLyyUXR3Rq+NMcFSH0cfNBnQMC72EayQBL
v+KFOKtw9wsqpDATDjqeEMRnLFNW5DUUtWD8L6D9GpE5G/hy/FgNPWxZrBZjQ445CowpmCRAnE7A
G3AFeo2Crg4vjnUjbH5oVHxfZfl+i5Gb3hUf/PcHtmRQgO8ExqDp3d7KOH3wiW7xzgRjGQ+/qP/l
8Arb99FwggEF+CxeP+zhZ2hsxP3rph3DdOzbOcLEQg1PGJH3uS61A3CUtf8dmZdfnrsiD+de3K5r
BbzXQGli4zlaqYofulbxv0yFl2TvhHQzMNrhPSqeyytXtnh7+POTUPM6RV+aMJdB5BxB2YVxfFIh
w3oeFYdYV2oEERwcFk038hzyyBzykctSzoRX2W7eZNSewSlP951OsXhCOIENvtOwZcGd3dPp8/tO
H32LwfdfboA6trSLWZgvybtla8nWRnG69Ho4Ds9VB4Nsj5eqUxTQ4Nxja8osEZr29E47ur1pO+sR
NNjCt9QNeyK7+hjgjc+wSUy7Polqey+sckJqhAR64MXAYOWLG4tXY62I56fsFfNEW4FWrWtViz3N
2kfMjqxCVP2Qd2KPQsklBjI82BAS+sopjrj44qnO9epHzbufXqV0n0nlierPMKH5aMcA+jrqL35C
7BhEVFJ+4/mlebjCJdU811cLsmSLA4q1nXu2PW/u+ko1Y9lGSnrqwMlWVSpEFnK6eU+XHkZ1GrtV
J9cCMdmao5DhY0OEEJqTAYUs7jbIdXjz6pTqv+1+ZYgaeNNHnvoraDrtdK2G+XN3Jy+taGN9gvxu
On73enUd4l7caXjgpP9M/WjuUZypZC/n+oPBGRz9/XM0eV2goYpu2CglnOrcQOHvoRLBq+dizHjh
dxZFetuBgpi1ubSz7BW8vxwi4SwZDC+117f9oW56ckA9gRWWXyjxvx+RUIrZwIEOn4mtWFoFitbN
hgJKzpf6Oov/ZQXC3ma1Vqxzde1d17yhuwdEnqAkAAqQetumDkKqboXk8hjVP1DOGzvY+9kN8ek/
qxNjbWyuOPZKSrtv20RloQYyFdiomRoEeCe6ffAgjo3VS2CJipaEpvhQ6mqO1ECtIAybcxqWPDwa
D/RyN1SbJDrh0MgNSe8Ge4KhCjYtNB1zhFtIn/KtNzOGu9peSvnHl1Ap2/QivUBuNFTcAcFGfgNw
23Dbbgs92dFHikJfcJxCZbTfnDx3oiuSsHWKghT5RFXzImxoLyzoLIanYI2Y0JausHRZFE60lEON
rMBaPfSlavc9b5JHhhwMY66kKVo7vPyncmf3mLGoht1xP4bRcdoCUSXgm+5eZqdDDdeDMI1TQJGD
6mp9lnIKODgq7747U7fC53hAlPtILrqcM9CyFvB8ODBFhpMX4H9p4+z7qgSJ2sXCtiNpRKElEp0z
zXDhhlSUkbG+6U/Bk75LVXxzvD3dPIfO3ckA71RCN56KON/+JtBOwFKCpgG41na9aEMDbLKbKDFJ
cvbCAg9Ep8gGXcBblTaqPzqtmjEs1dQaNAnRprhvU6wG3yuLOXx2gLKxUMwQ1FgDGLpsfTKmGfrH
fiIu9AWjcMwPDcZ2foXzIvnvn5pcLw/jrJNCST33Uvjn1R13/b97oT0K+ZNkSIo2faA9Rjh3/PPb
a/a+kLtZ5a4qpLi4SVzh7fDdoO5s5D/5p4trFDJLn4Z9h2MwbjpdRK8noMg+LyJNd6Z6l9+aicnk
c551kmGjsDy6lm7RRXvoNzJKBQ6amVVTu/L1Zxl2xKGcu3BsD5gek7lOKy9AP/mu96RmqLYBEmL8
WOps/rZ6Jt5aBggYRuMW+e4IKXOefg5o6P4DUzCjw3nldYBH2ToOVHr4BvxPkhKzu3SJoX8y38Gp
uA3FYCHnSL+Qu8+wGBCMtl70I32y3zAHZScf1Nk9tSrSO5J3umkiLuJqRwIMvB3+Ux4NeA33LaST
Sex34f5ndHOsCV8LKPW4nbEkz2U04KHVCRR4jaUaB+dWqhmIf2pX+B0TmkoQQtL0GSIjgUcE42mz
rUiSnFORi/yD6wyBM9lejAtwp+eP6gbkG3qP7zzOIWYZYDBJ0pHyAPg5MEjr7pn3R2QQ11FWAZvK
g2xcK3G/qgr8JUSLa4dmz15mC8Yq5wis7ug0lkTBx4PuZYKP6WEH44FJ2Rnl7vsbJvOCBT+Azqsd
28DQft4TN6FkEiPuR0c6uoNDMCAPI8PdvoBMlIXX0nTEC/+EnbwUB0goAC6ihwOrmVd/rT8ihLly
vN8Id4bjfiqtOHis2vBG4zv4soly/dy+ry/Md3apLnglA573D8TXtD0rx2j3ocW/Vwng9UnA0v7v
wwExTMdhccbTFCgghRmz5aqm2Vg2mYX61q2JQOViHHmyZFDteMq0mPfwHkj0h2vyCWDUQLMbMR4W
JN/sMzrBscnZ/yo46BXvHL2tLJD7Vw+nRXUFHp+vlagATSLF/tUwWst4PhIyMpBk0vbZ1XLFGw/6
WXux75zvr7F0uaCRQ3+eD85dr5e9468R19PHYObWTSrQIefWqE2eIgx0u68nXXku3xlBdvww29fA
z6HHYvFqRmpJ3+dj7pJs1Xgr03hgg/xPRjuzE+cgfdMihvYZRB3cS7lGh61PSPkFWBZPtjrQaG+8
V+SQWfmRG4nGeUFCGQ/9vmd4S6c+5Eys6Jb7lgHohlJe8rgfTQnPDBOs8oyD3oyjsZ+HzaEYMyBC
C54JHBKCs6kePKBPtMoxrmH2XlCTZQyR9UBORZRABiKIPxoGigQk1IdSr2pCgf1u3JcVBClgdwzs
r8JblbEUOdSzdIkGyc1Wasfqfg6wB9WZpN4CxFVjIoyfm9fkZwZgt6SOe/NrqTjQ6ESYgXWsrQpH
qyIqMu1lCDzstACSnZVqrMPHRjNd0U9xZUCWFQwzcMT31rLUYCJ9Uqy3dtNzUPg955buM8xOcR9d
12IlegTPpzwrJL5Mbd0NJ8vW/5tmvy69H7CFiv2AyjDrZXPwWDNJicR78ELRpHhc4EYipPu+WHYI
++pphgv9MH6xkM4F9/8tLN98QdrMC41Hw5QvIloYD/J7125p1OKw3umay2Dzwu1+uQEj9c7j8a1j
I10kZbRj3iqqG5oDX1dJdGYj048RYJEdeg6y86+f2FUsoPvc2ONJr88fAs2vO3gaT+38829F1TDM
7296kc2k3Rl3ewxAFu66AIsiOcqmmVkrufX0eP+sHYXEjgxSpt/6oanKJmT4kZV50yJl62rmXfj0
lah3wlDgHrvGsfEyO1GIWFH3N7ozqdmCYGmyKYXhVrCLMsOmlxy+2n039r7OGzj1pGNaAfoovYed
DUSrMPjQD52KkIG2W5k/prAXHo6kJUA9E2VkyHfBbyRiu6u8bvlqy75k3gKMv5JzzsXL2b8SK1iz
BW+J/2J3afTT1sV9LLKbMg+dYRwrcgI7IMFO+SQ7dkcO65Bxh29WtDwGLigICHzvo1FOXnC1buRT
RDBLOhARYiqoeYvf2rWlUD6wYGUlhr+32Vl4GAH3+3K5fsiMAhxPHYlplVY10Nkjr7f3UFfQMfHL
I1jqDkirsTCFfyIzzDArqABiKlp8s21BpxWdjYSxLpH/wG6Mc/1N7ZfuBGtUkWR5tEBVsIp16l1T
w0H6cKhATxGXpzmlqsm63OHdAdZr5Trdzab8ISseOOTBiM27nOPRqrZauJSpifFdvr+OJJTu2Afa
9h6awhZ3U7on8Q4a00V7w+penDkscw6lbWsKy28LW2Ij664L0bqxnZ1euxd+RTupB/aLo2BNnb4Z
j38bg/f4u/akjUhdwmNZPxJAfSbPkatIYKOnwS3qgvVmpwllZRGZtvPWsuuYtsYTMhnOzMkdhdIU
nakr3rAsFt/JcahZ52LWJyQTBpowo3T8BBINzbF+ADW1JKXpRNzeti2eRqLuBoxSqlO+y96juMpW
XFGMLtUsJRh4nuVBZSK6RZvz3VMAlX5ic48H2OGUktR0xVLhsKfMUKJnEnuQ4+n/bF91MNXgh5QG
mw7qX2N4lCbUrXBBq29/uQDqKw2ro/LFW1TSwQnIAP09Ge4QmvM88enGzPhgMHQK9lfwTkedv+DZ
JFWDxqr4NZ5gvQJjgZ12kOZDBYDXbaMwHXz+7uq6dyHEylkHomEZLde5vfV2WoZwYGuuYmAwDLfK
qMi/fQQjblEnp+KTdLNXg0krmtd/ui9PaQXP/dxVwAxlU+9uwdUv70smXOKkBcp/zq3yHPEEzFa7
tQey5ZwnMDi2SQGmN8hU1FhHfMRtdtMN7i7kKhBmRV+19XCdYDNcqgxpGQfexbrrFMB6RhCPsUE2
B7FGVg3bN7dvqykLv+6jDcIAmWqWbCpvMWnbzq1W9kW9T9fAvFk4FSfkGLjC1ISFcRGMUukZZ5Mf
LDaE35yX9fhaV2Sn9t28fTrFTCQqkDnTPgRlU6Q2QNMG8ufFpZZZLVmkTT8qzBW4yDakG872terG
vtkZg/3sYS/r480oEIQFfSwWEsxfZbXFUiAzx1ZgZMeSyYsxDWHvr7JMeuLPZv64a6S1U72B+nKd
2VC5Fv2Wv/slu0IiZMatRjRngmE5w6PQIX0LbKalj2oPkLRrh5ZJeBz0ia648oEscOOjtFSYc4+3
WUqgZOPgUpxzLOdsVMxkJkb8dCeeNbpmBapQx4JAR4DAWy8yX5sd5jahRYTkjLoM+Hr9wC0Oh/Ri
0Uo3s1+DRdgV0Kc+um8hitjhQZdgZBsH2F1oVJcehXOoycX3tg6s3hZsAMEdS0rtuGiiQz/r6iev
0VsLhXmJHQRD6uQqFSkJXK+YpcceUPFJVLubG14IKsU5izjedmxzYPGpVkCZTlcRx4qk0kpBjQ7m
FG1L1DPRcY+H7ALPEHxGzwtQU+SP5Xh3SXu+9qrI6QYbmLhFPz9ahrbDHIbvXb2m3w53HB2uy3KK
qXzz4fZGysp7aT1/Saj4aTyjMolmdR0Dmx8yLvInbMiLvu/jqaHA+TSDPPJPOh5gPq3be/eFpYEg
mAKgwlfhY2/e3hvV+3C3j6kXmY6DkX3W3zU4SmXy1J4Hf71qnKczZ8mtr+YqKyy2IWRDDPro9wTG
/o7m3IAPYQWhfQ/8Ra8orphD9BSz11pNBSsN+YVn6fCypOFUFSN2a1+ui8XWGU1a/OGcZ2SQK6Bx
pIPwg54qjUOlr44xVTuqThBCsK+FJsFa/f/IMnQF23Z8O/KCwEAcnVXQ39kA3RwkJ52iKMZFqzuE
DbvmR5UY4lrT8rETiBT0aZ3ELBnTEMc1kLBhDW7zxX+c+cNGGhX/woUMdhbkJNFksjZAPhVdjbK5
iATYhgnw06vtr4xr1OVqrOa+PryqhwNgEmcV+swHnbSEkn6OYhtJT3j0I/nKsc91EwIKTh186OKo
p1pClMqwVFF/0LUMiPUWHVjx7McxVjzV8JFFX7SYh6NWviaI/LuKwXKUwZI8kiYvS2ofG4WuyTQT
wNQ3sfgqYT5dYvV6U2xglbv66k/lALYeezp+o5MEAGZnYZ7MOhl0xfjBdoq6HNpe6a/wJBtwsxUo
N6Z/GleN6jnsgG9JazPdUoIMz97FKKk6iNhdywI/Mvyb2fnYmR5C1Aou2ga+WY+mp7lhFS5IyqnE
Jg8IxnMC6PS5dJ6XqF7Um2062hxkJcUvwDA8vEqn3FZl0aJx7h1zSBLqwXi64z8CpSa1jKWjNwjF
4dPqDKZXHFrGh5TO1ac6IhocDywWu8ce483ZN9WldfdWXTN9RBrepRZsrntJ68h8jrfID9DD4Iwc
ol6YdHiZ+YFo2OnBud6hpSk2krXpmZQCw5mWXLgQw6OzB5TLXqRmjXPRNtuvaTHUYmFZ6NxpZFVM
igUdydCIHoj2+YNpwBIVnh1UXmm5WI8gYWnaSuxzdFnu9Gobkk03C3+UvRIYFLKbKrZxF249tZYO
0n4VoAbTCA8jMeAaDcIkzBhMNm746FMvmVEb8mF8OTWYhy3odx3t2R/jYrY+oYp7Ed5o6EhXOsx6
J+wzIOINuFzMomDG/4QDkBjf5p752MK9jqCZgMSSrwLN8xNrHEqF9fPLprOCP4Hv6J5P1x93anxc
zrvju1m+7vabACZ8wvAbeNaqq6mGh2JwP3+P44r613c3NRYJbePOB3W7m6s32us/UyWqNFZFNDg9
3NkCzcH9RPpwCn7fxRyPPIHmhNPjAUnn1sSENeMkm464mPQkE4CF7+t4CeCWljrJl+1x189zidk0
HmM3hwXJk/RxacEf9B6xiIzUFFtr2Q02o4K45XKzkUDdXUyNlXYXcbFWx0O6ogd5e+larljKzf5T
IzagN0+xz6Yjecb5E2FaYm7AtfKl185TzcnBx1LWAkdp23RiezS+HsB7LM6UsxNevBgzWi+WqJWt
VYtEZHvNYPUMpiyOXeN9IfXIG1JbZCCbtsW243QwurLXH5bR9KWbM0YPpT9w3W9HbRrsOBWFQIbX
eOFBVzvijAlgLiL3MAOjVAF2M3MkWs+WVRKJ7zptczz2MmW/Y5tQle49rtxNGfZ7qX0/el6oSJJj
AWXM7NZe5HpFa38UfHEJEplyIJT4clUrthGRuqG3J5PY8nYw7lOsD4zwepVdJ1j+rE3uKVy3msEy
sxFeZTBq1sMP415wN1ml9cGzFhA4vcWrgeAsRsJnZ48yUR9fGxptzjaEktJyc/uTED8iAjrOjCA3
EaXq09vM3+ifHTF/vkuYfBRD57iJXTzCvEzkb/3EZsc57BZIL9OK/qQ5dySdxpbr/6dfo3nhKWP3
ImUXhrxDzUQL7AvgS7SRJ9gFHp4huyDJjYLl23hWANlxICjZchcSj/yZ/PmPjNiBaV5GcepcY+/G
aN3yJh8n9sW5hjCrvzJAFCfc2XSn8J/vykzBgBIZvURpjsoGjkIIzxAnxqWzIwz7hebFyv4VPS8i
ogLAJ9yTKzpDxuCDtloLNVgIfAcih8/K6BnsNS/16nv8EDWXZOISEHaPv3HTziy5vCjVrIdAfnzC
6+E2z1CpZE0PHur1lgGEvzgNc+zcfQFAmAHMhlR9QBVic68GlKmNAykaYI871Ta9FMbtcF9M5aJ6
MtH4ZThV9fMnHnGPEUnIfzLDoUa3oLYnK9qj6CtxXAeYUKpxnv4jCkS4b+MCMtB2g3ZG7bsuDl2Q
2z/MFFX5b5fvzAQ09cP1746z79balpeM+puR/xrxGpwem5qJlhpGYdO67xZcX1Yqz0ASYvG8qQ1X
4rLmMIoKRs6W0DvEvbDL5MTOUnvLtTWay558fK2Avq31JaKnP408NCQn5vynfbW4zWw02wmv1J5H
waCTSpHZx8opXbVhWLKwAh9sbZdvXiJMiGnbz4kSkPk1//7YXQN4Mr4HtDGxWqfmScsA/T9em8QP
Xjb8VBSMpYQzRnswsqHoqx08gXkMZSpOJqJaMw5AfE/cdH1KDmWSoA2tIKOK02s+9ic2UAkui3JM
X4Xhv4pkS2PV2JA1tdg3s9L0ElJIo0vu2l4gDV9p/sR4aTmjWcxJwt9N8YXMjXKxXmisewDuXF04
9Yjz0iFYmFv44yYPr1rLaxc/koHaq3wbsRleZwhlFeJ/zNODRFq7nLbjz15p+t7i2qd2/O8vihFd
+v9wF90tLQd3WhUBvZH2OGzbHg+JllufA8lKpoCe1LPNsv3JaLVopjb0YedaCJqHUTTJKfvyUz3p
n8a+1VqUNmARvioT30Gq4djMyzLA388G73xdc9YGAx/1Imv2EYo7rBl6HME7RMglxuRe8yhW3hSi
dZ+78d3625kZE0fTQCMQqivj48kI7KpQ6Eit2+6lZQR5LuuHjIBUmntl7/DCs6iZLGQDyAvO+ZTs
UvykXVdKPk2rr9kFS/9yugCWCBzMfr1+YRO56FU6ko9+DeoySAWf4tvCLDJVM8767/nLlGoxnjfp
tV9Ma9owPbOOkueC19QVo3d6STFNhUq7dKuffwGGhFaHU9PwX4/yqPhncNZOUjN5R+toS1gKg7ux
ntAsTMEijlJi2p2FDkSrsr2b4juDgft1UuJ8dSgxHZ7zLIJJX0/rdKYuZjKR6EzUowwMWzRdJRB+
EmkxsD9mN8YSKWkV1Sf7l0ApsqH6TRalSlr/TbT+cjPGoIco65w5iD1UxGd19euVAcqtuVJZX7Au
l13vl/iPm4ugEA6FxO1jypbVRJNvzUvE3jiCuCAtOe6kffBiQH8rVBGcwDaUWOJ8tdkBDq8djAHr
2D7z1cZ8vh53bnQrvw8RmvmA5aT9gRZh6yyRN3515G+E7gF2/2BMyVhvg/58quTpvyazH/zM6Uhe
r+9tmtDpWHoRQyMSr7OOh5ei0IsHx6YPr79tP78UmwlvDBOBaGHdK8cSqn4CiZOZE16nY3wCL1MC
s7SBGgyIfrIKib2hNt4g4fC64wandVruHkQL0KooUnCcDYJZdRh/zwmLCYdOidZiUhnOA8mqKnBI
12J6Gn3zq16AR4c6BQCaTF/Y+l1b+/UXaoiSkwnW2GDxiWU8Y2fABamQgYpef+FIt+H0irQXZ7//
0liBNwhcFnXbu0VSnjzssrgvL74ez4W2QbuRFKRUvi+iuDW95RWAASBlN7wi/B5S6vLKLDY6zoT8
27E9RZD1KHJc8LLu/bRHtPN1CagqsAUzlswMXmRENCbSFzVHPdGiaBVIXnmoAJAxy5es+7gCv26Y
S1jbHGx4DNsLzrISbAxIqR6BKQq97qFOMD61sJge+qBByqMe7gaUdFGepwSKl7AHZJeOI3xOhGMB
Ms/hp2KDmEhZ3IU84cVoMxt03WsaBnOwino4wgpFpdIny1l2cIPQN3Ug3OjOUAoFXxA5PLaMvuuy
MW/kNYgxxOU1SLrYYDbkMxOvQ8FbYJCcZNd3mAZ+rGM6PEx/S4DvvtiinqXebg4jzhJ5JY5+CRzN
8K2NKGzbz1tUUcMhhMmqt7mSqjv54RlyC5kGgbOOfxuejPpqCgBxVKfPTi7UFHamNzJe0zqReUzc
quuvC7Sw+fB4xci6ELneezlzXuP5MmkCoQ3a6MoihMpVF3LpC3DFy3Df7rTQ3FJecGL550s7R/z4
i0w2Jxu+ulEZYd8u+qL+ryMtSr+AxDppZxyKOpvymeISUA+nqTUy6NJUzn6gSW8p+H/ra0ZZYKNv
9wKMQtBWAzVvlVX+77diXgdax8vexBZsqcXhWPqyq5xKNtqEKXgqT7nLUZ8gBJqLkwiTZcPghqCg
hohL3L3kTkeWOp+Z9A+Q5sG/bFlqfc8S1djydoCa6D0orTqCXl9f3OtL0cKx30egcRjoiU0I3TLE
jQm5tGwVESdbom6X0spEY6TGRIXD7RbnGfB1KyWggXrRSrGuEwPIC/u7kxtHIsUYBgr4TNngG8Si
Zynf98uuvwL9Lg4JQOgPyqhj9LUWHBnXHm619+SJzBo6/lcuptvEOLgJpupG9JBRZ2cnObLbL17G
TM9mHnt8qq9VcRtQ8FudJ57Yl72a6tBv53RPYJYAzkn6Myuz7yveaZSbowd2pGwr8rdqOSGPVbvN
t4GD5bsc6zzPOrM1T3LSx8V7Qz7tit4mAfWlPTGi+08zqGJDhG+Jac+p/IAe5ZuGLNXC055Gs7GS
qFgbRTr0f5VySIJPK7irRhKHsEkDZZwxH5/K0Ri9TYxYRxULKeGxXn8YSgrmkhzSJGdq5w28n5je
qAHpN7MQA2lQg06t7AZGodAr0pAkiOfQos0uInGLlMIJOnfw35sneWdiP5zWygjJDgwWDLXff4NP
2yI9cIZCEFkp9BaEWJq20C0He0mVzFpDO/oDrbZiIP6scNeWiC/tFoD/8ls2WyF6Cd/cFq80r8Lz
BhVJTiPeTYKgO3YSChVq+bO3QLRn+1HQT2M4jKYkK74Z3CpZLd1L2PSRjxxY50Y27oV2XpNhrghJ
FMT2lJvHXDu/Q4PRthR5MQv6vpAKIjlV4Gyvfd8tLzf+HpJ1KmPyDcYciwx2yLod6VTsqSFbV8g5
x2Uhne5ipWhd58hMqpyHW6U/+nNOKL4yg6PoQxAXrSpzvI63QuQpcsabL18bMOIte2BeMxcJQbos
A4gpd+kG7E97fg1eqbB2wxqtEAw62IctkzTdxjI6uXgfmIh5ZTLWfbiG2dnGYj6kKOLB772agHuG
JOooCkrPqRo+jAbIs97cYuX0QpQLPqtsmfkPHO+p7LM74UW4lflMDgVSGhGOeA6UlCZcQNSc16Df
Z4filHN0Elh0FTKy1IZB2PYlU+WJtk0+4Mkj0ZjLMBMutnPcfAaZZk8bCmuZWXQuXfKqzbfKATLW
mb9Y5dwtbVBrHLdeWd6o4rjJVFMiZ7YE1O6FY6AY8wx7ssbp7T9/Rmyt+GZB7DqV82xHY/f61j6t
hHBWdywVzXxGBOW7zJOX4LVC7kyB7dN4fnyp8cKz6nt+DMP87t6OxcEvlvm9jLtyO9Wky+XEWYcs
1HsIRTMo6LSltmlJeZBCv7v6k2Yxhig63E0p1JS6TcA7QGwQnv/xP5OyWcR8c1Tn5t7aCJxjz9jF
6dw0RNFVw7hNxtpjC9FrO7jZ3KQiZy7ZhWrghVhaMnprrr39fk23PI6EkWmdJACaWV4vcVCfseZs
EasjSwShMNBFoKMnGG0Mjg7vZl6K9NxeThm/iDaCeE0LXxeeOpk0JA1h4zNkxqGkqk7oTdL8INf6
MV3hxpaOhzgz09v5keK3qYRLLmBlpE5pzAqu1mVQrXqN+PXFpxPwxIFvJi/S+fivsf8x+Ows92/+
npwE6gTaF654gp5Md9zkTCd/zvK5IcC5nepIuhCPGe9Wua1AXPKh2wkSqQ5pWtMDg5c16s5MGGpV
HphWHJ3D+BH9iCUgbMOq6sinuQMKQiR1y41mUwMz1UMIG30NPk84ibmLuU0UI8p9N/KTMVCQR5VG
B32eRy7j8JVFcPA4YaxTTlX6g9gXRgJXNOMyhzGhFM2Wf+qQB/WNX0ia2JsBJtQbJ6mZVBrwW9/o
cyCdJvxVuhfrEjboobEqp64DFJjRAJ0ExT7Xf8m79vAkz3QW2fU7RlgJf3LkvX8yzh69W1lTUeB7
8liK7sqILCp69G5/OWTX7pcIP/FTC3T4LIErz5HtguSbBww1/ozHvgGKy65sN3jomHHk7hdAZAet
DT+28psA67mXvUt37g3LskbVLJEEyVMNgjDKoUeT7X1fxLNytP2RS4HRtelH5Wv1fFuo6POrr7My
DsLeCXUFAwiMghydqhFEy/DVz2PKmI4dePl8Bi6LAHBULDyvgKFHV5Ym6LFOanm/aJFBjaWD9C+K
JuoeLnKrkPrB7Jl439lxCM66JKua3ENKcuNAueozD5n2mLyOBCOtbg8jIigvJ/QGFb+yxlLLL2Kh
sPMjkhXaweXEI8PiZw8ERs57yjc2OEyrYMtGSAs0Hs/UurPu22vdzqW2Gvxxn5GNkgvRm55cNCzj
insN32+PHdh4g6X+zfGIxOtxPbm/uuR4JNAq3+6Z6loY7qy42VLcRk9yeT7oDOiwWmRkoXqoshNW
EpfFep9hNKuXx1Oe7jg6lnpJm67kVnPZfnC04hrr5qK+jXi/ZyVHx97xb7d3cPnPfLgQNhpN0AmH
DSabMIL+T2nHeIMkoIt+U8pyiujvemJRZC5Tse8eYkpPAaMqu8sepUAaLEY0mQc53bn/qRtLazEs
N7Bso1ao1eGo5RWec4Pe72eLQP4pQEO54ZKZ476Zd9vguNDOtpfCa/s6JcOtCOw8SZWoUup6QtN5
C1a3qeiw0LU0jlYj6TafGOXXqV3zqMl1qBo7XmPapK+15xtljdG1FCdIwa0LZfxhI9vK9ZJZpIGg
81xYpgdzUO0SxPayr3tYcbxJGuabiItEk1VaZ886eH6c3cq6m4GH2pFLumFP0ctysqOsOc8jfzXL
eOZ62AAUvnD9q3AvvWnqj8S/eE2mO+55+DEXlL/yinxj0yBfATN7dP3SVArKP2w7EOaJQAsBmBXe
kbW9RYsJ2iVRg2tqExyq4yZ1kOkntWjLGZudbRarA7JAgei9O+IzNNdiqYUVy74fML6Z7PRFGEKp
UNYQzn1u4KA8i52MTBlAnLOUdUDmpZ6EMkrS6mTBnhVmKlVmtgKAwqNZKRMMtYhiEiJybLpVSMfq
Cmr1VcgFLedVo8ig8w2jfbX/Mr8KKnRf9X2s7oHWthhLXrnmGCbQLGu875THKvEx8azKtCUpaDYz
oLS60G1J/sdx8o4LlFDjJntWogz/49Hd9kuUL57/yke4IdeZDCndtfkKPIINDn86M10kSs/PkwC+
7xSVG8QIHb3MZJJwTjXbsUnTEMLJuwvayS1lojuaO7Lz9y6gmVVvXDF3B9550niLDMYjIYfHOrLl
+JrJpylDF7l5XZKS/xFpCszjTYbUV01V5dnAJEN2RWpea7IJUb3aVcMcfkiheV2thkGGRPOiIFTn
yL3Ls0Adk2h69iNdQFBFYbsth6B0vQY+qao/8ntGesPHqyjmu3szkDnaDwHARvdrrby4hdyxH0/N
PojMaSikUyYgFPueGWb8PBV+07Mv8ofFoh6vxXenoezXndD/ssSH0yYFMp54BqRkT4rZP31wldID
D2voqqv3IFBOyCy4gWTP3qIp0qM+ko7tBDE21ibo70wcg+nQ+SQy4Jg6ti9BFuLVvWUsSoizO6Hu
5H5L6qMoOY4bQY3bgJlMoMOkdRuQcHKtrkf8jD8XGzhgd1MrblvQFWLvpLlhfibecRAC42oFUMzg
BoOhPzO2b8r0DOvQawAZKcycmNG7+u9bhTddwzBV9ItiPVIaOEEtVoM1NQAc5y3OddVsZAHFTIS7
cjSjmnHVaCBO6z0tW170fZzBs49QNjJehMrkIEeEGFKMTCt/urYj+uaw7SuJM1lgsZH4IrueY/DP
9NOWrDW4Fel36JSlbvcMul/tTRZom/O6FbvLbeYWFbuBHmlqZUnsQg23yhp9+Bhtn46bvOFuWlBI
Pbokz/ofx35ImrVSpYlNELu5mQSFS6VoPE8Y6D/Ue6ANal8b2iPPDEGeonEF4AWLmdch4gKMz5jV
awKyT705JPz1tb+2rn5xBzc4mQdeBH+aNPXrYUveoUq4ydQnOZ0MTJPzGtXf1gX6X8l0674+zmR9
klqmqt3FXrfjXMsnEX7m+caZP+DF4NLO6zdYzdcT82YI1izmS6aL7+rlcigaDtWJ1vkcuiQ8hb7G
Rd77JgBeoNgYUeCkx4Z9eOBlAXXfCgCOgn8scP0H7w2IUJsoqo0Wa6F3Fp1c6fo90UJfs5wwpwv9
fOvqO5JWk40TtW33df2fdh1tqrRcXQfwUn6CSsUwMzCqgvBayTXE2eHxaAQq1A8UY3urLSdNvBkM
ef6WDkIuF2uWlO17/XZasUcqJbSEMADf12t/fHT45WwGzTIWXDK+NReQJI5bBBaX5WnxBV68Tfzj
wRx5sS/sQ44AbxvNfWr5LzzHOOkP7Iucl40WUxJtg62UEhRNEC3quUAhSDwP1V9lqHU2omzisTP2
DZIUwUnA/xRaVdX1qlXT2pDvYuNmJybYqJNA68Ind1PkiM2bP8qXASxBqC+J2JyczeCEqKeYR+Yb
nEmG/46bsLUUiMNieugrGLJJzYSDiaewbjFE53AnTDqGYKbTzktcfyLeaS4VcyNelJHOYXYYp1gY
gnQgUv+SNeP9jt9acfnJQ4cnnl08hcKVuen0zddalSaIRDt2lqZZEiVD+WMetDIRsMkn2AWOLFd6
npCDJvdVDVai5FfI/HttdKr8pU2hqM0KUdMkzJQPWr77efRe3si5xwSLDgge2Hn7VwFaygZjBhUn
0SNRcJHLpXsaQp7c3Ii+0FwWNdutQUfjAFjCWm2+afKs+RRi4Dlv1uFgevxpFGFKG7ZWUNcvQh+0
HU8HbSUPpon99XbBVvZ4Sikp4toQSujfPylsvb5V392boGdS6MCa1XQoBxO4O64HGDvccS4nSQWp
1m0QWybZuerDBkq27NyGGIJVznhNdSRRyoUQbVvvjWDerPrxhYgB8sTLTfUa4emZDIPqi4+on6YV
Ikn8VivnxzEqIHjBw/tPnX1oy2f6qTXgvLVcCSTnevpuPDUgstVlaxokvsuiWUk9xe18YY2cb7IW
5yLvKcHfc1EIf8z+nPsx27zkdj1mUoh6DkJ/6kvod3g0zUbzOSLaMP8yuVM7WgrAryJ4E/Yi3W/1
fUumne8Y3PVcqemHmL2+YlW3K7TZBqWhHjqiBQ/eJrfM0a6Il/Y0/SJNhSj6Iwgf2KEUHXt2yF3A
2yVXOwQrPW7o0x1LP64GIrH59ykIm68ioUDqo0KBKmuj/C1lDAId3Zfj6WYJlguu98Ht6xXm1IXK
F/9yeGLrP6vYC3bH2wMHLHPhDcIQptKk1xFtQuIoWM6zk8drGCUpTovQD7FIgH8MzsjHoW0ZhE5B
6gpHlj7IIoCuqt5YMPAnC35QypDxsdWcqt6uosww706+k3SxHVvjR6OHv7usQ+0yXL1+HJVtFTWx
hEGAJTxAkAO1LQnkdklbHCFXeQ0w2TV7dLpNTVJhy7CcflfXH7mXF/RcewRwbFDEf04VoRMWrr5j
uUGoJRAuGTb6RQz4fxZstRo9wZaKx2zLFnq7tyo5NBDsz7Oe6agjbs/pQB6RfQdzL0X8Vx0nLu24
w3YelRIoIjlvSbndv+gy94PhGV8KD6qWXpEIUAzWjQ2KoqNuJ4zye7yJSOiUM1A/pUCwTvgCPzk/
IhCMyG+eu+OxOUbleoxWoh7EOkREav8+bAEn6cBAZVKBqQ137oY2Srwm0KQPIfdvGMM2Qy/Gv8PU
FZgwUPpHSNAU99zn6his/SzjMq8RUdD9JyktsjFwIlx4QltTpiIctHTXrjeWGFi6dNkp+1UH3yRQ
4eXxmy99gdEWMSODdWD4Dj7UxLvSjpeyESg43p5SURbD+gDro0/5UtBlpjtUlczJtTaevO9zUBjs
r8R5hcqpNeIuKuMz9VP+MlvT5evgk+Zpi0/kQlgfgWPIQkzZxNIXLpzfUYEBAbiIRvXNN5lapR9S
YF9KMfcDCEwkf1i5tfzktZx77ojoITZbZ3HKkmNZBTyfHTxVkQYVOHfxTTlUeom/1nbnkpQD2KGp
WhuaF2VLwAyCu71KO8fN4JV8XGSK71aRqOA1IwjeTs/BNH2HQiZ4RvMpGSoRfibXA1okZ20qCULQ
w5vBFrH7sbhwKj6tmV5XF9yZ7wF+v+CbO22gWfNQ4DcUaj6HpcRBd7aJICxR9KCI6VXLUyPm9JoD
9AgLxPboCvQjXMijvm0az3oSkDwfmQePFzbFOW353LItQ57ONlhl9RIzyNk4Q1RVbb4AhEjESD3h
G9k8aZ3kcrXebe/p8dghq/F6TLwsy82n7cPy2osnvc40HqCwvxPW3H8e6bARVBUgCiZQie2jIevD
h89Cn/DDafpdXKmOAROMJx1JToRsLoHxJZXwEwqD47exbkyfO1vPyi8yMcG0ha3yqSA9Mx7RHfP8
NGxnh28XvYwppKDsIkxdrdLwVrs1x7sTKNIt4MwBFvocqRewVU4esXnigS3yTRJsNTjbfKY1wEXB
SvAWleSMON9mt7k3h39iRPR4RqSzYY2MwdF4o45sZANlP2Oj+GUCCTNUqY8ydJ8osLa8ebIag6fy
1BTV0RG00KPR9/CZqTTBCMUgvXvgZyTrhse78pYDVtuhw+cZNCu8ZHeP2zGJSGrq4YEEF3uFVNKO
RTkLtSSCfgF0stf5oSDynIK1HbGFDM51qxpg8rxhq6KaKopHZOY5U9CfeEu5c4hgYjP89jNzQ6oZ
AxFTXXu9s54gPGk/18OpQ8a05thIunL87BDZcJnWunultCHinwYLpLdUEDDYkXdUCag/RqHHD7WF
a5mO5RVGUznLWMmYp9O0q235W/clk+jRoibwZIGV6goj6NTVP7a47JnVGIR9uYwRXRVLUok33ebS
e0iEHwsImPg8iq8oqoFrrQ9+qHEsZ3o9ys0CEopytf55SZCjfsU+K7iCWFdviL3fj+kop884CIBI
HaI2JJUf07ID8kdkFNBTD1gTbpz4eRWh7eXLTpLROpH+2da+jsu5XSev1Aj6hUfwQHhYd9nhpbzS
yLGEjzRaUVfykeFUjdKWOY+j1wi7lZFOpy7c3ICkvIh2H1ufw52eLvdbNSoOhaO43ZWxtk3KCwFh
cbiGYdB8w+d/H3HKuygEiNyAzsDsUe64oNK/6p3TL7hAppofJtFQ5aq+wK4ulW1zSdj8iguatnt+
vTVU07JkfNxb2FMKl1cMgrqBm68Iz8/0LBpQ4UTz+b0kKhIw2XulyTri1OIf/y3FpUnxoECcZrce
iICe76lfaomtXKBrf6eSaTgEqckXb0oy5+SVsW06hbHUx+ApitKWXgMk8B0Kys0eeyJsx+7BjLow
5JeG3FlELIrq5qTPnk02jV7rzVHE6T69Nb5/Ds/Eh9h2E4qZ06wiZvJZV+ACMeHhAC34i2XB8g8q
S2Lx1tX5IMPeVPe8jltyhAqyiQxHQB5sVDIiHUotrETVxJvgoK4IIHgwQF3s9KgJS9honH5vxVnA
V5fWaQf8NP2mCI1TcDhdmDe29PEU4bHggiyf+/Gp/G6t6og1UN3/FETj9FaAZd0Pn0oQsuVQmfc7
qA7mDlgx2a54+5UIbLRUUyqS03YrHe3YtAVjrG2X04jDWvA8WZsoVmEesx73Zyf47KN6V16kyBUO
WwkwYjmb49AcBykzQ1EcEMe/N0/1PDfB1t/9DkQyTT2RmHU3cUFwR4vzW0GHy7cmS+AlMON0F5S1
LtEXsjV9USJ8TS3TtXwLBhtWJ5i31eO5fR6juDgCN7FUDHpS0BBDKLfqNllQwm09XteXyYVpmyV5
SzODIxS33XpiNVhXswEb+egCR2CcYCofjdidLk4RgLfmuZDNrEaf2oMg2yt8DnoSX7yzZlmboZAF
Eyo6BDfXc4x3/oVsDKQ3oN87jB7gABRLe4KUI+fpPMKt4Z1JwaqhG+Kc88v5vSfv9UVlNOzQo826
BRyMxWT65XC1IdeWhO7CFd8RsSgloAH7r6Tij8Eo5WsEAzFkHLLQNGTN4cfjRFEkSM4DUQnGbRu8
lqvo5zQBu7H3wQCgeIcyxZx5CxILtsinV7gsSUDQUkIBtqBz5lZemcs8Fz57+jeKtXsHp1uC5Pws
8xA6f+bkkmlZ7PrmGqdyEret5dPncvpd0p8ZlTR+ohHAUndDIt5aPkCsddqi/JqtLzKxtCyIpNAN
8O0p7zG1DJf3RJU41y0yzNEWjYqy3xdzy4igipO+fcpuCYrSn8qiF9J/0P+UlUE67pdDTUvFCka4
t5NbDXcs+jxpS2udPgI3y1ffN3AovzZnF2v4l9ZcBHyVt/2RbmZfqs3TPbx0W2uNtcGV/GE182d1
keSywmqmKDEdwVFnWooTN5RD5BSZssVM2DI00jsy56Y/BC3m02SOStFMb62Gi70ialCxDncBkROq
CLScAcY88owtPfY/DNSOxkHaq/MRFjU+w44SceJMsmxnG/lyARXbSJ+uOLjTLhKg7wXZ4/nWFKb6
Q3eS31op6u9QyD1GcAIl0p8VGi7ULmh3WF2yFVr4NKgcq5MDWHx1nuRBffzJu384/uTsT7RBYonm
dGPAmsBGF+DkcOXVUTVVQM0lr0UwYrbu9Xjeet2FFa5EPe/jAxZHL+Hn12rgv/PUZoWjMvd8cTnK
X7g1y+YspIzN1TKBJxnUtbaizZe1h+sC0H5456kFwALO6UNvlqXk3NRlcP8puifLB9K+3l0O3Lix
9RhfSYhmc3p8pbE9kLdXXbSW1cDY3r8OxOjLa+wE0pEJwvsz7h0aUBeLdHduhAgoLYmudCjwYWqB
lhnf/xzqk9L0tVwAwXIW9+n2leBG0U9w7Q8Wd+Qgqj0yHl7LUEQ7KJBgEQbYkGvV1Jwg1grYmjnK
ZIP03sxvmXr+Mn5P3oh+lkM7N8dng4456HP+5HVQEtFeqydpRoXIjBcqBoDtzkWTc06xlCKE3oQ6
2KiRqkYJLVJ8/mGKwUe1uBsHH8uiP1U3mqoEIzNtENDozz/Fk2lj7DrDZZEVmepaKMXDGwcobdt+
ep3oN4ogJ7Jhptmt3LvdcrIUxeSySGtVoDUulbah9qhGEfrF8Z4D8eqhYFPZAPHgEWO5GEi0ZkSa
Y14YAS9xjiXSixQSmeX8g1info/Du/nlCh6e7ZUkGbliALJi4aamd15aZfpob+n8vCjh2nhUeOGq
VvXzdOz2r75f8zWNuNDwjaxyLDh48FLnyUVfDzXFgdH2ewjv3/MfNiwYPKACixrM4wKtrUECaF9n
8vvK5hvAZnQjwdfHsjF/FbK5NcP51/A8CGEgn/7TR2RSvtnsXQzq9SZIYi1dUAgHjaHoa1xWrzud
Cb57/ow8OCsqwO6JbjJRoYjwr9T5Df+XHUJ4O/Lg5JFATv/yY/exgMMxRvZl6DRj412htDeLujGo
GdlBfjPwryAgR8viiJkkMnCdthK/D1wzV00rBNANdCVVRhLQ9nYQRmMHh1aqn00jWU2FkpxGsbTA
X+/WrGgSgcKPq6yiue7UxGQjBtPa/27/1CNyfl8LuhDjJQyvjYiHlgY3Zv7cKOXBfExSfqmbekUt
VH6Pf4EAq4bzF00N6jVMfWPpJTGhhHIJC8bwFJ6+ZOOLSCUa5D3Wpc20DZMjp9ZfjdY4rXGVaiXy
Tt7nWeH9a3h5zNb2XOlbZCqCOQbDAsXJ40WP/DBFyQ6Ovv7+l0uw+10NhtpOa7rGbHzE4DRsHlyD
whYV0DbydzEUz7GuajrO/C57FEN8TcNl1K0KEnQRTIbOBT21WQ1nle9VfpCMTYfbffioCgTIKEwE
50gN5JKqBxkg2kpD+m0s9ex2PqOZTjYDxErKU8ZiVTla6s9FofdMYhP7BpUTsQwpmfB33nro3Vwv
u7yw7ZnwlBBVwqRBOeDJPNJxmWBeYez+mryo28Kjw40Sf7XPeT+fbGi9cF1w3ghFkmOmpWytJ0SS
KZx8T4AUXW26q950CPSQjYvpKZKoCym4k5RLJi5F7rZBLHql0gw4a1KaW4qD4lN+bwISV9twYJJY
Onsf+79AYPLFGxb2T0DNHEpUlLFJK/y7KL9DcsyXFmnVF0dPCYF9ryza189/x+e8fJLM6GpaJ1kR
LpsimcoW30yQqS7oHGL5iiRAe0/6lro44ARviHGkEVbd189xOpjDnmRho0gP1/2Ru3YMD69o692I
ST81/zzYxH/0OONbk8CozIyc618T2wIsB1vy8l7T7YZRTwi1yLHYfVNUgwvSEgp94rtjCn5hu1/B
ZMMTe+FA2HW2Xdoj+yNGMdzs8BDjhyZRN7yLydMUTcOsz9j13yIrlNkG13xtoZxrtZu9qHm46fUD
P9CXEzKxFsM44JItKinw+MO+5Z0wdJg5vM9ULN3LxpMmWtA7oRePAFPQCL+4tOhqeH7rw/5OeRVm
26bP2bSN76Xd0Fb/B9aJ/Gl5ed/xl2NNLoGMk46gReY/wiMrn9xCKS04MBcfbX0cXxyLedBPrr4e
OhQCI/sqU5cVSRfC8GYpolvZonxwY4AG37JyBcTFHUNfWcBzDcd2Gm6rtW1zKPfZKOd29QP17/dR
EE6UnezbcTh9GOnD01fzXr/7OhRHxg9X6irMgp0EdbRP/czBmAiljMbRXwi7JmGCvfm7I6ClGIP3
o74FzaShCm6c6iVFw03hc+KUXSxu7HlBP693mue60dZBLHcz6YRn70s5nIdbwYNO9GaI5ujhQU1V
fnfVqfTFFzOpeGEPE9DbS/4fmZOwi3PmILcXs55Ul8Ch9ZijKKXmCAYEPUK7Ryj2oKRc52hTGnX7
QDOHqdLRS6G0K/LUNzx4mDm3gcQrdSy8Hpn2y9+QcCuNccbbMZbtBBHSzhXy/pq6LOoc3RMKHA97
42aF5aREE+lHDWB5+tgoGpzWhLdsvcYDLbtcyY1JjN3xXYnnqCt2X9V2nfxCeP1RmHCLmevRopn3
AtNLWfEGVITK+ji18DygDYH4aoNUAgwB7crKTKkwJDqkrryFtrmD6mCS6aLDYHVUusoLhAqTwSzs
mpe4PMQhoA7UyOfq1cbbimhOcq7KGskWvtqC4GS0A5kEAx8H7WbfoxbXMc89NL98cWv4tz3ZFtgP
gBDm3s02V475zCnbBreCdRpDLwQujGgCFrTV6mSqIyA4m9qZ4lB8QbYrk8c7hjBU6bcnp6LG8lLz
oxzVk4Slqr9tQ/Wv1ievd7bk9q1majF51vg2vCqfxAWF+oWirlgGlwSZX/6rygNIyNLnoNGHa7Hl
MF+w5wVJLRFJ+KzY20RD+ZiLul5rTfgEOyRbxrhbWP/xK8P66J/BfStYuw8nDjbDwLES9tM6YWXy
ikQdZH4fzi7hOgXQCVVWk/1WgmyPYv6EaYkgc5ev0bt6vQxherU/7JENobQRD2mOiND6KAjVqzA8
ky5NM5XNi9Ct5E1hkqFpxRMlJjCBH24LjKAfLXQZi4rucW2Ye7ZqFtNviEsC6dnxiA/rBoOcvMZ9
19doept2hGKc+0Zd4Ulw0OYbAIlYyJNjnj/cnH6Iy8UhjYCDeVEedpGTlXtfOla1EXHmAM16DaMg
ZuUwGxTrvduiRXIS1Qb4NP2mBdVHyyZl8cFoRPEUHGV6Y6Ycl/0J9ppoHM3OAxDdYIfibxdBAtkl
ynB0UkGELPeiBbBBYcKPTHT2lsZx54KajGV4k6GYCTtA04I1VYcK45tww147pjG9mvweVTUEXD5y
b3l+dbWDRaEaY+90b0MLgf8VjSVaojhm5posgSohTo7gxmHxayANtXlIgIt3fDVwczOrwAe6vzS4
pUK/LqFwJjZU5nOVhtFEMluFQL5IqM0eAM8Esn0ju7oCKzFEUH6txasZe5FiaJCpXCkLOQGCWPS3
y2Fj07fjKHad5g0KsiHaSkFPC4UUk1YciCL6bPhESGnJAAO6xhA07aspXlzOHcwdZNPW3j7j6URF
vz36kFhsm8R33ikd0mIaOVdL4yGHIdghsbemXFPh1s7u8dyqCfUUF2wz/Dn2T6ATx276O4KZ141a
pgp9f9FZoDVpMB6jskNYwmB2S7Unit0ltvRDaK2HleehTGlXmVu6XoU8A94TkrNcOG8i5uEWhM37
BHDNHljcmlFeTmPSvKlW80a6T996v7eKNtC3TPWJO18mw6GYD61JdOVT93p+VELaZWBab9HAzYAq
k7fw1EjTnSUCES8qDkLmz/jHejrrmqEF9mwwsnS1HNNiJuEug6ETMUuodYJBb/S7Wl4Nc65uzIZz
/uJOQ9fBzLnbTF/qyjnjmOp8lARzQT+pps+diKIzCXkbIa7RJ64gyXPuLwAQyuMM5TgGQTTrin8P
bbr1OT6C8KKKLaOQWvPqybhmdPleE9NtKLwvEUdFfHBUYz02Xm0VRabIJ7xX6a4ZeeXt4cB9iCPE
EZMHm4HZynuaQYzPs75+7o1c/LuQWmtnZk0+++K8hS/bZPo2HziXTabUhE5ov7FDg9qgJO99g495
qX5ILFc6lekeKbXvXpbLlbNJLbX8T7SGdJl1YY7uZeVAotjSSsp+CuISKnAQcnYBXNlEoOTURiH9
AUmwIlPs/fvCzfET6Wt8P6symuvHyZ5k2UHvmrA9iJ0ty6gr6BL0BQUO8NODtc8cSXUTg2LVvYkl
9scF1cRSCOuVcimEkCC+Rc2WZvo+NOv6iweg7VKCSF5BDPYoMl2NQoJVTlMrFJpBXLP9HWVNQXzE
lWcg3NWhLxy20RbXHWzEulftP1RhHqGrhDjYz126qwAqduI63Jqcj6gX0FaOCfsbQBMDJmCjF6pm
QTrMTROPH+8AE71LgJXA+WaeL+gnOxovlFsqWvpDb5PaRMWsTsFAmWT+ar1l8ivLh4tuSE1KeUbB
Y7+fqjTOTUW/1j3To8BWQYIkX6ohaBO/kywcx80xtbcN1fJhUCGiASUNKm3mx9dCfT7JYa8YPsg3
JdegK9Kz1gDBP8mgZRkxx4vk6AEYd6WWeudpcdfympLoAScCb2gvh1OQ47GWCteqXeJC+VRlI/Ge
xu57U3yddBvGXCyNVyBOZYtI3v7NSEvTfis2Oi4XRiKNYqxKTuAH6hwDeyd9XbqHTPGDKpC0KBB4
cer4+zcEfe83RRYqc3KeG7RxqVPotMcS/aO37m+X1p0PrbBRgz0ecGU9AD6818G5PgaDbKCbSaTA
43DxiMMep98oxi3HGS4dj4pUbpmcZgOX80IOrastc8Sc7QGFH7Bcche0mkVkQmqltZjjMeqXEGnW
8Ftcl97jD57JIzz9j0XR6szfz2bW/e0d6hrCg0z1/qp8GMc9n9OVhaTiZicLdcZvpxSPdzQcbQ10
bBFULPfg6g/gxf6nXU/o52dJ1FI2ytABWClNAnH4SwtQYqniuYgLpnkg9pUKvh0wMbb5W7/pnXWi
j+1+dXRtGNsa5zWV6S1EvVB/CwG/JaJFhXzEK+uZnB5lATv1tPxq4HfSRMn+Zl3tH7PSGsbQ4/GV
SPUocmxOaBnZ9gYsowF2MtwTdcd63PXJncud5Rs/IWVWGSQ1rGV4kNMr0xM+VD1qCbtuxOqNJcS/
DPg9PHvtBgiUk9GPekUhLz+LngWQ3Xb6sS5RrKnPGZvly04dZUda8cpB1eZVgo/WvFJfmIY7Z+xl
7a5XXIXWb4Smd29gPbNTD/C5eLyEjSdyeUHalbP+DTRSfP+N3+lffWRR2VYS6Eij3Jj6IfAhYLyq
LEab0J+brjvX3+3ahYVQkgl/71sCYxec276tA4/Ez/HKGBSSukye14T+URlwFacEuZ8XbqUoO/wt
Czt19B6rELBachVPgSsqKTSFPoJuadqUG6BUE24wc+FyWaLWemO2dtvw7i6gYsMBJu9TtGPVu+2R
OKs12EkRoUm5j5h6zbXzf+m/G43VWBonfUff9A8G6mqKzK+HMk6cB9viUGeiichml9bfJz+AsmD6
Mv/D5g36UJaMEhTmBN5q0yHX2vYdgQ+Qk/ha7DYrhxgZL+4GbAnWA2kQ2hXzEB8RcfMSP/s2pXtH
TMyvnGQKWDuu8legLIlmnFpeHVL+fncw/BBJJGaE2xMXtXyfkB/k9iTQrN91xY6VAfnD8Jll9fF+
+Hc4nEjZMh1UMS566HhKZQR3ivqAYOL1itz/pP9JUyzr9wA4YkWMnuo3fL01hqco1az2KtYGc73v
q+1agOypfLixH2ag0GAtdcFxHf6IrhTfLa0OTmhFw/yCCNc+tWCR6tDWxPGGwPlK7LZaFa7jznUY
Qjf+saLENj3jE4p3BYoxN2+P2Pxfs4bDs+vnWSViqzs0yX3D0tRn5/ydeBBsXlySZy9HL9mwwMXu
xREGVjHZwYkkw8v+EId6JAvMDxApl2XKXKJQJUNjT/fPifM8A5pQnkSBMTsf7cUS3f6wybc+VknN
l0mCk484Xt03IgxjOuf6HHWRt6GWs37AFAzE28I17J29gCCvmaaKKsi/Lh4BBdLtFXnlTfkBdnDl
u/UMOS6wbA3igG+luXOoBaGyymkvWD83I67bI5XhpBHVV0rven/Z0p8P0JqWiTjsrdMh5JdVt5dn
TM8JUEx2hmemM8K7YCfp0q53bhPCiREtvqZC83Vj0C+c57KtEkDSkAjRsm6dJvI0PxpndICRi+jt
0Zjpxj/395fEck8yhwor5Kwis89fXT8vPFWlwgRcFt/vhRxJPWFwixHIuBIMzmuP1fXkZckaTyeF
zbbbJK2au7pGWesx1W3CxLPKOUE5xkv7PRYEdPR+3FY3p0Lof+WXFP/wU9dv3x2m2vuffPzVDsX0
KnoDIw/JRH9C+HEHdktRmlDgdOftTh7+QF+7Cw6kp7aEkr9TyKjWWZr5WM3s09S/P05BxCwiO/0d
VvfNtXOi96/4FJfVK0nB/XsGRLPB6gSLh5XPvKu8TMO91T6cPfuBvW/d4gHQ7FuCXx4oz/xaFUha
75zoodSa1Z/yt7NixT8PwfUszRzOqpX+RU1YSXZYPVarwW29BEApCdme2DFV2BD7CARPUnO22wQo
NOST6Sj5arWy1L/2aEYGyDogHvKFSbPbZjWPBHLBDeUqyVvPuvcywMcyUr/mItZSgHm8H4izEhgo
aHz8Vt7y1WfkVFhz4p8dptbnFS0TgXYDF54yT1iE/zZz7ggtGw5BGvpbIB1J4+GlPPDYFOglcyi4
QMVGpzSFOjxlg+KeaCRvacxM0osa6WQT/0/zlOZp4FliA5MFzWvnZHZJYCET3rCNuB9IXRhpL2fO
z6Ih4DTwbKmMC2CRMqmEoRC4OaITIKPQCS545aYyrJXTiMbi28DapZUpzPDI9g7HzlhVH8UZcqF6
buhnQvddDPX8C3cPNgv34t6zufYyB+Nnf+Q3vXM6tx65xNmbmWi37FEGj5kE8zbI/g7LOxvbfRqG
CyvujCINBeQzMim8dlBy6hr+XEL8CUReI928zP9KBm539IoNDWhi192zxv5CZq4CvLdn/IpkseSP
pDW7gb7f9EjVJa0Ah1bvSmb+alU0On2mNnmqtCzWTvgdewL7iWeqiC+Jo7LQ5Trh7oHFYqtdjLyD
5x1GnNThdXt7IkFE0rFgD1BMoks+n/ZErJohhfmx/laRXiBCXoI6DvpSz5KWcqfpbCxB+mnoEdOp
+AXjjRhyOeynjN0oE6FX36dMZnNNeHFVbnHAvDE4kTLTOmOqgYRDmj3Pb8cRjchyHtWQSxT3nD09
SgHlEroUFy2QNgeFpJkeyzQONFM+OOdWi2VyVHifqpqm4zOz6Q1TPoqYk2rqvCp62RLl38NA+UVv
XHK1Fr/uWCCz3eigVw/h1GsKvzkeEZFunQBZzf0AKG+YvjB6qL5jGB6Bg39T3v86fqpzeJMUnXJ7
MnMQbmUUnTNaDHSFYWxAZT66RBM2XnKrBNTdMLmDp5PbGbLXQR9KNQmHtGbP4SJZfK9knCLthMju
AI7ad6QBSjuihv+yVkE4Z1WmTaDNqMOstmx3mbvbxiLzniY1JVzCkfs6bz8itEVPRbsRvZeYjaSP
OOEG8u8Q3BROvY+xTRwE104fvEOSK7ullL+jQdR24llk9lzKymZqkxbNUQ+r3vc2LNpQ2011PIA1
hRnRqQnDbqCeION50/DHs4DGVMsKHCKEWLn22gcXszQHWwyy/dLIZ8IupuG+dCAwBS2qiFQ1AN6W
UWcxjvZnhnzm+wC6inWPIbaxP1H22mimtzr+5m6u4uM/FSSuEBR/b5pea9vHqgIaYJpGjMdaGj0S
+jgdkRyLkYO2E8XOMVLGar/F4MYZGtqU9YM7HI0chF8hWmFM7kJafMXqjiXb0ELJZQGSh+VhxV/r
Kgq82atZF9SVmlK6DQJFBjTKhmo4q4ha7lxvdFSlk8UceDbJ29cKH9UZgeD55VistfMBn+xnub1d
VQivDygALjoCmrt6AlZNfQnvEoL68B9L5Ehmmdb1fd0jtmQ6+1tui5mwsptU2ZR0MN7MT/KqvsMv
A1CcFmI43M9MSRYRtSPz6oNp+cZhuKLI8qUin3cMgGc9Dl5pTaI1qDH7YVN6kcvX8BUkQ3P2l2Q+
9K6gaWuCwOQgYH4knnxcec0GKV0OLY9Jo4c7DWRl83OfP2Il3U3mvhcyFbaTU7B9FTUZKOhAfrOe
Wj8sdXuptclv5GnDkdQZtiv1oPpK1Zp+UVc3NYZvYn/Yjr7xi0F1yVLbMMRwjQOu7Iq9V8SziwXG
SyDp40cKBgoEoSzjMaE92WbaL0qh80kgzH+SAqB01/hrF7KnMsBRgSxHvdGBVS1MEhhVC0jWMV+s
RGa8HRudOarqyqj3qLMSqiVmGFcNa75Dd4wtuq0xcnMsLFz+yRrGAb8H5IktOIUdTIhIATe5i17h
1eL+NdjWIBA4u53cSpf/0I0YW8X0uJcRHPnoNauPZm6ArGuM4l3shSyr9k8P3pKdHCRcqBJt0M6i
tTAZWnPKckw8fchiVeQsPSaKEpuu+ZUx0iVnUqhNFTQDGHkFtPtU2TtNNF5bBYUMa9PL9yRr7L4c
vZeOPoDa5OeO2VZQohn4xn+IS7f6X9D5ccVYg+iOzWbcT/T6rGCGYLUZW4Yydw0cE6Er9fK5bwOP
c6TZ+dPJWsjq3mDDJw+DxCkOtglVfT6mpdEsYeUfDfc4pDz8ADqaK7yw6hGk7bgCNfKOPdkDbkUI
z82oHtoqBjsKzATt8ctRdtqFonTob/kQlxLeXZ3d/ybpASQetgf6ksgJmeYPDZ2VWvM8yrvCcKyX
7ONK7bTP1H+Q7IzFpzJbxOGs23FtuaOr4xSAANrIZ4tDPo3CUBx/SR4Lv7qyVS0pAEBia9cNbE4O
Ow6TJ29EJm4PIDl227r9uVZpXqMWDrEtpHOY6CAS08YGbD7T0uOFRRxN3e+pRSMbXY/fKGizz0JW
tqHSZcR7y4y7zicFmdDCXctDjkTTs/mZ12OG1exK92mgELTrFfYbIiTvOnF6iEtdT5FG6ybfc8yq
CwZ2jPU/qET701N0YqIIIm8NgibKWzHf65KCKXQWYwF7ddU+QzZg5JNcbh0Q1haLdYrgu3hJ6cgZ
WZzpuOy5R3iHgJqLgI1FwY3gCH8M639cZhJ+0os1EhSn26xUjYnp6GHZ3oLmxp/aWY3WFsH48yuE
mFFyHBICIyEc+5riNArCcq7jy4FETTLWmapE5PolgtuYc01ag4hZ8tBqduj2bjWm6mthx3CqFoP5
JxmaH8u6bkeyuSJNcVDKvjmSs0PSN8FYhGYKqhIXy6QRXQWBX5pfF6BCg6mxWd0GtdHg8+xlyFkN
fr7lOAXdYg8WhGpS38z0ddIqLawt7mHYmUmtnfIYf1zHj27ClccojH1seGGZywsyQ50xRTC3Z7lO
SfBSmszJh/Q3xTUDkRNXsaKdUgmb1SMEuHy3Kj36C4ZKuDQczgZ6Efzd8mh529xCzvMw94FV+1cv
2zGBwdayD4FvvwXssBxljz6tUvbKw5f+GJjk+cJEj2EdiAbwgx0MgQ3TMDDwUv1qnlRT4uHb/m/G
4HuYi4ZpHQGilzteMQ4wmzfTFMFJ8YXDcbGLBBJ+RxJLThlcPnF1U7X7jxm/ea4ADvUdh7EDRK1N
fJ9snaxZTVhgc/y19N5Hbk2pv6TTYgXqhHLKYs6SXU07qH/ey50Q+Vy57QOMfDwomFoELIJLU8uV
Fo980UDcpJL9AAP0f+zrzwBlIbIIqRrNwxA5nddqJk/IyiA4LyvSsT7NBQSigXHW+vbhwB0pwTP0
UVMwyuTG7iworu+WShoX1IFeitnK0CLIaZqG0120YboSYxA2f0PNrfnr7BiKA3LO5butChLuESfK
YYPA9clzoej1bn/RUNOKoHw9g6EHZbTErKXXLIjKf9wZwU1zZm3qaqX3Wm1Tk34GZRfmgcrF3/5m
Z+2jhipb3m+43xU41b4J21ccbq9Rhzy81jceRkw7ARAMSh56QgceDMMhX1ag5kivv9uGedDMMGv4
+yhY4ORiGqYZ0nAEsiF8koBodjqtifmBdBx7E1kRSMz83sw4ndiJFEmvGSqGJ5ttFlx9wAYZ3Sgs
KxPkaA2ZsoJiaskVec/skwW1Lzb0sAYb+PLNPr9lNsbQ42Nz17cXwIj3RINd41Ahdc+YWl/AjiJR
e6BGwcrpE66cREFHON/6c+vj8jkdezLXsv3+b3IfNGxV3pysACXv89EucD5yPG3+fmo9jPLfn6Sf
fz2LQEujkSsjadKWhDyEbIHQmHb2ma+d0VETXWVUtOjI7ICwiCg/MWCW9Yk4C6nCoCxlOXu/LCZg
CFTXpds7jg+gpNLiorD/o+tgLd/TdZy4oHy8W6JGjsdHE1algWlMXtXjChZ6v680TI8qjV6XX230
ysk68mk+yituPeKJUtkphxbprhFVFq97LbSUcJu96syVphHNMrr3QbQnKnOFt/zPCsaAWFa2ffXK
9GNfIu3bOCW+2Q0+c0R4TiUvNX/3s8fKmlirLtBBXvdWicQXs2LqIDWWMBtcGyWKE01g+B4QAdZz
pkJjYeQBB5r9PKk4Gi+32zhE+LcYV7zjy1s1AYNSKYIg4v3xcYcoC3CFgSYP8e3TeUZaXo6NZC/z
hMrR5Alb9unTM/6m+9L3mH5IeOFXS1zwtwSUSmm05Wqi3wtx77CEhBGOQCu0EPtLx3r1ykTx15yA
2SiVJaO4H9qqsBe3ub3dsjOkiD6wgssAu8hLz3LUx8a9LxCcBS6XDbvR/MqBfos5LdE1XSaboMNA
UDy4Pu+9z/8MYuXqEJ/Lt6eP6vu6230wtwJ2QoWHssKk8Uew4wr3g9SGxnUrFrKZAwYZ0ekzXMFs
ATn1KNbX2tnhY2l2g8b31m+f8H1KGtJ2XMPKIhwQz0nCd788dvb4OFIDAuYmL9iI70P5n8AQW+zh
xhQxFB4sly/KqYd85h+lgdQZjFck4252WwVR28Bx6SRXvky2lEiXEcZtPJlmoR5hKntqP1pbbZYf
bVH34Ccz7v8JMb88CxSAf3bPHsaPBxAoFrYIPPIgibr18UGbpdVECKeQBIXa+ydz1Q/btCIPFX+X
kvyyLWW6pPy0zCfc5FWcmHcFdc3csRTJeMGx14RoYoUELOtOHCMXYEDv2H+haT9gKmyec+0cYgmq
sKzIauhly2rwLJlmNI/LrGhQz8eu0jSI2ONH2MIonAA0K+sxmdl8YUaNMOpLHPBhvW1Rm+0lnObE
v30CVaBd1+rFmYt4hRovby1XrUT3B+dZEREx9HqSL1p1di02XGN5HZRl/tBP2xG0pYz58cfnlnbB
VIThoCCpFh1oLS4NWMu5xNbK94VqG6pEpGhQuRXem55yjhZCxk30udFo23ovSS5gBDt8SrI7VMVb
v8e3c4TXOGQvUhnKzLagweTy6RJ6MjEzCJm0GwF0HIIRdACoKlCP5hnMO3QUBiEpc7Tqlvr3g5zL
Jz4kFooHp3UiFHDyj8tmj24/DtYfskmm/VdjCRVxZhjRZR9tb2LbMR0ho0CyGaQBPrJ17P8ZQdQy
GUWqdcrtlRrWcEyVRm3ytoLsUiLHkEwqgzlDsst7ehixMr0GIXwG5yKjYgQWC7NiKOQWr19f0Fja
3FFuwlDPHhxyj7cd6fmdzmopI90YsVlpwOdoN2GcQbccl4NSefRkNBTtQ1ZRh0s3vmIK/sV6tjjB
gk56mKrrbcuIKseXmAvTBwmsahG3hRDCHUdur5T5EBcXG4ZSvztkJ5bwaTHkVm80vnzmflpd32w9
0q92QLevqEsh2oIUM60rfP8NOeh5V/xh796HCSS/7OvlmCyVPTQQYStPIrh0Au74r4c7Sy877y2+
tD4kaPLD+WOF2T/e+Mum2ILuXlCYMB67pVyNwsxFhiQcF3BnmQrizVBbHqaxhvp6M5uU4QddAqGM
JUH3uJXF4gPmRZixMorQ9EssRLaJFg4CYn37d1rTXE29DBSCXn5Yf+joCv+634OmOMZa58AIjPh9
fs4Q9Jk5kuQJVsECrtGL+p5Blz6vayyZDuuULNdRXHWnsDygKkDqXfFQaiAaxqEUkA9VwjH2PpIy
KlV3lTHBOf3y5lQufQZQRsxLvVpLe3IZQcZfJ0Rtc3IrPkdxBwhZENi+IEZbreBv3dpesVukV/se
mVvw5bT4L0gn68DbK8VrmShYyOAjx8Nh6zNg2NONctsfnyyXNRTgploLYI1Gtg0fltrYhs2LYynB
s4nnCru4kZ5TPjTGx7vKXuQlZB9KOhBCZaPrvWeLYaJpSE4NRhM7Y9ZBWJeGCw3K4BEiXLrIh8zG
4Uck959JJ5a6dNjxldsQ8CuN6L63SR4EvyUyTJ9K/+xntMjqrnxEOck/5oxeiNZKOWrGfYflJ46x
O2eQCPo/tQnTColB51fZB4vH3BYzt8LWxx/SE1J0sZdbPottMMTqQqA6DbxBNRGfDsAnWLh+Qieg
6dNlcVT/i8rFhaA40yf/SDkvu9NYzgZ3vpTy9QWOA1/OMFkInPQzFMK4wyDQa4/wV2Gt0rUo7CUX
qQSBBjhzz/DfUyJWGdXqvnC+WEyJ57nyxsyRBCGuFm9pM9eZjkzOZDklt62VSDyXtcmD0JhkNYPb
QATKJ0kv7be8eZ1BkHcEWS61By9enqiiUBgBKkILDe/jmjI1r6OuvvedbAPI0javdOV2dxr85rnG
zSzmenDwCyh8Y3Qmm0ZW6Aln21IVeMBqsrCQNAbDmoGfJBnxddaItUH3uWI4HQEJ70pttgxDxYPH
cM3PIPsiwrbIcnh08FHAIox67133P9V7YURCf7GK20wXiOmQwgGGDkVa6AYYf8M4r7GnNgihkX9f
vJmkG8NFeniIbaFjEM9AnhbTXcoTmHUw4cxlXAkEjI82u2O57dvIEj89jt9L5SQNqbeMHi05WsxP
ogCoSt48sEGnurLiJReUHKfbfNB7+14Wh7unnx2y+X2WUt+1HvOoUVI1csweH9B8hoNPVicIlCSJ
N928zsAQVGJLOcyNpeJbXeg78N+7DOgCkrpT12iCzgGtTzwD4gyewNt5Coy0ZNEBZ3vyTT96cSom
2MmOBfRoDvETBQMF0b0+vn5h39ByEeutVW94ENZYrPqr7/WR1eklK7oY8jQk3D7j26Z9YIWCKTJE
b0Nr7AW4omm12ond4PwWN6DkhuktDRDoyEIlaRYMF7ZkZsrWOqd/SBS3hGY8qqFEzNr1qvRP7Rhf
G5DafEVsStpnmCnqjuJ6Mh07tCl+M4FwNC2ZjBOq9YfP2GdjpnSq2JHBqQrhXWDEgIl3DFs+hcH5
qPMCY6DUfGPjNEd10y5sormKLAaP+1jfztE81PqIXwmfl6De7R0iijc8Gb6QFb/YIoqw348smwC9
d3JEgK9Xmx6uzXUuXhptDfN8wXM+amvzWuZdQfwfrqMKbpkFwfPx5329p5+2LcglU2eOhsoTdjE+
iVmRv9NFJ2ErUTbZ5jqAvGgSQ3B9H4QGUP31ajdA0+EEFQd/asNeUjqX+1+x48j/hRcl8RmGRA6W
04oPDikfl0NYJ9zKxOGmtvLK3xsAtv5qhpHnDaaKD16Aq2jA4uZEvlPOQDbc7cAmy9UWAEH9ARwz
NTT49KEDUVeE4yx2l/KuiXSN6r+nWDrGDQZOp7Veq0wNWiIQkA88aYOMS9rvcWyTVYeFaj9ecd/o
Wi1pIFKjx1KtEuduqMDJc7HnG4Sqcud0jktf5UzwbLVKI5C14+3Axm54Wd7JFj9vsWCkfargnWUI
ACyreL5TGseKsenZwBbDpLHYLcUf9ZnkMiL/gIZaOy40tN1YBOz2HyKQj+T45KctJzKsbjcypF8o
SC9N7BEvNQUMhxMnUnU4AH/VhojpCBRr0a4IZ1+yES7RM9cb7CBZAOIYK7jPq1gzZYSHOcAn/ZgG
ZycmzWQ9g0ylHyIkwGDCXRkODOk+semq/E0LPKRk429lbHUQlywHM88aoeXPiKRp3WswJ1kc2rEm
c5g/ccTU8DcVsFG2f2bZwh6ZgZnOqDjw+pjQ38DSKsxSSs+4W62LPFNrItkzryFh0eO55ghmlcP5
EhXEXtWQjLZldy8EFckOogSsSfnaZ8cE3XZBXyk979smEteJiUeI+4Uz2/IjsXh27OHMqeAQ8WiR
LgyUxQ14/ckZ/+b+vEnh2YekKurfXYLqsl6gwQj7tYHlGzo0oLSR9DDUCSeqMBNKiGDeiJ8OpmA9
0FIApJQDH2A+52KyOVoaDALTgDueGUoNu5HTq0zQuZcTJM/EDfZalZNQWtzpObmPRDtMc53GZ4oP
1WZO9S3+ZiO8S0q5omT/GDTae6kwll9HZcQpuPf1udBcv8+KPpin9+Uo77mmzt88XeiW4oAVGUY/
zT9eCSGlZfEe3WTgplCCJvTCyjA7R2dcbytB+7yiQyo5g7/mE9aKc+0OOx0rOlxe50bETld/D/yq
D7wL+uuLOrvzyXMei6eOHqLLR2EbIbjS+Y/KokFE+/DjkRQSj6eKInQS9W2xgphnV6GAh+HtuPAM
J8AIPx5BF1AM+nJjkNwDyKnZcdiMuNgm5Yf+J4YZxdZ2IkatznqEn5x+MiFCYXPPZa8QapABXuEX
dxWgbwifHlJ0I2sh51xJ/bJXSdzMry0lHKQQGC+8uEgjb1LtLC9H15TZCgjOLGj7Qti9Q8dsi7S1
TZzYTqfDiHWvG2ue6sy2yjS0qbjeLbS7w4LeZCHgM4u/bLghy5LFDAqIaK/aFCCpad1iEq+2JGKu
AniLaYJJIcRfE3gebmIX9w8jhj3JoOAJ2P1ofb+VRwAEGiQD0NhoWbWgeyCmG3Mu0MB8TDt/gWSY
8iYGvesgcJwS3BWZTzhK3fCFfkQno0Ebx5MQqS6NsNMLZGEC6Rt8Vpxm3ta99HWIB2JngPWFxxyn
axEUQz6u+FgQs4V3Zl8PrLeEmsXdEJFTrZ8YYYDOKphRt1R+ZOa4DaxeYvSYf8RgpA/bWeIptDhn
JtS8ctngoQ7ycmUWn90aQobRkCSAqW3q8BaZ8ngrMH+wSom730IJB+AcmWZZG+maO/2JH/hPB/R/
sWI+mjdFXIhTeaE05lZut0ErLptBYOx0His/yNyCamZBHRpjuaYkFg9ctTfCwPDR4qEEmhgw9qjG
zFQtCl+Q6ip8sA5o74Zi7LJA+Emif0YIv1rkzsZRCUoy+j/b0Z3GdRbS1mOKhA3kxKjHndiDnpjN
zqeTL17dWwt8+u8TDDNbeLqLRwmhtLKTnnTbIUaC8COTwD1DOMYU6tOzlaL2tFcz8w6ReSQtnNn7
AwQPO+2QhjEEtXHlgBhNX0exy7P31gr4qYlgv/ulTIWtLvYm2MHt2/qXlTRBWsybD6bKCWWTWKzA
Ig5eO/3tCBc1vkI7IvSTJ5KxrsD40I4zAEZGgw3DENcfCyUeE0TV2TN9uEQ1DlgsGXpBOMmPZzg9
DDfS2DxCZjsx4tQe8KuklEDoax6vJzOSLcZo91niCRGVrV9FoP5zXhcs1yKYrC50LAeTjDtuOXuR
xCUCbleWF6wBvnpklF0b99AH8H9hZp7ZKJTHsBq9Kzn5XboC2J4xc4UkwNw0x82kdLeG0tt+BgaA
y+u/y+3GkyGUGYGh+RokxKUtKaVrgS1KYtoPIWw0sUx5qXRsjKkqwXrzccDlJuTZG9B2Unp5Sq6t
a6pZTezEmyEfoeH6zyXcuCgeut7np1z/gnVRKUidT5LxjfLsmY5XwRTwfy2deU5mIMV0mlGmCa5p
tCLfc9sKydu5XggADoxuK+ca9cJeHTOYIfbXOsQkKy8JY+5r+f+yKjM8B2JPwQdJoBoI2cPcnICf
fKEIYBx8AuMicK5aIP9Yp8JkldvlADWJx516k9+yvMhKROcocq1IvmxGbdo9CaFf5dND1/9yqLNv
UWF+NRElGx7hMeDJeAh1qfIIT2jeI2uOtRSBDJpbZT8gP5pdmvbRdzanRMGHOkj52lJZuJBYLhMA
tslHljfxR+RafrJiVAfPZ2baR39x7XQOwmQfmPo55XnwJmdTuZR6k2fd8r8GnEKG4DPrlqNDHb7+
yPTb6tPDqL0xQwhB5wIdBH6CisBC1x0XOOdkxYtAQ6F/ZUFY6FdiEJ4zvFcW8P+UyDh6WRb0Ir8R
405YtO0ppGYbTnBiBZrL1PU/m6l+64lNzSFvUHH6zgJT+f11pAdO7PDdfpUKnHWB0e0ql3uMWLoZ
KAMXooBYJib/dXdaezk+t0Js4nGwkorLJn5lqkLMHuMDkJ5Rht/Kkwnj6uWrb7mJwZ2v6Eai1h57
YH4hSDIIT87E7qtq2nMAXI8uN6+gKZsceC2Fk7aQ22+tR/IL7AZaKhXozoE+1ANGGiDYLYyamgsd
cqI54KclEggPPk4SFWwdds8hj5TWufWS+BI4/WsoCgsOjeDeF5xFip/YmdThSOD6CB+r4Y1kiXiN
NYiugdSQdvTuob8AHNJaiMyTQ4ghXMz/CkvsbKAqNLjv60wqAQDgC3GnKRLUamoq1omZG58V/l9y
KLtAmVqcy4oQwWpfaZnBSeCjJvwy8r2yGwRZ/oy1VQhumQQz1IlOcXzCAbbjXuDnAESWnWZrAbA1
lsmY2yL+fk0sNns3a72OACEXI9dbbNvT5f/8VB7jndfE6hEx+BeTmA49mWVEcu426ej4nVafocvO
FA4vqo67Z2voMzaZa6siCfsKb8E6Yx9vHAE6wYt+HGeXsiYxwNsg7hOZ+J9RwELx98Ke1EO+YssK
gbVuc0twgr3G5+o9hGLPDY8pZWtW6G8sun430JMNNLp5pVwl67+wVdZIx9JnjCs0yFwA48Ocbl+N
enfLi3HujP6QSZPkaCpyo/G7scTTb3c5gDRV3XWOtzW8sM9feEj7KqaBP/IzON9iLNezOegh43bm
A9frMqFUDNx+LoYKlCAqGWgxJABUsL45Ms3+8eulPuhbXoMJOzvLGvwFDQ1MYrHh5gDONOhAvJRA
At7Wspeo45U8SY2+j137Ysk3k8AVtaSuU+DY9/yEfR7xo6tg/NQ2EAKiIKvrCHtSEYG6Gp1M/kWY
KGpO96ZfAM0sUqKsrQphenkZCZSgALb5ZKyDSiCthSf1RcEsZQLPkKBmA5MGG8IHW5ySjSuFId+R
ZGkgV2Lm6OKxIX+SNEg9JgRVLVp2oqsa9xQqlNGAww/j+hx/hjkwqBJQAvr2F/DipD/nVDmuIUxa
95c+HIZaswpy6/BXeLD64ROQbwDmEd2oPKNONldQ0fNbPp0UMpp612X80NNepps3/V3C1GoX87c1
SLcEjn8cOf29ozeA2TnqmNux6RzHh/HQc+smpXb3NdRmk6gD2JKa4U3l35zsI5zJDERCYuU8WIOJ
TFsMScrn+GGbls3i0b68hrTlMANnMoUD/a1yF2JuDvnEPUpoQ2eRbeFBAxZDK8GTOQsE20LhuuJH
jUcPwNykSLC6kvU6FEE8Cdote8xIaCYj73XkuojiBsbwzLp0e0nlxk0LjzJcuZKD4SbQQlusVaTK
B0BRLxWRBHS7rpEM/xe7dzZxvOpypmLh9JmuBbEBrHSlVqFfFqyprMeCKj1csU734iWhfZYnhZ4t
+r575PUGcpLM6hSRyZl9PrHt2ezFWtkfVW7bRfTgF/nBFxNyL94YjtAWspYc1lLoly/L8coQlV/4
03HGg318DDhs6qy4cLD0pUU84bhAaUeNrmwrVAkYuliX9SIkXjhte/qfuyhrjPevbYc3+pCW2X0J
e+XwV7+mJx6H95rc1yVjociwSfgVi5l/9gTPaEoDXBEqCb6MIEQMYwilZ6WIyhdDqgZu93g7tJO3
CmPSfU/HBrZOxq0HGeF1eVzqUaDvciZ+tHeD9lyc/J5xMjxTB70BAnIj+Yl3XpBDJMcSSWGEo15E
YT/j2DIyc3iIfkEqiUQUBpMGdliXbmIRWTdaIAG/QWvF6eSLfFvRZPZvRuYyYwnICRf6Dn8Tzla0
swMtQsWpm5OsdbJixvySVjmAmm4sQoOldH3CwhL1LdW9LZoT4s6C/L8MMGZASl4sNsRKOzpzKVrD
DwHxHeWoORiW8ZOl7VlXKMqZLuk9N0nGCm6OTMVrF4PSf+Jgwh+uy+sqXh660m+8WCmjAk6KbIiQ
+T0b3xMlURDFKgojJemzSZNqMiy2Yc2eTWxvUA1Fd8YrVSw3P0uazKaLMN+yCv6kg7zTH0nZWGmu
RtdtEaoDWbCiopg7HqeV98KvffHiUBDamX1woReMK41K2KdILvJK81LAbSEthAjV9Rd35/m9cGe8
6DEtNAcV3x35xOuw04MDTIz3BasHGUOIrljB3N10RBOxrOGtQ+N0APzpv89aZ4U/GQ/3UQZtSHB5
Bfb6nmAq6WFwthRD4Hznyt5JgoPLEUrna9ZqHqwEJefEY5PjdrGmLo2CvKSYUa0NGGDRFjbe79xc
ppzbCYSSeH+hckI6Gm2fRO6KPtnyFMca1U+DkiBcju2lHtVFpwWV7Y+JnbnjV9KjhrcHKs3U5Wju
Xm1+EPMWvSfcmdmJDk6Q7Hx24PyHWW07uHslsvhVlIu2o3NvUO+njQW/NMSBnDlzuYhdFRbnVS4U
DdIzw9ZpYq7/Js47C6xbJxEyV3W/KH/McGMG5oh1ReBzdXh+f39AuR5BgIOH2iIklWM9+mzJYeGR
pK4ZVksFJ77FTfa7KbkIVmx9ELNGUeH2W3QqCGgsxNbvo/8nRBWv9VcCQvn4n0zLzB33qRqjPRGV
sECinzO3lfBxLbD4H8B7JMSJkjled2OoomBmevDwcEqW/TUbQOiVPULF3w+cMG30EkkMQofyiFHJ
NHl8e9UPmqz1I9RbSf+R40z4t3K7O4Gr11VR01MuRnUOBqTONkEc1f99f2AKzAVElUTXDdCYP6/3
3TFZJywP/GXkwq+xKCi7MTwo5gA0zadaIAG4gn7j7gK6Ayg5Tj5s4WtQN0/wUrdBPLZIxoL9V0xW
MokPGLNhbL/xH+fS7dAuK38wrIe7wbLd71QYly+F/iSiZWfutC7HBEj4EJnEUCvngr5mlzYK9/Jj
shCpp90hzh8eSgBzPXUQy2CLIRf/vHr+VbbVefucRrN24Fe4dEH/SgXzoqgbcfLV7p6v9380wpFq
Mv0eCVaSjw3JectJC4RK8pfiEiHdxoYtHdIhxW5GByMt4x2A6Xfxh7eJxDECaIPFyGusbYw3FuDZ
DYUDbxPIvuCoFdmcwUaVF6wYEGRyB1IqUz4R44Fclyd4mLI9eTZTeTuNS7H45tXCMdL0/3ipoh3k
gxrQ5pdNAElSKrqwpzRTgOPY2OpqhLn+SENsdadeRblbBVdAa0edzCy/nXVwjtGfhjxoAOFnNT15
O1QB59S/WTMXjbe/Mb+gK/9Laq2pCHXwzPqc4wu3+xNL52xurajSYqE5I9lLU0un55JnRP7wXD04
wk2K+lXYtf5HWz291tKykb5P7uL6SN48pMnCY5Zoya+9Cbejxpp528id1aqaJg1DPuSc1Xp5Uafp
ZdE2NuvYrdikUE9h5G18HM0XY8p2YxknuunaEwjFEsTArqhx5Wstt26vSB3y0TyDYT+cKa6Q82XR
fvlWoKoH76bd/P4IlG1GpIlh4D6Ce/mql+24LNYtvzCfCz+0YLzqoKhrUbEdjWWDtnUaelQGxy1p
wUj9QKkM0UldHYRzZb6vrcwVCtizEb89uQiJ+jKdMznmS3gtVAbkgiXxriXL3A+gN02myCRgXVS1
HPt2zEvw7vzLo5rJKfBgpZG2PRA4rrCNXefq/Jw3X7hXvvlVajBa7UeAUJ+hhAMmOl60AS+nAZXx
k9rSDr/p6c4+JxM98I+JqZXj4oNrpGh9040QWJuNU1i9UeCqI/3z4ixLsHjCFfFrmqQFtGciuX+a
TKyQUKjfIGgNsuR569BLpCpRAif2NzMH7EutjEyqRxnH5Dz869LWpLI3zgCPdKgCXlPg6HemZW8t
EQptAOtmaRbt7P1IGce2yXlH2GMbt3+dWw8e3LSHbwhuE6/RmEH0TbYkBGvwuheQIb2gbRQeOE4A
02dERmM6Usgj0wNSE1vXwyDLG+fGLTydR0fX2TkOhyDUtdBQWsq9p77urPdxcO2qkWRcLrA+63H6
8LG7PD8HaJIadLZOHBaznr4BZnSG1ITwhYLkUn38x+WaVBwh81wK94B9UVQt68EmVc9AYZKzpPm8
p6kLUKLCi2G16dn0CPuoW+xQzHJaWBUQz4Iqu96CCg3nrQUVtBhD/Zt7D95+yXdk/2W72wgdwc08
9mPcV5vCH2DPDeMTR6eKu3nvIJqlgtE2YGIPsJqIXUKiy7NpbUN9TNEcTRJVJPBWLpFwK8foABOg
1lTEnG0ab6n9E0leoYDmhpSq8Uc/hcSUvDX7tdyAQdk07yl/u0gI5wbphhUV+tpVs9K8UZFCpa7S
KRZuc931iI+megu1m5Y9fey76mFxq6TKbNQu1W0vqLncwnDKm2UrEKLyn9e0Q/KG9n8DG2wd5x3H
7416KT5w9y+jPWYYOb3AzXSllBnbnKovOXuObYRymkA8QfdO6NHpNHVMbjf5V0E5ldxrpoWhWjVy
Dl0HVxxZ0usneiSdzz4QVlNYO2+HSCDzyWvsSPKTvwcaxXR/c5+DHzTuBbe9ddCLc56K3vnsDwNE
i7QnV+ifBOqyBwfMhTc+xhx6ZX1EQUid1EkxIrA6YjReGCHlVmCUONEqYqWHyA/5OO/UoJnPJxiR
jpBMOAcVE2Aa8/jQEF3Y1l3eQdOinBY35qxwwG6xQp3YCGtu1DMYeX1fgQd2HVGS2J4k18vnD64l
PFZXx2ma5dIV/YXG8fD7I+msom2C8Hw69HexlXVCle7EyYDXp7IS+RwKy35n3EdkRCBpkJk86PMw
Bq020Ue8eKBo5igSbNbGXMoGFoo0zB2Z7kTXYaEN9G3RM7lqNGqXxrkGg8zAnjc/9xU/QgKAtR1v
4VGMe8fxBmwbit1VFTScrQzPdqHHfIxYlo9rzOC2zZQk52d4CiZTGD7wGBnUqm7PEYvm5BXPuq5U
IhGnwwrIkKgn0gJanNsopufK/lBlNaH7gmm8Qks2MfgsM7y6zjn8Hh+WIuiABgc8fuc51o8++ybf
D55NYHq7kUFEpOa7vvkM5omU8ydVLbSmrcWM4oAGHVeWXbRAmkXysXdjP/pun6dJWGEQuAFksOgM
9tnfs9wnLi3qvsDzNIjYuMNniwiHecrNV+jGlAKSnDE0+uQwGVW137+Z5XYBVUlVu7lHF38j2xK+
RyvhtzG6eYcA2rggDyALyRXlFVAdF47fLgKoSPWDE43nEnOcmRKFCr927x8r9/yEd1zfRZXe9BHe
+JPDkj1DtOlzqd0BZ3yD2KdT8y5j6IadUQg9MHdHQ3w2s8lJGujnDgklfYyVpxbIlFODsyjsSrTs
n6zZrD6XKNZRxApU8fyzBf7LHg/l78TLCtyYROBZIXw1HlhK5/FIM1cMSODoK61zFCB9zgNpTeOH
yOStGsgP/BeBGQeqj/rkdyBdrB/zYvHa44r7998FBUqTGI5JFVwjbAZ/EGHzZFf1ooAVGysq70me
T4cLJb+i8bdVXKM08ngol6G7KjUMOWzR5Uah/iSk2ZLFAuYt9STmz61Pfr8U5IQTGYTzetcS1Whu
yPtgV9D7+ePTU1FR3zZXmBSx02433atY7jnDIQXoaz44UjYHqkE7kTVjARNNrDGmxUU2E36pb9m8
HqmzieMQgZYj4IaDT8gArI7pF5vNdTSW86Fnei06TfZKdbu5K7m4KKTe4KcdafOQzuLselOB9gq8
5IRicXQdHS0bePXwOffwzhv2rmKJcCovs/dYhGh9QlarxkH3johx1EjpsWTyIvbb2plyK+d5ud2g
yo78k4z9igCFXxyw6EiMNXl0BeQs9n5iBIeiB7oFxvHZsoxVR/+zPJ4DLc2tw7SOy5EUL05XqyQJ
QwQTt1gTBWBXnyN9G0GG17WMGhWXk1+4EW7f9jyI8CkROwJkZw8LyXipFwnO/3okmZ09pLIvr0mW
fe8nmP8NigWIbB2yRTjrFUzwPTo1ClNZ2/q9dV/4I+xmHu7B7al/yErL18le6Mi0gYeRq/0E7Jdd
Wxq7NkXeoMlLLO2UL+YmBNxK4dmOfMq1oOXnsvnEzIsn7oJdbF4InTl7YLo/4HHNAUGvAyt7dnIh
LjZQkCZCX85x2vki+V6ufzoXqmfPQJIW7HCBz5tw+aDnSz4vq7NIQYuBzL7EajAIpQDTYTYZOX6p
3ZlpVrlu55d7tSIBQ+1P0/5dTlPF12NKe1i2FLlI9Q6zvQg0pgVhwrlyKclqkZ1QOeWdVGCq+X5Y
FoYdjKfx3wh5p9/q+rgkwJciy/7E/F8pmGmbfTwixZJZzGgY4puxAYTvoYmZCynkgFdN4dLGnso9
UrhayQeKBd3EM2FmvIRXUQaKEkcYLy0QODaKa5Lc2wKU4b8/2wbmuFsrcOQMbMgP5klbf1s8fx5m
I9/nijGPu1H1WuToceGdhVmMPBNTwkXRTmvSutd1aas3cathJaOI7dKSHP6XErvTNjNH5wu+Xs/W
HPUaZvpDe0w5gCAco73R8RYBIijt69ZwK1LCR/y1Z9wFVXO1sqm96YZEVyWEDtTbrQGiao/Wj45n
ML4c52wRvwXCKleUOoO/Y0tb6+LrkJ3uAOBgKQ77xSonuibBldiWUSZXMyrpi1ObR5crF41R9pwU
bz0gaJ4PQmloze80AXYyDZq9L4UxiaSHu6HzO9ALtSemDeNclLL8fnrpjewTUZkHf9uljFFyqTJ3
Hgy3ykXwirU/IEtRxHe6vgKsXN8D5tZ47xZ1ogRmpYWjkC4X7tdoSKicKnsMylvVEf6pSuWzU3Vx
zi9P6SL/gD8aDV+mr17BHvqoiNDp7pTHcyGHUEjOSjGctieVZ6U5JkWry3Y+iVIghtzDKFpW5bEw
TOeHcYwbQLPxJJVHBP1pp5unMmqgk2hWbwo/ijasBrrQgdMsYL+P969ZcKuhbhJwRSNkZgXW09L4
5RSBCXk3KMkqaj18MqhvHj0IaLG9OZw24LJj04PGWNO3xHsYLfrB8dnRlVmZ806CHzRuLiQpHaIb
S6XFqXtqjYhGRunzPtFvSQ9BJ3phJx5tjA3DYqO8ktkas8vxB0iB5NEP05UQ9NLN2Cbw6IB+0N8P
Rcg9m/CR2JZfCpAUtzsggJ0rH3p+qD705qQbJTnFWG2vOhI4zoBiZBf5JoDuYvHkAduROZgg/vtc
tPneRxlqcN0ELJBeLO9YL1NjG7kAR9OXqJd3OCkbz4y5fT4jf0pEzsi1caRPUN3XWca/c6du8w/v
KWyYJC9DNkvLEbBQsfh6TuifF3OVjLKPp2b+ejXo+z+0qTa9NSEyn3rsVMCTHC8KDug+ypJcxRRl
YLqJ5d6/p+R/RPsvwO0ZenaPqKruQ7Ecbye0qK2Q8qxKuzeIr6ojdO/5yHPWPBRcZgKBfgxwqDOV
k69Z/L/ajDo/y3VDwjrpevxMvhOqnA//KGy41b/Uc2nvT2YqrdVAVfs1x4IK6LWEAVR0tZqCUHjI
lcH4eH1EoLdomSlsl/XU/cR5s/VWqOpcRQYzG3fAH6XFCQIm3reO9b5oA/XZGrI0Drr3RslBxX2f
P5ro3w2nKbmoUdK+uJK/nr0PpFIEXKqjVd9r19K6HYJ0ROiVt4pXLTuF8GhpH1FohnZU6DPpAw46
6233QJ7FrynOOraURUG8zth5ag2kvrbil0S+mav2hVv7RU2R1UlBdd5WHDIpw0C0IQeiqbgLXaTP
B0+KcMnrs+q+zJzxhdtjNwscXAnNu+gWZ0U1hhi1fGY//TLfPRfzUDv3Sjqw8V7TPKbEv7GkaVpe
UB4Jk6Pt9Ghz5maAi66WprE4qmMA+am+mP13lOIZwOrsDT0v5TAI/So2h5MwwHuZJr3TfTknGD7c
BZz0QSmeAFC18IMbLz7KJ4h5QG2u+GVrCehO5+S+xv05jY5pwsbE/2jyGZxIq2T17+voHMQr5KiO
Q1l+lVD0MfFLDTaa75OLkdsIgp6zCBtiWIT9Xu7Je4juGLOKXRQ9WvvpXgKU+LBG+ctIBgP3yBBV
1RBJ5yqgdA65PedX5wNQOyF9KrD4pT5zE0W2ZerqtB5fk/+UHcV8L7s8iEqjJJ/S6tfNAXcCe/VN
++Qsj5Mge+HDt/FGrfZkqtS5gOLoZT0qbGGUMxdruqTPEHkKcGpIBcen3XkSjmqCLeEQCX7lbSbH
2UzmW1TsKDmsHELW/BRzHghezOLkyPcxb7OsGfpdQYiShWhMbyzIH5cJhcov7DYcVYGQbTBJDf4j
sE4l9R+HxgMAtWQiupFo0NhLo9NKP8iFiPHAV4l92qoQAMIHVF2EuL0FIm6EHfsag0ctlS3XxlYU
m52Iwqw0yx4pO8UjYCVVULxBRsReV8uU7RdzydM/sPu+xlte5POSJXNUvuh42kkmfZAcg29eWMmQ
nlnbOGQNFmtpmWk5Dpiz3hlU86W0QxqW4WSp1v/aK0U9FZ/RiNGhPKvxI6hfh2lmtfZbA6NXiSSG
a2HCoW95ZfJPpauhrmPWhfZX50UpbNYklz+4B7Y+QjoaB8vYB26E/Wuf26AbqL9eJzN6uIrHq00d
0IThHjpSRTNOKGw1in1692SILzoje2U8S1HwCqHs8EYa9eoxkG4oQKD7qhT84R7TRBfESdHHW8hA
OQWwvkPdJFPKjBSU6SJMNUUMf9//mZ8fXyVcYiiHhlf8BAJKBR4VcLoarJi7JDbSo4EXZFy1FFvj
FsgFDLgjLOAtgFBJzMeczCikpt1pomlMcVk1nHmZOkfA/DjiCBpuA8LwmjmsKhLVaG8iv4g87VVF
UxC7+ngboUy4Hf9d7JItaG1wOsIQNvWljXgghRm/mEHgzeySd0i8Gr4LrSYBn7+EeogXMFPlBdlD
utHUN76dtAf4QbIoYHKpulTIanq2gwtkus/zAXKzt1UrIfjb302Y4DIn4G1fvtCaC1xI+NcpEIde
ykKTY8dQblRERlfZ5DriMgRuTQAHcNZ+nDgzA0i+DsOJc9bskLQwpsc7hqAgD3FuT+M5+ghQQKMy
6IVia4mFQ6niU9UFdwsG3zkl/WVhVQMX513jLhB3rPxlnN4xWK0fzMgrFSJ89ZR0k8LBWdSJc96Y
dNJ95kVjcyWwAGTxx5CQq+0pe6ig4+ZPlfJkHSMH/RKjknUsOQ1PDyE0vczm1dWORhUcGhQvAaUO
dDmmwiQ2K1RxEwzW858DoV/Hfp5wCrZi0g7rG0H9ILVxKJT0waSDDvFEP8UzlTYPE0VTnlVKdFHO
cRfDQna010lCSQ8oIcFyrUaiTjmV+24wFr/mkx8tiWi7xZ26oD35r8Yme3fxh/4YD89sO0VMg3X4
9ooMFdeZozcJ7usG/Y/zPyznOq9YidPuc1geQbIwAvZdOvornfvCGMjVrkQF9ru7s+pYqXv3rtNw
RVACWHkJUQ6kHhRVLVGJ14r4kHXstJkM61lqLuPCJGtYaMhy6kWibF0vx/SO5eCoAl+js+8mvj0m
omIoJxt3QA5VvqWdXZWngj1U5NG+SUc19ebpS/PHx0Lp/OXGAnkZofe5O162SbGRVTS6wFme8CvL
V8NIM69s+XVZKKg153ydUMowdgqtXDOZPsuRjsXs95SzhYRsijtzXkf7kt8A4CG+f4QuinTigy0C
AgYl+4talyXtO7P2hiKsAlq4wVXGjbTZ9fehNm94pONsocDiS9wblUF2pX/c6ML2le7OrEk1x+r1
4pPFTM8E+agmSz3YZO+sRQ2TOFbHnSakIiStD/7BOjAonSs29i+eaYegE9HFPACieF0FJi9exOXn
2AU5teKMB3O2eg4KyfF3ZGIeajzLHda5KIYKs22pkZgcPybwOupg07USau6ffd5j6A4Ja6ZfMB8v
dPUiIYFBAnlsnFwiEDW6AH/XpccKMHwD8E+6Gpn2PjkL8U5WUeTaCNvY5A6oXZ33cAg7yUwtPOJW
08DjiqhoXt8O49aZ9Z4egKQnQ+m+dKFnfvnR+x+xvGMgASepLEkKHk1eK6bCC3azx1rquiOEFKh/
8Gjtnll/tIhy9HTabj9Q8dZsLZeQ1GflRR+wc/bOOmU2BtHt3tJsUC5BMvZD6oaUOFKNKWnQ6dzK
zwIe+CnQawU/7l4V1pkH6oay8OxDu9CvbCm8/55Fi1YTIVvE8urS3X2W5dkUAjKzV53+XPHVNJbZ
qO0P7QiRp0vcJdUbNhl1l8Mmbtk+e/t3xqpQPsiJD9uw5lzNsLcUPy0xucizqMwkC6AOyDBYWh/D
7kxdW1GmbANBMRRE9Te0ABg5yxsKmukuRfiH+tOSVPAcRSHiOErTkqvVaOAIsk0Ec8tOWqQDOzYw
TAZxBN1IHZXU5yj1fGSppErMSyqMV/pUdHujpQqgCxjWRTsFPI+ukrMB1ezWi44ijnBnDtPSXy+e
ssa2lXno9lbg/ggxHFgKBus1acs9C2bgTJ9H05/T6Md/9O9BVty56T7oFYy1KLzoZfroFJpd84ng
AvYQOS1lp1kThWjHau9zMf8sivP7GT7C6Fv/M4i5vgbLO2APvt8EXnQZJDmQcmc9bHp/KZBle4FP
DHSEX4C4GrSnEGuXEz5SHS/c7VplwWd2sUCVH6CdETIN1oxNaRsadXYqrYkDEoa1RUrxhpkW5vVC
ODSD6Uy97huZfOhilElZm2gDdmSnXWnNPOh03pliVsqDi+wu/i/XhGhkdSsNJKc88JfSuakIAE4g
XWi4iTCXGpsG+x0ef8hIbmhH7zhoRIpT1DG8GTSvh11awllHMDRCnbBlUoeMZ8BV0q4J0MNxvTP9
pqNgfIF2AhpgGveNXrJ/y0Qsek7P97bg6jyxGnJrZ8m5pMBZUYw3wrvB4H6NIzNgAGkS1Mm7sgdt
Ej0A+/3y9ahFJ+qYKDgli9dDCkuy/ulhoop9aPRGZ8cG/m7PDwG9BQQEf+h1KlKfCeODLvSFIP1n
fBnl4U02lxycRX0mOtlG6OlAdIa+CDYN3uAyIymLq0WPqBR39/WUvIfZt4D7hCc8iGJEIV73lCSH
07gNdC/lg0VF+qb7uGMpLnhBYbAVFTImVntNqFtkvtAy+3Hdit5YEbeG1AiHzhfZYHJ1CWI01K5n
wlhYef5ghfzsUxsYbBbaZP6DJ5gyAle6yIjBnBIXPuxSO8tgkHLbvcXxporwQP8QZnNaIWkgoKVv
RZFKkfLjvoVzXmkAsEUKpHyKsIOXfRhBQAYTT91gOdJyyIDV78EIM7G9JI4DkZBNqc3wW2D2JSzh
9UwRYevkHpiPhTjxeTEDARB2C4RTkJPJ0OUGhOkwopus7TeVRqNMllwcgoaIPumtT/1jmne9KJpp
J4ih2Dq3PM9S1zRID+nNLlDz3ZWLKxZjIgBXgw9Zl78IJay9I4EGBGxPJimRQjEisUpxNcGXh9n0
jE3HB+wa9E13N4ZZnCpASM/rMi6YzkY2C103qRTQ63zSGZluiulJfEd1VLGbpcAXiJd9vy/IcmTu
f4ht1LEENaBvO6yjKwABwbUEKKis2q+Nv7oLghIJPQzpTMk9oP4P23WXC3i3pEY8FmeSfcl/HqDc
XrKh+QfJPeRGk+IKxGgFlcw0wEYzsTjawqSpnpDzk2lv1K0GTwZngE+Gk6rYY8ZEqWWh2hKGw+1U
HRRRs9kSuEYgmbAm0qPBvq+2+XEnFtfX/A/DnSsSgh9qLh9aq0AKvedczQIDy1nNmESNRkRhctWH
4mOhnaDNeM3j6ra79Zqh6wjZfq8BkTAxSrF9Aq+Ok3ppI+5DBiVru+uXK59Crhoegqo1QpFcupv6
gUh2VTLWvjWemUSS0mJCsMV3ucLhaxub6b9GRnsH+jZUZnLdzbI7YNfRiXk8vx1UsOZtr/h5UkJ9
Gi5+1IAuSR7dmOMqx9/gxMPDXYwTfKNBuEpCBeSK3VbERdtKx6X2weilaxun1ofwlbHEuQ1LNLdE
GWKK8Omd1BjYorSB4WQNw2LQzxyN5U4iKZzQM+2zFlmw+wFWqRBHVO5ENsrU7Cw/IlNhFhKM3jSn
bnHjN4B2KtVYk+B6yEttmh1EGFLyxqBHeE+7IBmwdib7vzTC9r0NC6ELUU+DN3SxpdUBgx0LFtAR
JOd9S5yUKAYcy8L7w1DmlS2blyJ9tdmGMM62ROBWl1DFipE4qeFvqrkNA+UaqIhUY425Atddnn6T
TayfRcAEyEWlr6IoDU5p+7dQmmc+jDqEV/dEHTIDW0Ii5mjcilRHosq2tDZX+w1FEZENc0NR9e7k
mn7Gkp4rISRWxxRo0fO4F8gzxa8AuhujO3KHLdF+c6elE1VCCWQrdJCDN7TG420x5IR+h4Azt3sN
GDdCC7cKKLcqgqG0WrXhOSGj9U+jmKVL0sUOv0NMG2CjAqUHMzYtM8NCka/SRNtiNlyhyq+zGDLF
qG1+4biV1+Z0UKsFtLnLa3LcpW57kBF6+cXkyEcuHHJ8TZf3jNBoijGp+GYyvD4Fqu8PI78ZySCC
rRxKRZN0cCzhf/fFkiYi+rtjfUwNJblALpQ2zhbOi0EGgQaAJoXYYhM7vveom5AoU4Fs1o6VYr/P
aAM3Vyfy3fiGBeZhFsxi2URYkgfZaFDDDE5YNkEIb2RivoHcheXBL7Cn8cO0nhe+F0PkaUT3U/hq
hOWe+ytQvpsrdeQbB9zriuV9JGMsW0m8MBp9aJ7diq/HExpL4Ts5flfO+TSnGngtgyr2SQh+QZlo
ZVqBeuQwiY+GaTbLgLWZu+lWq6UfEJjinkcNpdMByUrGE0vC9xp1jBgN5U7hVJ04ZLPfD0J3tnoV
SESlbUkXe8HIPkzt47Q1qPPkI8AM1ytU1+F4q+7sOMxs/D+qVFyPP/EkPIlf9rRQLTNOdHWp0oPz
+H5cr3r7VKooCxMCFCP8v+X1pp2A1n2ztmK8YgXZGQjHQPmNNLVMAq2B3lfR4BGlX6oFjlrYmsn5
cM8OfdqB0/FI0ygJUY2XVGly9XuQhNS3HtT5cyG2fg6A0Ytqzb4mTSgXE07jXwHan2poDwEafL8n
TfL/tc4Wv0j9b9aUtTzAX6xV3pIhdkS7msXYFG5EqDsc4JdwEfGa/TwfmO/JIvFWn8everPCqhaJ
u+apTglV9JoO/Kf4O+G0Am2r5kC8Hr5mClXT8L+OFM1QXJF+y6ltx8raHQh+ET60b52A/OQJwXSl
q3pqFh+VQS0W62vt/PKbdwFA87AlInhiunHDPN03KGmDmdqdTZ5oZwUJeBorhYO4D1p7Yz8JGTuI
r8cDRQGxDY/vmuTtNd5/MogCQFIxtKdfsBmrfdsoG63bRqqzSKdWSXad7XQyh5zLGMg9PKL9MFn2
C1hMrtkO0/lHyOGr/VwVfYX12+jSQLoZrwXXyBulTflAniyVQTeLLtMpqzVaD3y0V/bvQOK0lB21
ur9ol7OwL8uS6CfdvJ6sO3YnWVJjb9zKcixKZf3X8nsdgRzaYkGKiWS7VnM8IyIOOfi7c76fe+oz
Vn6790K9+8NRR+XkwE5uy+08VNQnyV1ECUSFoF72axbc6gHJvXI5Fqe1+0N0ZWNp4AKuW1LUNUjt
/GFrnO1DA3HdCOjKhpOIs9ReS1lwnLUUnzRRAxvohRRDRK5GcDhXKzwKVIOm2SUQbZ/QvOpCUWGF
5ZtP9bJYK2gmpPFdiU2Y8p0jn4YJPprt9j6XlWaXIyWx3az1Gr4oa1zpqt4NYcvOp79XtcxIRmG4
AfWcpKeaAT3x4qhRMIOc6RdGbCMk7LeExnWm2DFm2CqlyfoyxBm6YkRxnf6QsuyIE68alTRp8nNp
kcyHYv6kloJe9oEYDR7WbCzhZWlO1g/qnJTV2glcPkkhCyL/eDisU4yyTiHZtG2XENPzd0f6FL+H
H9VXLbebsNAUrlWb+DSwB40q75ZxizxK1UE5BBvTR0Oc0jGugaW2xrNqRqBRLPX6Tt74gMltydgW
+uy4ZKTgSqACrep4VDKlYh3QzEULpx/pLy8Vy9UpUfioYNNdoIjElu8EzzvvQoYgOX9X3X5FWlQr
ZcIFzq67p+ltb0o0Xs3gFaGiGOlJP2X/qxrU5/42Bf4i/DPh5f+I0zGmaFReZG+7RbK5qgW5gBg4
l0VsOqVIthBsgPc0NIXsiIYv8L/Tt5HVNi8jKVkfjwVBjtiubnBtOWY5U5wOdeoBA9b1BLsYURUh
yVGemLgIUqEJFjVuSZzhalo1113vUreERtyqt1FXQFmrDEHj/M1MqbWVgdh262xb8C4ZWs/Kh0N1
iZIdqwOfOTubg7AQmOOmT250xtypXOKbDdIbPYqIab47Zr7vNxzP9PwwzA9Dmp7rWwbQ7Do+SF26
+8o2IxlCbCXOXRxwvOl2kDlOPMVLnF49UlhFZ5ae62VaG/IV5OPHtriJVS0W2Ih3OZhoKb0DQxwp
VZwI8+CdmKOEaq4jZAj9nvelCnBKjRF6/D2A+ldywLtv9GUbZ3qNN7ZSz/tSkeyaPLMQ2CDDRNAo
Aw7qpQJ1lSqzMQQC7U8wL4xrh1rqL6di90pY4gFJ+xU2YRBW4SqOt0QYDwHKGZRTDUCA9La+IUIV
NR598xIIYJtfCNcLWkWbreEuPXEFfRf2ytMxvzKB1aPLdCbO2nHpsOyB3i07RTEvrPBPM71Uel9Q
/EJcZ5eH/u6pWGlWkWb39cnCHpPNDewMF1gQianX4YuimwMzVyphm6UNZSQDm8gP9wFwUdx9nx9K
KKZa6fdx9TaH4m1tOGNh/wT0GjPRMd9g3iAqCJAuuTfL8+GacEY5OQxy8Ujy2yKWwLBuk+vfmkIj
7+1IVTvfMtNT7m/q2R/BO3xr0qKjQrMZUNNiucXqIDdqmBkJX9U9M/nH/RV2FiN3V0D0hmpJ0d94
yOFlme6LIcCRqscWdoTnU5nyL7GDX1ZNcZbOLIl3j6wkVBYgU5wI0LLunco0bvNavpBD4+JGGV5j
0/KDX+7BqzlJOzCE4er6FVcyZO6B4CC3hcIBVe6999c80bHeOpfFRM5Quw3L3lYK4r8XZ5iA1SLT
gKhZKT73WUjiyNQEaXxY1MyRHKA2+Pxzu/AGyHHCMXJm9G7yGSwFLs+cNmyajJsLSthu4BJBA/y+
rTi+YtmAioVAQ6wVdVjjFDjzaqJJhwPHt7ftAdoTGyrRNOke8vxTxyffxVKLO7vICDJCfYP/vVHc
b7Fr3eofT6nxLS36Yaw8cheqVnzJjCnARwZZfXc3rILUWrX3QRbtGSAz+2PIB+s6gLDFCwblE0lN
odsk89uV1ZWUXEdIqlV+bXAmwTx9TazWqmS1OSNDcuB+YBh/91I9xIWEW/HCbYk/74D55i5Srdst
6gA/Ubef4tVGAJpVwfOYXBFn80ZILN+UUKCPQ2Uz56Mt0kg2EzTGROgh3T9jK3Z+2IW66S/jo0ts
MbB4d4CG6UalthZQtPJxRVjMwmMojdwh7jlGOlw1Meh9xVrv/qWslhO6UFe2/7rzIPq9WKMuIDY+
2k0gQqGwpjtZcSAO+se0V33lMASEwJVqk/mt6et1/BUQ/JYbGkhGBctOzpfbTzlKgDcjnhzdSwiq
7n2vC7Ae1o9kCodvOSsbDCBXOU6MLDmo+4SOZppwvbKDbGvXtG6QYwoHnT7XSKLmOa2KgmoJERPA
JYB1hAHlonDoTabMgxduM23zrPdacjtPm/CzOjXAwhhCHX4D9nx2eEYIgBFyhO8BkJJTxVeMyYEN
HLXAebQEuhCSFXxTd0rzsjLwLq7lkshMSEI7BdueiecTLiKP9kc8Qp1YTLxmlkHfWlMDa8zHCuaE
f73Wf+TN+ELtBURxd8rEbtWd1airmko/zmszhN8kHGYTcuICQCAW1xCrr3cfqXhmjMBZlzQpBVUC
FaLvw4PHuiT1fJrqdDlgjJW7c2/C8m9z4PBglTtXw1iBtd5AgoEqNp/zMdBlwm3x5Qxv9M2peLc3
4BWj6pcBdXabn+wHxbdzTysxy6j0W0w5xNNaoTjFkBIrVY7kafz3bgFtJao/rzW1JT8vQ1YWrs2+
vHFFcsToIvmfCnf7/vF/B/SQUiHD7e8z16E4WiuaFPI/lH0zYmjof5KNVkpzq1kWXSoYZPblmHqu
NQo70gHByyl2P2wNBPE6NJtNdU7wKQeKm5HY+wpOKICTm77XVcXlC9tNiSNtddKuXkT1W/T45II0
wBKZXZpdk3TuO2YnR4VGToqvSMh3A2KhIdtn3xvSZCsrKXgHPRqJfE7MSfKu/7PZZCS5pVgjz7hT
327BL48ws9GPDZd+ZkMZ1bmeUEmfWR9FARxCLR7m6oYyK4cDz5KGsD+DDsBkbSh5T/8SoeA92z1C
NoQpyXHTPcKEjo3AIzUN/gxjyNN37tvPd/FFLtg8jC19Tudgv7hkfv1A9GYA2bNjdBwrNTDvsT+z
sfpANsyEAYIMMO7zqxqmlDSySLTfObOj/1Pya91PtAAG2W+bphNd4B/AhXak/soYOgJ13bAGZBZ5
NV++2Ze7aBD+dA8u95bWp5iadTleulOGLmbqp9LyyTUUgEDOk9NffAEH5x8BHiUxbGxxA+XQPhBZ
Ikr2VvvoUp8ADH/GIpn8/DJm+UOJK1JJJ8PcKbNo9MfGsX9aqX2G98jOEHXp6FLhx1AQZfBEhL0N
cNJqL2FBdQX+y93uxNjeZnfsZBqd/yVpskZMucCwEiVLiVFg77MbytjL+DSbpWOdnyQ2yUHuCyWr
UBFxiTVLTYNSeW8gJ54bGCFgyIldu4fu3SsdgaNk3uIfyoTq5PvGKjiPBoEao2drWzvZzs4y1uSD
oYdNgMVaOXBTSjsiL10GknKEpqIAComSSViJQrG0n6RD+Pj9cubOZdW7IGCUZrD/7WfIkrJ/L1ER
vrHPrcvryZxb/ltVkS4z2KXcwbQlKzUKqXC9FR9jMWvzK6kRJno5ksCJRRwdryXFoBX8+pMgdp+x
7tz3Y0DC4mpqIcXujMjEdQeEsL+e+um+gyaO3x1wjBharHKRuAfYIM0hIrIrmQXyJO0i6QZogx8/
NhmeA1/nl7UHHMfC6uXqMTcaJ2q/Fx55ind8S26AIhVouuM4BiOYTwkrOB6BWZ5YsGF7+5s5+LnP
bxETEbXTOymu7/5uzfK2c80jEUjwnyrO2xDl3VIOH9K/KCGxMKuRy0ukU15pXPgBFR5wF5yfzbTL
6uLDzBGeE4kHuDk8G71xCg3eQNoFF2SFkkXgFXD+dg3MtUmNnKnkaMjvjW4Hf3TetSLVx2im4rBr
KkrhQ+BPO712Vl8hjQ0DTDYegdb+r7q/8Qgqk28PmTFAg9DXM9dk184lY2IoMRM9xuyICdAzUUkd
fdVWx8oWg1kZahpnqDyeOyyd5Rh6wa1EZzr5g5pVGyi9lvYZA9xsT3/4F+YMjT8hMYBDOTNX2x2N
Dy4pH9eqV1013OkzA0ZGKiEk7NU3onJ0/gB5fToTfh/ZRmBcfBckumfx8PSJOZAEU6htDOM+ahFE
3DP2b2ePiXfV8cdl+JOxupOqngcyMMELIKRuz4ZNjIZ1Q8B2UpBso59/m2oH3LRM+jzWJrNVVgNc
N9T9ywQXX7uJ1ii/xPBFo42QYhX9wRbJ2jcJimpwY7WPrGMqZv5wHhBfkhfoauI4AaaIutN2dYyj
YbXGMJW06McVeXHJUUC1/Noo5e94aB3t3kb1pPFWlLEA/UYTNKNbaNiYVOTSht23U1M+I0qYVSk9
P/VeRlDRbrYnRXJ1gHZ2+9XSExI42TF+3rkatgKS+8XJW6wjKrGSJFJnlieveteEhV8IgakOQ41j
R/qrRP1zrX/0AmjUKueX63xBDeKJlXow5/R8E/MibeFksZ8VTfNj+apxk03W0+YaHx72khoweyzz
BMGPs8UHePVeCIT/RQpun0PEr7alZhmzBsr214nFl+GBpBB/Iw/5aIKAo6CYlJ0SAdV8sQgjYeqk
cJdbeq34hZJ7GuGOhDYQJHuIasr/03DEfWabz1YDLvKUoxYnURsK8PutXP6sOenwAnZj0nzgI1aa
RkQa92HRtv8g5WRDpp7GwrYzKocmaIJc98yPUiCgnlloDhsYbJybZHId2uvcqVIgJAfD828AiKJZ
Ob7+WDmB48oGn2H8h6ZQVv+dtz+lT/RGGYfHCM/2V1KHBpdHo2nXDRBx0Rz9Tl6St9q9QuZqJRTw
+mevUTN9jW2HucyOlmHuV5aULX1lIjZ4B5z/XVdA6I15198+xSqSnAF/DQ3zixda57mxZib4ors+
BILUtyKriKYzmvG85TTsWW7qHgbtuII+RxAuF/+Qrd3Y5zPmcldnLVa2ika6DifygeYAXVn6RVbA
agG38YOPy89wFcd+EzTZVmBvECkWnBggaeevFvg0b3On2ZmfPYxFEQyoORwai/M11k1ZPPl7i9NP
ffr8aEeZeMtKxw83yrjpfucC20jHUo+qeEvkTVOR6dJ67C00ffcx08n714KXTYiB07wLZMca7Fwr
93EI1DRFJuU8B6ejjy5SwMisKnXX0LOTnuW10fj2/ziAarbuydAHrDnV7qE/pHaVsAJZJOLbBqqQ
ZvDddUGLc+kcabEg50JuP24xK5xKVqWsi3AWE6OW5O42pC8robuQk//B37NvQuMB8zZA+FPEVrjX
qfN6/GtGrPo1YkARX0pC938wGTExmspc/r1Q8Yp0kg010k1+IZC4FDfrpSSouQAaK3YYYhLmE4vX
X0lhdYBLxyEmj1M+Qhnh4xi794qUcHJL21SHifcazroGEY0FUukBqEjfYqiTjeiVSaggvQ/M+1I0
+almbIi4fhMEuJnOZC7zcDaH9GlGKG9d61cL2UXmfNwejWJuUwcfH6rFZQKUKFn6sLOGbgksfDJL
nuIateAsnrpzsQHuvElPtpKZb1b7oHeX9BaJs8zJb/zxypeF8bsWLcRclBIseiExHSdKBkIG0oYn
E99umJiyAoM2ki+xsClcei/YbTgbz6fXJxATStc6Mpi64XXRBzKDm0jS0JsDfGk/X4ndhZ5jDQzh
OtfxuybgGoefut3Cu0tFXphcq7O+SNQKTfDwLOkvBNEMJMXxo8Q6XRkowcE6MmweJ/GfJjuHBJMD
O5iZLoQORQXbr/lhskrTTClMenov3zktXa2LyYXKI5JACE+Kndekehg7qezT3mG6lEzuXNL/PGPX
vRH1TsdfS7/drZoLG7IPLwljR+wd/aZlzVZkkDIuvKC44W/JpnbyKwhxwJP5btFFHJ8PrYUklzDS
vjfZ5AChXRDWhm4oh8l26actUpCU88h7S8PRO5XcIG9KlDDhqfzaMBJrBX6sQoxpPAYlr9xZUGac
mdu6ixnHTGvW3pVg5pvqTo6axLc3eCsWZ8l3vabOKZiSXqSDY6Oyhe4z1N9mqTQUgtsuMOGaqu6s
yNImmwieLKlwyAc7EpJOcgQiaLOU8+a/bqIdWT9E5azPnYhzY7rUUqmiJO1nSDukKmpu5ZRpeLwO
t4w7cOJ5TGY0ncFQ3i0sKlbT+WyW+ekvQhfkp/ouAiEIsZGLAcxQQ4WMxfQlFGni1uu0Ol64AwXZ
vLAdMd2FAuFJDnWkUygm3i5HiQfWs2yS1wbcn4Wj8WhTEpho6NQX7iJabs0hrpUHmDnvG1Thhx9v
ZDQsHw4VMKXALTYPNHj/MJFfl8J59mkMkER1EW0JdHvtX9vBOpeLrzSEFftPm86OMFNF1yGU3oCD
cfV/n0Uj0AE9A8oP4bdY2XRh4xkKuPPTb9dX1+HBctXqaBCjv1cBfIz0TnCe5tA9rzwCZUrmucLD
+CpYIbwaxFlwUXxBMpPPka0OlOEw1K3gXJb0kWj1NmM6oOtdK896HXpNcCdMEs39IRMjVb98wXku
CMOn++L+c/uPQhYh3a1HdQb3XkXJt94erLpAiDebGhrKN33cLJjORR61DSFylCurmIMWFEvSJs/B
uOxsk4AaySB4cPAFRdKy5xLV2n/zStxKlTzF7xYvVHYQwleO23bq8pyMaXX+eP38oi7vzQ2S4NHx
vIDWzpJpOfN9esxwj6wJVL7vTbEjvzchrbAtUPRGbmViB6gPIo/R9fRZHWCcej+bVHPGDzZgWL6D
X8YzNu7qsSBcrNv0rrOvh/Bys5L+x5PGxjIiRH066vVTi3h+3/ZJYO5YDMZoSSLxY3y/0Ff54xLt
hWS+lrXbewYoGy+lqXTzr32ZhJuRxEZlPQ/p+YEXEbbDQ11HYG/aAlckk2Gm0VaAJpoOnfLmuleL
xN5KP2M8e5pWCJjzf4gbrnAEkr3jKX5SfnaSpXLqUEvQU07cRujGYIR593rdukMcc1Dr+nvJT5uf
Iph4i66Yu88QVoeFfzgpN5qw3pv6UJ/6/99LBsM8rYaJKY0UfLLmLF8dElK1I3jaFMQ2pQh3EnAc
+v629etYDUZmtjthcWPs/BsRjInLAcCjlIZXsmkUbasKxhEsK56fiibFZpYiaQHvsMrX80L0d7jM
grKcPAKYZ8gs0taqLF/nan735qx2eje1zMQ/Kjj8DDXLRF3CTTdfiNcuXZ3hXxMh7NbrnwR0KJMq
rw3+Xr8mMoktmW7HJi/CHkkqOkrCXEQh1Cb/dPTb54qV4xZZgwoTrgWgkBM/HKAdZc+wBuqZbMHj
QYM6tbDlQoDOJ+hu2+UkjYEMKe5066GwKSi1dms0YSR8LY57/wbXIaUXyHkc5YGQLaZnhcW3B67O
+RWaj5xL3C4cBfZMqjQgMMDf65GOcJ4fVMF8nt3V0mh6AJd8Z9QOsmJaVgmRpr19qRK4rXaZCTWs
jt3+N0bvBWnxeCixWAG6ozyVM7mThn3oU4Rbg7LMFsVdTyevIkseLS5LOBPDhhFAVxzdM0Is7pME
vUl18ozh8MUloJObU4gxFVnYg5WrSgKrrx1mXX9mHIFX5Hwr6Q0zRln8cFxYFGDKolTqavSZ9lsR
X/8mBbujYF770lETdBjeK1nsBZeXZXI5PxWEZJfrG9bZmz2gFCeTP0HU6pzE8b2vYYh2rtJp1n9Y
YU0JGdYtIOYk8EUjmeNv0Cy+oLRm1HLLIVqJu9c6ja8+rB85miK+Gm+f4wCoP0x9DNAXvX6kHrTn
Zuczn4t33uAKdeuF6M+2kd0Q9zYgV/iVE5+sLhs1r9eMIWjvRVp0SShP9sW1JSv1EHKqBn13Qw/g
tAUoJeAs5PKyfH8ALp29K1RKUn9nJTvWXErA8+7MD1BMqdaO77UtUyT33IrTp8fdYWTAUQ5ubm2E
geHOmehnMGT8a1JfqqGeJTHgjD8lNFP18HLxSh+Dm3ufvpFEEDQLErzLfCjwVWwl+0aA23sLqkOV
/3uh9wuCXij5FjPx6hbw0tSMa65wIcmzD6hHU8/rIBQHUEZdhE1f0OszptMB2MnFTq1sV67V5ru9
XXTXWJ20dpleP92yhGxBykN9P8asxKNGpnAKWPLPq8GvKdhhTOJOGgk4nzAu1dVMjMA2nAqLW3Zj
J0xzYX9F41SPa9Gy8qQgajFjQPdJUGeImPCuWmVaI/JqDM1PDwLw+ePYcK3Slkm8evDEaUeFjgYO
rcTZ6vc/XE+rKdvAYeGcp6g99H6kO4B7rJosabNpHGM93agko572t5VnYhYqDF1sOm57N2e2cyso
ZnEYv4Brf/MMbtw3VxHG1LHVSuf3MD29Fgox1ELQ7sJhGe8rdc75Ia6V23CXT/t9zgDtMCCcZM0X
FjW48acfs2+tR8u/t3vd8s3ZrruzzbCC/pU7/QNrB7nsXkJ0wYUtKA1ImQGKHXoGgW9UQfPka8+n
anSw9KZxSwbDXwwmL8ZWe3R37PzviY96nG3FV9/MnpYmsAKdESrQNaxl/jUB05LbJsrr47tXLEOL
yFny3exjX73EMRPuWsLEwy8RSPGvSLizCKVdLRdUrzlUByimJh+yIw0Lydp9Bv5yY9kanttSsupd
9CA0oI16W6eKqhJxEWiAtXEq9MBAukfVuNknZL7hhE4bKLOAeJY4Iy0VLTJ5GbKOf+WIzxwNk9yI
byfs9RyoFYgN7tHksxSWIFO0ph58X7vcDJtnU75zQkk62z47OOFwx5lQV8TLw6QnIW4s0DQ014Qu
wZg86UxsASBkw/d+hAldo7a6kTepgVbl+tPKtJZiH8y4H2FnQi3+yuGzVfuEWJvwSvOfNwZhwnU4
bQ3vroYvgTVseuWlulkJZ2GltdbRoFvDBaW6+eKKqnocmRIohywifJmU0WfLpsTn6QoKuL92U2Hz
CtNvcRhG2mQD9mRvDBgynZtR+BvHW4gFW4MenqeUFMvxU6uIcLf8ic6wywct1JJwQpu8hznrX2vR
Wi+m49xWU9ArJUmiBw5i73uD36qSPh5Bdrf77GkBTibtiPbAaRQwXHh+T+MtwibMTqNjdROSh7+r
UP2hUMeelePKU6bjtQaBDyE3ZT5N4A43W/lrdaEtvlDXjS+/txPXw/TtKarAcQ0U+Gx3PPuwsjXE
SK7k+7gi8N7/Wdh7QZtJmJuXYgrI/nChPp5+XGW2X7LT2jUOq6PZiD1FUI/RcAPqipc4YzaSHF0P
JgG5yYZBlNmUl830MSBZSx8aXFNyhey/Pe1JTv9rjuQLJHkqhFAruBAu7LwktRc5WX2eDxc80ycF
YMe+TvhD+o15Mb5g9sKzPwcqbZ6du1Vc3bWHGnY87tVSBTJGW8jclZP8jXH/RqsZGVm5dh2Lcp8S
z5SPYedyGOw43jznFSP+KrMz2bOGjzhwbRCogDQ4skK4s7Wmy9/mKy9P53gtBjptIsLppokxIOrm
hDh1Xtm6uS5ispETIjK7NZF278KVhp6U9cNFmzgB04W71/EyRJSHE/IRQy4cwbgKpsXd1FtqWDVT
88jokIWiLxCSjtxApbjmeXcGgHbrPmtt3Gi6fUj7Z/txj0WPpxOCbU1LTM2aNKeS49DcAM7hJiW8
8vg3JPGrvjqhSVqlmHFEtH9KX8Sol2Z0NgYMZOK8VBOyt0cScLB6EJGmO5bO88uav33EC/CODzkW
GWJmqZXE6VUIPPxDqS8VHB4ijCIqNyPqqWzKT6CnAjE2yXMMv1M4u57y10ZreJ/mFHg9MiGnqGHG
xawzw08FlkQVMY90htLELDZtqNOp7qD/mCyTFtG3xd2u9lJEpQE728r5Z1aK5XcFnWECAlfGsqEJ
T6ot2hnA0MGsi4/FOcrvQUY5DYgDQND8iML0+ntCvPB3pY3h2pnveKXJmsM5djKYn1OKUqqBB94t
SJVDtcnbF/qm9AtW2C5zVAgOeu+rgTKfxlH49eCYCQSEtVQLzKO9btxeE44AgvgUZMPkmiozNwue
Q5h+D3LsJnnsQNF6SJKOLrIiHTdKD0U1/AS7tM2bb2S1xZ5+ZJrj+++c+Z+mw/rPAh1e4T1LMm8o
m9FwEamDjRwdT/QcSu9P5vVJwh/G/ZdFVcwtH9AtScDDiISIGVG39MkUQ+jCh88ikewYdcRHiiBx
DS1pjyrEYve3HpR7fciagsED/PyD9zCWJ3/zwIPf7psgwRvoeIk2ch3v5Eo9Gdf2z6rzA23ygh04
SytCKB5KmFbtxn9ubEt2FnRc/cPmZKVKQa+c0jfumMLyYwSEK757TrL/yMMZ2UsMys/aXZ8JDNBf
99z0Q3pqpz29id0HLI/KHiiMlcfVCxFVxmXwBht83yxyBM6aCAOt1Ib7sdD/cSNNbFFKhZfqocUT
ST6z9uKgoSWMr4yu7hh8UUYF0erlZpeZNiTJ2sSyljs/vbjNKgt9pKFs2fQ+9WZhdLeXlri8lb3z
rAdWrtiVy0vA4XBr0BE+Gm7OLH9l/RLPF8OCRMPR/NfrPVDQDAvZTHmTrHD3WQ4GWKsPeg6ZkvtR
L1yE6uWW7rzdR/F/EolFaaKVEnurTX010jb4gQikCQAmnH7Wzju+mYFbjwKO0GE6ONp9ZbpiS1c3
fIg+r648o3O/7VIMNRzmxWjFwPqJjbbshF7q1RTVOzZIKvUhbV/0T4tE+bBom2RYBjqfMLvXj6Gm
gQDgzAuKaUEx5HBBgqX/1nXTL9XJxe6L03ich0RlT8idvf2Ak/dqU27yUQwtgCZHpLqFlnZo0oQE
xspiPhYm1ntEboO2410pvnGAeAoqWVMdgbGMZQXNVoTAbQqunbO6Sd1ffqn8D0yEukrr6K52cl6n
EsWyW9hfmbVSDd3h8Es+Ex6tT82W0mX3W9DRGEIkgYNgY2Qqt7E8ohSGZNPzlteGk5torIuXgkJd
HPcgQWrbXoaYWo/x/MziSKFAeDhqagbk/iW/j6cfSafYtiHE5AW41Tw/OVEhRJ07Z1nxkJO/LmmK
7yEtNmvKr+jG1usp9sgn+TXcWS40SabA5StWulRrACPnApHF7yQYKt444N/b6dqj50efBgrzuW/d
bWi6hqM71FiOXH8g9ADiaOYYUYzq8X3b3dU/oSnKLARhKzedK59Hn+RZfCSbzRxwzgRGYwWEFfnJ
VvNCxACCFkO0JKN5Nl3E6pTvkPzDHnk24cODUokW5RK9K9xu8+XFgwe1QHIvG7bYWYHLVuTEtY78
bK5tzcRNlVxLjphvArjwVVsfifqJkVY42wcILxNAByVVkgP8zNeJIvsuyaufabaI/lyKWj/Mh7k1
6uaOIdmyOyv4BypC83dJVgJbkLylBekO8pdZ9qg++5yVOCDV5SLRMRRMTtpqqZHwdx58AqJw6lr9
R6JD+vK+dJWrhi/UD1hg6Sqanhd2cF2QRwt2vtdhBVL6y1fYSEMIuJC8KF2Wx5DNlJJsYhVteR19
xXgSQhvJYdposDsub5tO98qUuldC9jmu2IIWRC+ZVai9M5EslP8q7PQ1fKpedxurJysDBY0gR+lc
alHIFAglNFayb3RncsBxxBfsODN1L5yWbmwBtf8eo+TImRh5XW/4Tixju+X2B+vt597HgYiZqz5b
lIJ8esgz2o5YUDcFKc/KhSihrYctNmkCVSUvC2x7ls+xGvAJ8MGBHrGC9mxFjl06Wz++E29mSHQE
mOioL/96/JCwKGnCG9wJ5n8IgQoha/CD2ucRaw560UcDiNb/upYp0DF1Gja6mvqJzjPX2Pcx16oP
/gsMyFkAmZvXCcZfM0YbytTagRaB4tETMex7ab1APh35lyFzDB+AXJgIvoxHyQQCaYLTdCkBp18C
z1cguqVHAVnXvqT2RaFwcESSt42tWsU+KicamP9Tdkd82y+J5C7NvSuXemcrBV5zWDm5bqMJERTv
SVOl+6Jx5ia0ApvfPdD+FLANYBwvpHigLV0RY+iXesFOiCsvzgbVTJTAM1TvRRo5ON1OzxSYBicf
TLUYVjGQbxglghLelcpV63gBeZAU3eHpsh3agc+RSxlhZD7zVDgaE/TNNRXw3SwmXzprBPAu26MA
veREleu1Kmh+xIIPz/Z4C2Cyk4GcYRfWLgF81TGbrzL89/m6NU/80XNzj+MA9JvJvBDBJ0VlC98b
enmus1jagAa5z+W7IH0U6azI2k2GX7NQYb/+gKi4/Nsjgz8NyRzKfq+MIwBQcmrG2/DpxNS/6bXP
CE06C+N9mcfCIavzbEwjz9hGxcYHQHfWJpx6rLlEy95Cl/N4BqdUt8HLz+qEN6X8u47kAo5EfDaO
WkVImVYhR92tAzZxJOVNM4xR09pqZCWPdfrsn1Vat7Na9MzRUTmue1ovTQ0V9HVlBD9k/KYZ+hHa
00h1l9a2FDObSgylAGtrUlYRzH8gLexs8wzAxNlff1IF0/yyv+I7KscpKMRNItJ3ffZ/WlptAsYr
nVE0RRQwxMtjGowCuHatThrp8b8vnMuvlkMYXYZ41kv2Sd3VKIdMT0EDZyG13OB7QniYpaFxpBXy
jCCiKx5P5vOc0mfr2DL0rNKS3rlkrg7wJehZGwHxQ4J2IZ/dt+DECoqkGSRLCj8nnNsBYxbneJN7
uYNoNXpq1+yoJpdHnlniO6M5g3Hj43/1hGBlKnbtWKGs5Z57LPTEVW5B614FGhlNU3g4Oqa9wWyq
TRLdNijwT4y5ouMDn3Td2hIZtdcKLMl+Rxen3Fz1eGs27kbLOXOeF4qF0TXM8rFcvpNrvi5KVEBG
xwqDwaixv7f7d2gPh/dHhyfDMFFPEwaYZ7YudRrOjm/gULvnBozMIs8CKdZyoyh3OaP3QEsWqN1B
z75P0SZg7ooJeksRKa0HY7t3RHkaQ4skhS9TXIHAYvxUPG3Yn9iZoGVhxWYHqKANnSzpG8gWXqo/
RdngwZnfTtFl0qw1WgnuTFSbhaI67uv8zHHijqAhTdF1BmE1kU8YHNFJYwF6OXhDaE6lMLLtGF9s
m7r5W0bky8hjeZi8MboJtYRofWS/NS1J1spY1nTKe7SNm8XgMrGTxTFyA8KlFuDivsrBU4sTkWk0
alRcPsMJGguTnd5ZdGdY4HataQoggWORjDzEST7rmgwOZOgpmYoDlEDKC0qNLlXaEsIhN9Qy4K/C
0QbKHCTdyXcErvvfhgvNG2QrAcnOx9BAbYVdPeQHZKLNGL1eDdn92Sno+cSn8CAzsqzYRnD6qSK4
wwr0XglS5LCZdE7qIXVfD3EztRlzB60l2p7a/zYb7qm73A1kDvSvu3MFLTxv7AWglW4iIM/7NnB6
FVihpQ5eGLToxhAE2jAvE/0FLEPmyfM7izCqk4DwteiiVwIOc+7fZpIEBkUZJsY9fn6A4OSRKYA0
BhliSSjVxABKNybl5B9RHew+S81EWbzocgZzhu1xcok/vXprzbwsHFXZAD8JYD11Kz8FxQegpywH
PYpoleWDBQlPnYHvGb3yFT91XnFc9WQ8pvUk7e7uKVc/PdEoJe/9eeY9gfmFht1nlk58QSeosYOT
yb7U5FiH+N/d30NDHTmQizFEtMI7JxWgVB/LgHuV/SvGvrV6zYr5YXCpaEy0rfVd6GaI1/InsVNi
oRRu3Sp9633TBqUoQJ1q8ZE3YZV0sa/K6DvxVaucKFJxQQPb735qF6DPLKXieUx3H1ImBr8x1sVV
GBbsE09RYtSh8o2a6Z5LHGFXHq0WnUZ5zA0EflxMEaxK0t46Soo/yfMddmaPDDUNrVThLIGaC/a8
qFBP5k0DtwsmRgHbSJRSvNsl+AcTbdWl63Z5+u3X29N+lTa7jGa3EyvtvyB/3gZDzb+y+jM+HrkH
E9508YK/KL3o5fsUxmVmUo+NBB5oksJlTUxGUZakVSXuvwHkiqmnSEQ7v3GRwIfKW8aHnEg0Obj2
2VIhblu7BVp3MV08x9Wu77KgD+tA+hzKfgazims6OIWqYNDzdEzGZWyuIUKCQdp6Zf0HwZLCHY0m
BllTOlgybrcbkHaMTbMpTw4RFboCs4ekEip5TnvrCesFoCrD97/n18U61L3QPxheQLw4qrl23k+q
cz0OtrVuoO3De5nCoxnvTgTJrAgBYpKQEXkIAF+E670z7qRB1l52e9BkVl+mUeRv4vFLHjfYCUta
MxtRKzyCdUylKFwNzLcsuqX2OHfNNgjr/YPKpRPzSzpHG5entNkLdnL26SE9TziuzEDwXBtA14JE
5ilowtJT+tm4+a/huurzIZY60sO62NQjhT+mmUsLoPpd7+2K1BL6RPeVnnwpX/98cICTQG6mYqN4
D7zo0njUnz/vZrKRvtNzOy9H8T5CCqy3QcyDE7KxScr2GLb+pl1ZjXW2oIbn5dadlz2JKzydBRYq
oGT7IlifcWJ/rWBx3G5sfahN+DlMBM1wMaAbGtv2+RoKVp+s2+PWEEOqDyChixjyNmGA9DwEDS43
Zyf42wlisn4ifPc53nloWjVmov0P/qvzCX9U7pFjPGDUAYIPOrDzbmWXLkSD9yilsx7hynZlXkX0
StkAJ5mubnpx8YMvbJSk5lSy/o1DFwrF8FNzGfU2HqllMXP66Tvvm9eKM3d20q4XdtRiI+cO9xsp
WRhiZoIZgSt5/0XeIJcFbFskFUEj+5MbB2ei6NRCxkLUyAb8nIssWnGMvGU8ZIUyB911ikE7mEe0
8uA0NS942CathckkgMZndVGzippl/ydRcTlXsCN5cdi8WeSCfK5CucGJjvEPGn3xqDuzRgoCyU0t
M1nzuDdQ6OmV0XytaOBHDhv98KZcI/BQvtDbuAK++se6PFlVQKfaUciZTswcPrCQVCDB+z17zFTZ
Zn2SrhY3xlSPvHIHU3sHPO/EdOQ9Pruqk5lDbLjchXc7uTKPyg35vew4lvWMVzfxM3adOyQ9F9Sa
MfopVRHBzp0f0Slbc8RWetRU52a3Omnas0g79cJcxi7ja+ditkOKdAOQWMZQ2k3DMjEeQVWfIeYR
zeylJaaz2MzfGgA1d7dRxk59M+vocWJnwnNYGPt1MWcB5czlMUBBlrYdVqTGCMQTwPN5i8lwa0Ci
Uduiva/GGHDOVUubBAS8J2lbHFZapZnIdTKNBGUWFu/MKgElDnjYc2+xxhwqDMPHyidrWO6DIKUH
QUwsQqRtTsfLbYkR+TrcPZiiBE1ebNjfkX0422nXCr9GBf1ZE5IvufyifQ6TPwPV7EC2yZxJaY7t
wBMEwPUHMQsGYZDZyl+DCKG48shiS2NfKrbYXZqo9LyLCpMTBM4f2RbbULZIhJ69ZC+9vBTM5B5d
4hiwLKJSsG3YB8noeGBL9vaoG19vAkploiqQhFE0N/Tm+H7X0Y+eVhrJOtUyNfC4nDL6hFQ8xyXu
CYDv1XBqhMsOpHWWmN0mBW/Rney6FCzJAVR+DY3vJ3gRWQQdhELelUTR4hmWrnAJnDd4LjZ9ZxZQ
L65BXRKDslMV7rmmD6fzULgr7bOyQPJvCE7NA0Qvraq4lc14amGNKm6sl6Y2Jd10yMAzM83zLNQI
G7PtRNM/3ARdZPtELjD94n/EfVJx1Am65gepOA6IkEjH3zlnTrAHqea0+WFsF1xWuZzfqM/YBerB
4SH/cdaKhZI1J1+YmSlxuXiyiD+9aCj02n/Tv7lSfo8yre+iyFYi8WP8cLBl21/vaCt/F4dKNOeF
az3WKNlKqUgXuNRvLJZoxZi0iz+OEhfGelwvBcQRuRgKRMJKT//dEoCPr+uzg9+n6sUGcJv5L5DQ
JUyUekCYmp8l9g9+IdAgLQ/iV4pPwBInfEaZRhSFymflCTB98xZRsY3rSmWdRYRqJVaGn4EnqWit
DjLde0Y4imvBVVlQRoo4e0tKSLjwmG0/MvOuWJ2Xu4TKKlKfqXGHQxiaQGO8YLVJTYC73Mj/Wbx+
I7h5MSDsKLyakK4a5l8xIFPC0bvUqG4J+lM6UA3hiZyAYnp9Qzw9v/Pu4FQn2mH4W36246Srp7rQ
oS5LbfRNkfv+R6z8peuaqNdpGMObNzD83DzIDIk5m3CuO0MgwoCqZU8LmuDCRy84VSgCl/adLA2Z
R5LSt00wj3G+XwEnsDOwas1gSYZ5GjiDQpumA/5O/yDsb3Wtjc9jlGKSk5DTYJMrR4hARhCdwMEz
gT/WIBgIgf2g4DxV65e0awYCjd8PY6/MHh9Wd+/WGSOW1A/mfbtbtVEJoxghzijeMV7G78UXLceU
VMMRFL4osw4VCxsrkrslMWOvrIDjw/HLcXLioxYSS/lHn0ylQstDeuVqKtj8Pnl7avFRo7h5r7QE
vTytSRoG3YQ0kjkGO8wQMUMeFjDj0gKhaPtLpKVy2EYILdtdYEqfovTa6BuFUIUdWeW3IkG5/zZf
EvGzWde0vteFY0G3H+1wV/YizoPtd5b8ZRCwfGSOJzJl9QuK8+Y93ihJxicE6Zd3IVb+T2Hx02mZ
HvHd2pV3LQl5kstXC/cVmEq2NtwC/NEVfkxepGO4nUOZL8vmUdbj1R/X7byd58AFmOlRToBHh2K7
M0p2Ouu/CBpWqWbjF4cKK6dR4IVsixmG1LAmWPrx3GZTyS3u56XduQzqILtxGzUOHOBKicftBjoV
HohWklK7QNGb4de/6kAXT46VjQWctMH+nNwjuoOTYzrrm3oIWWOqR2tvLvP0BbqjI3ezjrk3mw6y
otBqvIxCTFtVCfQpDJ+d9NtsJRsMhfz7ivhC3Ht8EBv+CxzlIRxWxy/6EqVejNxt9rJe3WtfdMTA
qX19RzPcRX0G3Qk09bvgrcRcJWLfdJdL5SfV1euOrdZhyJw/Zpv5jqu4o3Vb+kePV6y1QHU2sY1p
ODLRkQkc/zsE6GKB58E0UvAllwsgD6axVj3J102sCqElUEhPIqJUJMtE5d93RwamcT81NPdsdJz4
kj9Szm1jVZUg5ZISyHrUm/rOiR6HEtdTVa1mSxJArwpwws3njneRK3K3DGOcpiej91VUzmOZtl03
9Sm1ALBEmVpz5Bt6nEcn0oSZb5ab0yqGdw9g1qxP+0WEiid2B8FyOeig96V7L5afALKsAaBPOK0Y
soDGihmsG9OIaN8GqI666v1tSInUqunWfumnk7YkG8Jcd9AT0myRvmluWNwzqwKf995s1/PUrtNE
RYN80GFRW1IQFuhveAJ+IzyEVikbSYRSl7dRN2xk0oQndABYgUgB18+K2skGswrexivLTB9XAngZ
4Oj1x2sJWOUTkN0YnHk+xWpjjmqueEBZMNZH8TioVlxr7M5W4OMWZBWx+D0tegG/xLmFopEx0tBL
hum3WfjEiBNnePWTxXfFUHzET+W93Aaw5ISRPvcGV9R7ZQdkzli00bnudmufyg4XaxHhi7fnXvZM
M6wTcSFS6PWs6bAzkUJIMTJmkAdbWPmp9zSPc7jylRcqUKLLUJgQG+yYtKAQqPiMlF/ai38+HMpY
cM9Y5CUCS+N9mvbAZIW6ZC8bbZaUwBxutpg6jDZ7+FxtRMwu0jXKMgilhdsZcRKv5kBai83oTxk2
z7o3Aq5xjrMIL2iPExgaa1WdvZqceUKM/1hJ89ZVpC3wZS0aOuKd31cUwuwVVmdonwVuURH+KVDs
X0uU2v+V6ZLIxHtLffvvbqH9vMUJmZdNkAD+IaTt2yBLIE5lzX83pBDQ/U+BjNpRz2L3cw5cRdld
Hr8oBWxGY2OQPDRr1PfDLyKgHbGPvWCCOEYBzEX3KlXg0hq2neRawfxlS9JP8WtPcdQOtq5oIq7p
0SffhHdHsZJSDYZ4wNxduReLChHwry3HAiqX28Rdi3HXujEc7+BDJ/8vlnMRsywyi/n3P17kIMJC
cf19IOQMn30YfsoDCSfJAuGdp+/3laQ/MIPjOxa+lkmdcHnLi8uHzGucs/JLQB2zV5X15t7B38no
/zCI6ZeLtMN6qb98YDu9C2jDadOn7F+hQKXn76G81Sm9nCaKDlxiNLrGRJVSHRdMdt/vX7N3AAuv
Usw0xAgjNQjAIqGPnLT+3MzlUAmI7yhZqBDy7O/EPjhTzrSPL4wpHz7+DqGr0a9ih29S3gJc6U73
L9xK4QpIdLCJnuNXPuPcBuRkmjM3+KLZzMKzNsKTPTs2HA6EfN3IIKTGrQoqseFQ7Z5bB2+itMhN
YnaRY1pnRJ0j8YCbtAG4LwcwDVVqV20Kc3Eb7vgf+lb3BDIUjERBHagtvHSWdI9hsNNl/Alz37q9
FdOzxpq8sgwGVsSNhv9bRGi2E+TdRPFoDIkGm2AH3YuyBgE9gMIpPWYhInBURYfU5ReqzRt3kR5X
e+wabdsonOm2zZbpK4jRvwM1gP3VxPVOCu9HO24v7rnsbr4OOlHj7wbBxtjMEOqIDiBYOJz0cNXe
ew/NA3bmjqAvbB6w14T/PgGTTUQw48PrP/tmqr+pcKc5SBDJJOZJxAev2VBiDw/YG+hoL54OI0qr
y9fHQyCBIZx3NpMUAKH3Gl1l0Q19oDYn6uro1uZdza9CaayKf5YiWPrRhkmI/G71k+KlXevTeJDx
pVkFYmYgdNCwzbadkoH8/DXhkGCRRCVV/WYkIca+Q/yu7VzbEsUnL3CeusuP7MrmxCijbQky/8ik
nGVel+d9gHfHbFL31GswwuJWmIP7llJD7akRSvP3/SN2fjTLOmzXnq/f1QGyJb1JTAs7kpXiTUQz
vNSuS33vCSn2FsPdw5/XeDMusoVv/kcn07mx/NP9Mjx6jGTb0Vld9cglS807PApz4+iNIGocFmWn
9eQpUYOiaVNgZ62Sx2D1hH3f1MniE10SdxEYzkpQbQg2USGB3tWKfiMHfkL7HtDodtub8QVlN1Ca
ax2Ym3vfoxbiRNMtj3TVvXPZLIAXRGuZgjTFACm9UcXOuw15kucKcAlab9m8S9Mlwck7dHPwXG/6
SqvfpoYvWNEOYpU2ItVAQQO4lpSPAZhqmwDjNymQjLEr78x/iUbovSR5ezPcS22q1v5lu6GImRiy
GU3at7nibv3ct/g4fzpjhjaMwWhj7MrVDBKh30/Pg0Ykd/z5dGJqzReYYXgGt65L7WROcNoekRWp
aV9MfcC5vlQLj2+iYIRVbvlJmrkfMnLFU6gICozGp4ZhQ5QeAvOtm5ZSJZHvHK0ELI8gR1l51IQa
LJ16q7Zj6Tx0sBsQdVre6XIbE+4ErhVqI2PMtl+qb6i8PfL41Sxjjl4kqUBdfJqAF/8MMMerwoZA
jMi5OK6yVW7Qd941ajDxx+E6ACnTTj4Lxo9MwnLaFBzbJdpjq7uOGC59oNIYmBCxxCrwUUfB2yln
E8Fs6JTBtGx+PrR+FqWffrZ7b18HfgfYSEUmFsTU1MbslB73TytnNPyZ4RoKVMB9agjSEEGSXp8d
cjNs9xnYgarUHM421Hb1V5sNEXnvP3RRKRW6CY2ZDUr0YQJeDQGzeGc6cHoV+Dd+8OXZVZ2oPgDn
ddOF2PGxgXKqAYR/CS2xR435gSF8N+O4tMMV5D4jsDwmoJOUJtVqxiY+C4ZUttx5OYDqnSEscZ72
SeTjI+Tt+Wzvy4uiVD5odYvuE7DZ+i0A9v1KFIZ8m+hIhxu1mF5F50lO/F37tX7bS/UAyXm3ZdwT
kfnlOSMmYUvS+sNDOJypCZtBcPMPdkdGP1qBxExdM4kgAodqIerM/20AFdvdMirDUQHaf2/JUCS7
LAi2pE2fGnHkJDnLVh2P29hnPWaeiiuwUqDu75WaH00mDUBoo8DmOgxZqF+AHTLyn0kRGe8/7Hax
AKoYdGwaMkNsZjsYCmlbP4QyLuMYGgRO7N2pfEYJp7Ted8ooJfvq/WHwpU33+x9htJBy9QhQJgKA
wLCcjywciQapTFisyYZT9XfbANEvfqCnW+uT30tZt58JHFJc7z4dEBZjXG13FCRBLbuW3LfmoldW
v9vP1qcuCgcxejKPo7fqk3DaCpwiuWcnvad476nFgA3EuOr6x0zud15KSDi9GdaQQK8SCnOFa1Vh
q+m0ThtJyEe8UTqiGkFswaqm//rEUHFri+ZbTv8wyId695fXioYEH4qbomupzbMkHhTnJ1oR2eIw
oBiwkcxPgwBdISs3TC9gn6X4r4C0FaLdDdUC2Vx3zSlGhrZZ2MrFg53aDzfiO4gybExlB5VItxKa
B8fb1p77BboxMM/K1rxVOvolB6AGxp76lC+RUo/6SsnCvebsHcKHQ0MWEtUOymg/dTCwtCKyPYb+
1Ts2Nlklm+hZ3odnlUXeQZ0rxj0urVBbzX8maYOW5XRbyrc0Sm8JudYuydHsQDCRlWVv7JiDI/0n
/5LaSmnRBgz1cHnUfbuVn2oZhKwj+iEgD5+Jg7U67K+wXEWvL3toeTZc+wO55HgArpQikocz7CgF
9KXs5UI/PGeXK2xS2Kv5//3lyYxfQ6U+jkyxqHWyAjwtSQ9Xz1/3Cfra41Tf5nUSDsCs52B465Xd
cAhcKXTivgrfnp5Y2LJYPdoLm+gxNUyUiNf8g8LC5d3NJgTtuwKk8Oervc9t2nJxwddZsBdyrFOq
3mGo1bDxEsqfhqH0taDS+ggJHujU0YywCW1qk2efCRFtk65pZH1iDErpKINMXVFSAit+4uIQJ4uG
n4CTSTdZ04xOEclUShIfdMUBtuxPhAr5mRMqhrnEAydoEnzfIVWvoKVmexF7CzXoQkBKjpbwajyM
0CrP+QenrPR4k6oJqzPZ6LC4KnSY4yPZ31omT+hXV2QfG6HtesrOZJ0u062hfZVji781bMW4ljOb
cnb9n41BwAFObg/FSQdl5/ydy3Ipsnb5xnqcjfSLBRSFeSS12rRb+NG1JZNf5uHxqPOF7pIxBRwM
ChqIQ8mVpKTgbgRh6+2v4OVriEAqe5h+rD0FfoOYcxmlusg+tGV/yXaJRPtdmucHcAl4BmTEpfZB
XiTzWflR9rqMFquHgwFfV4r+1o3Mc/75wcpu2l+p1Sd1IHsqRjjhWRiz8ISu1BscS5O8WLnp9YBD
emngu7XlL9yPKh1xjSouGugQihuQASmJUwcphh9ZUjERt7HuhF/85CPaL5HqbR0KUG94iqSIE2PL
QpJrymkzwrSyj89wReEc1aZ9daydBOyKGgH2dIHejDPP2qO9QyxbQusHNtdIXntvPCBKGRAHpilj
zMNxRURqKN3fyAvUSJD9Fk7qlehByWXZO0/zqHSaeR2+YlQ0ng7D9IDfGlEAvsKHzIAE9LVlQgsN
0PiY7pQ4TurcltJbWYsQ7TGU6HFARuggm7wYVrHq90cqnvawii767pc9gB6zSfHCqZ6vwDjnW9AF
b498g6pRPAJR2itXDsPsSu5Txhki3KjqqTCKrouSp2BlQILxzPK5rrchrOCnUZPQKBJoFBbrDEfy
1v7oGOrDqU3qjwKW/e3j81w0b6ffE4CL0ic1FxKNwNA3lddVYMWSxKD0+o7Nsf5K77YkCeEeOHQc
RrfIbgTfc0hgt4bKgfmWHkXNC1wQMjBLoqa3yugTJlCOD5r1kyH/c6HuYGaHt1k9ZfqMTK06CuYD
OIru1Ds/idZAoV2FoMXr/7TZ6NvPz0GJXVZxSv+EwfWVLlIyzFlprLX8mhfvJlT9b+ws9gSZYqLw
W35xeKYtRPg/btik2QD/W9dLCjsLfMWa8bRJMCW2OYUjL602OGSxxZCdkdJY6qFFuaZrpd6YtW0X
/hqqbJ/5n9QC0ogMGRdt0Tc0SyHZ79YRWVDycF9uWyQWDYTCTy7JjI1IB82tOQoFZCW7AUpgoPlY
+9yGmu6cbe+sacx1RtRp/1Hpc+z3fLnuzz+omdW1mXnUPoO5GmPNKWPEwAOzwG8HkEMp+m/pk93g
LWlUdy+XAA1MkOZB31E7KbT5ppw8beWWLJSzm+lrgi9cun35ZxN2gzTzTFODxk+6mXkYq7wED8hX
g+CF0ryty3Hewb0J1HEYa7JRixJ7g3wYr9E63nWKq8ck7C3/xXyZy45hb98dk9YJJ3r7973PMpmH
UbTsafgNnoQwjQg0SKzJyVeVkKI21kh5/psNYrs8P/fS9in0qTM4Dp2xWk1x8gOZ8zVpDkYAw3BK
bTd9Uf2XLEQObqFFGw/xA0TPhFkYvCJ/oUudY0PWH1EYUAZ77B0Jlo5UtP+Xk2ifyQp1VGkYid6l
fiPBdLVfpyUbptcjAf5+SidqPh+MZH1nMtaGPeh007a7w/q/0xz1s+EFipiQBL0yFdYPFHnk0EPn
GQnNdpwTJ7ErVooQw/PAgNtXJxecV7vXDzf4mPY3JDx95RZGHBmo03gWF/N3KFaMqqsYF//JjUiy
d18j0C2o8Sknb2C/E2A9WZMsjec2bMjffz00UMRegcbt4WeHgR01TgYsa625XIjM3fhc7wsZ5/Mc
pdPkPAfkdrsqVy0+C26xj1SqPjejYNLLCSlLbsFmluKT030W5p4cbQxojLqYyjCn6fAjvhUZ27Zf
8sNH+VAMcE8ZjtCPK8I0TT2DiPexXdktNdlSr8/DXXLjCh2qy2aPS2hQOpHCSRaE7IgVrFrLbI64
HQjrCB8kAYTPuf6L2cFTCtTQijm+G8R1zbGPYSqpuYpt8VEml8XyepZN56guw56EabTJJY3B6DJ7
3cLGzntYcWMyHjjSiYU8QlpRBZDfYthLf2HN/fs2xH52ogQo3Q4579OSSFhRvsD8Ww/3pBdo9+qu
OiCukSbmn0tIIdxBfnPge1bkZi8Rzk/5z6BfhCDO9gDHqVXqVzkRiNP48sWo1b2yR/gSswwrw1jr
Vhv0v92DIzDuAdACe1boRz2NJISJP18oaABieLrujGU2DAgdy0jg+DhtVNl2Y4EdS9MAqxXFJtAh
k+ecoge/kig+w046Xnhl2G/hXy/w0s73mQ8wZ7+akN98VSo9yLIwakuhkzlFgMt/v6nM9Cua21r3
Jb216bgtFlVRwy7EEhono5Bt1c71pX00QmfaV9FdXDh7iFwV28W75Iq5mVmuycRplR3if3Hty9U4
cd7zSHyNIL61mT59REferMnubnMnJaQapXdxiIaTYZJ+xv+F0c1wKpcwWfqZAY+av7QukKnkK7dr
JxqnXLIxsju3QDeqite06dU48viQQ86Pl/6rH1dzCwWhXwvxjzt86mracoEuG4tK0VHLZPk+wfj+
2Gvk9pn6Rbe76psGqttUME47vUK5ImUvJhFZKk3P4+814TgVkUIsjb2z9Y0aNsYk2r6LoQILmmIn
AUMM3/GfeD6KP6IQYB7uuUg1NbiVJvAwC1fKeFARXH815JXVg8hwLdYkDSSx15p+uvbWFtSCEeJz
TNzZjGRACl2zqTViU0NE6EG3y57tPChdXPr2Evn65TCqssTZlimcPTEZYOxVv70XJJfWhkp59Agj
EV0s/LcMiRDpAQbQhvpRFEJBo8yrjf0WctMiZt2n/CoaUoOAvKScoGS05rHJJp5SzvD6U7xIyxJz
aCapYRFlbISQxZnqf69reBomIOq21ozxzarDwzTBkcRrTe5BuIPcmfgQO2+veAJVcVk4qM/0DVeD
bj92e1/p1bf+d5VaUWW9ss3yeLAdbo34HkGON38c6bDulAMaWwvmP9IiAamzgb9z8Dm5wwlJV3lh
tGhsyLfkDSJg5zK28qSvLyMkgaFjDIF7qik51vVmyWxNh7BbzzmXlVgrt6fktpNxzk0nu9604Mvt
yXvWluRIml42baJGnQI+9byj5M/zcwtJzyUXBiUDGznsInhV0ZbqsIc4bV+/yCj2tqYGsUMMpSw2
ef47nYTwThlfVCtk4oSYmhYFuGXAZJuzw0w/dViLmqlIOUJJtyreJ5nG8gZnvc47A8oDQhjpZlSw
Vyqs+meM89qOCym4+zCQPXM5mNSi44e8w736R+pPvLb7EYu8Gz2oATCRVWEryRCIB+8MtgZglKUE
eP1O8uBB4EfwWTC29Y0aAnGDz6l7nC2DNWwsLJEEQEb3SVKp0dmX2vIdYGJdcUKz0w4KjXqLErGR
e/s6f8wO1IkjCtvc+Wgj1vRBO1Hqy+rHdbim4tBlg6+Qi7UvYYRwDOEKnHuyF8lgRvnXVxt+Tc/r
Qf13mirLJzkmphu04Uyws73iJm8oEhW9kBRWhe0dBfO0W6gF2R4mt1X64ViQuhL0j4LB0C5Ld1oO
/Nk0H38aEVKR+IBaPeNTNKKuw1ABm8SMi7IV6j78KQrdBmvIi5QnyPOC1J9Qd8wKGNvBoWrwyDjg
fW8+eWQsJ3qCGnpe7Z3QXYJtbZ3Yp1pNiWxZtx/xuW0eb/fwRT/blZnfiGdoWEL9bCpszBH7qkA4
usPFHZc8D/2o4yriHdTezyAf0szcpc2SfunNqwHbMp3XYH2AQm8JKh4zkyvCj4nmwosR1DC5JMJx
ZWhSj9trOC2jw6K9uzUl5HVKbEn4kq0+izlzn3RYdd/2yc/syuCCBOGN2LkbQjgsqlPu37NQ6fHl
SEhkyRtrfTUBV5HO+GeqxSAg366iXmHbtbIiQhvg461m6G5QTK0WDiWLiL7X49ZhrxtoVFtBbLvv
SSiq1CdDE1Hf6R0ONVd+wndyD+83BbEZ7x0fDCjaNCOxW+RO1togXU7BfgVeYuq9tJb4IIcgUqca
p6yBc/x0OQhtTYk12OPzxkW6xIP4Vfh7+Z58kyTyIa4gtIS/ko9eEtQhzuPj0Lpvig1hLeRGv28E
/SdUp8EhFqxeU+hQO1HaikQnO07JeyyOM1p6kkftHNEii6j3itFho5n7dx+h4i+K6i8r1ugjc0GV
fUJuqCIx2C563BPMPl0m4F+cQhDlxN1W//Z5RY5O2lc0vS6Ce7rJ4uYp8Sgpm5aHcO4ZNv4+U86o
qgyzYmPuenFVRSg6M20sT7bjE7TJfXtoxLC8xy9+Iv/SXqLA1eYGGci9FKvt0c6lf1IfsQT+KQFC
G4COUA8BXZ1HRr5wTn45H6zXjkQ2nPtfKLzqHCl2GLLmv4vP0ziYHpYFCf8VjV4PaUHgMV6Tl8La
tvVBRzFaMX1+OI7jrDQYRI2lvJoy4XqS5EYKJ9t6AbxCC5UICU4TmyRBPW1qPUIescRl2BReirrK
TGz3aZJD2ZQV2O/eaDKpEqfxSmz1B0QNMNLHzCTgPjBiaK6rLGqBYMoJnxQSZRPUzKE8FxNb7LVs
NUFYaFGaVsjRxpamKklq4c4Nh2RIIcQcrwZ/dQaFwLVIBt6wCNiBcIhKLL/VvVvCdiwXcSGfmI23
HD4HJ7W5v1ZOcGmrOzLVedQ8wSSnz3f7cyhi002TWMBlVEyCw7vIJ6urzGqSucZ2dH34Jgd7NlgN
J5QGxeCuiWdw6Dk3gI5jnqtsp4GjgHwauC4DPfWZY0ApieZp0L+n2mXUx9Bq7Pj7GyWXqYhyeTpl
uBMi2Prhg7VGnmPco5RY0mSHOhV0jTmQxruu/DzJ/9OdZObOkECLEE48K7MhbZQDJkhQvLCIqPHL
jBtZY67MuNWlYwKgwQaIT+g3uz/Lh48v2yVEfPJ+34lR2NE0CBBg00RrCKPmVC5jjC/wKOL/OUus
iVHXKawOWOxBwZ06v2rSyxwJ42fhXqWV6Lwd2xT4XEOENrZez3XN0kelyoHLWaVoFf+wqtNUifMy
F1wY2vRCQOKN4fwwk+Iao1qhc8WBNVZDeJnbSUNN697fCeLIO5qJXzo8tUqBUlxDX0JY5FgXhtOI
wtKHxBLXVOVTpygNujDzSBao+dsF8PIE9kem/HcUybVXU5k/yKEgV83B2628EOfHdUnexI0vDYmo
ajdazvVaF0SFODCEWTuvhRkySKG/I/CwXoO0hlLJraKCuayX8pOE+2NQqRS2fcj1CmjWpAQNvvCC
OCbp4HIMNor7MAZI58cjGx9q50B63WD+Yw1ta6winRgL/4oSq1xVHltgmPCQ4Kxm+KVv7+0NWTa5
E0tZy+WKx7WY3oYG0VDaWe/aX/Em464IKjwBh6bCmbxrdeqBydVeQPSO8Xep13oAH+GCw8atj5Ti
+F6FC8QkfvOUU7T+5wg0jVuNVS4bYIaY6j8TW6qSSxrh24lPWYw2sjb0ouWw0B0mn7nTzkleib6c
Ohu5V95j68bH/xOExcsAKhPR/5bqcEV9jad7bQ7/v38vYNvdVic4LYcog8GwyrFgL7XLeQNcQu6O
vpoCzCrRKSHeCUVk849DMTfnUvr408fLdxptmxrvGx2lvc/VqFFKFB4yicexLM74wK5+oy/s1xki
jn0BOP4l6GpFgozkHzxPRnjmPftU97GhGA/WAGfvcsTR6C0ICjpAAEyadmtO3ITb5cSxQ1T1kV1A
JIcUWS3244F84+Mks/qWxekvrI5QyNWSeJt6ZmZmmHNZ8Yp1D8Dj3J1zphG5yVsalfRQQ3TTXaYv
x0CWrhAWe4MG+PDGHv6hDnWgEcm27ouS7AgVcDV3aj/bZCVhtulaoJ0TUC4/DZslQa+oftqK3weI
fHr45nr49uh4qwb5hlknvNqxm6Y7293FdZpN/x/kktdQnyvYkZ9C/SQJsKl1OFZu+IlTgnQO7F0l
SyyRqmrqR4EECrWozxHIbnH63vVYp2HQyigE5qhS4kvuBnW6Edy19EQ2RHsDkOmIuRAdgHWyra2A
zcpBCN+s0y8ynwZmWnvA+G5dWpfcLh5WzXmhOwFD43qeNHXoT2D/Xz4GI9mZ4+2pBuG1emik/ydq
qsdbIqOuBY8TZqNpeZmUlEZJFTmgNeg5HzdzIOaxnZ6ygw8EVxUd43REZfxpYSJd3EmwNHhHKSG/
4UZAKn4WV3gquq22M35edmuUPqODa+f1Z1czNpn+cot6vRSNXZjU72d+1vYpbqzYFrCtDdeXdJbk
tkz/J6hyrQ65J079l1mycfQkUxaIoxyxZxH1plXesmHysI4XbSpcdtjpweSHA6Ns0lycqUi2i76p
qs920evawgxaEKduntmgSAzbTrK9ANDKVuediglLaJdACsRm+stwTuqmPUU1j8sU+uasVAxa9TfP
cvHIRwTfPUD8fuSmTq89TQwoXGbN2sG6MCqt5IfuMwcBB5gwBxEtsX0kcE86+Pmsjt6rwkTqvrTK
paRsDnFWWCo4QeIkeyWsNgaEAZLdb6B+ogv7VIGKHBnITvN296iV0xPWWKlGgqjliChlXteEwuEn
tE8k1KGuVzPfbvwVXOHsIODAztlL2YFYoxaKXmQVFBFTbGEDhnVEtACh/35NqmWWjSU3/iVjqgx2
Ted3mlhca43uu3PrKbqPteRW01XjCijIDIxiC62MV4oJjQ3OWcLaACwjE20xHj7hugaosa+kM9gP
EiHPyEDYiLUhccl/efLtnVvKfL2Y7oP+6NggWs+rmzOAzCs7nwlG6SfjVi8qSPUrIT/7T/Sho0nS
iLhF0wsmjhCrxTyiwvijb7bYyWkZD+hgjuxz2drC4yKduvKzGeEbQEWw8NOx1sKTJj0jG1yhfY3S
cJgYeZT/PypXqLAOxUSho6x+PKfh3eUc0oB19qBxH0Mk/pAzWX5dSH61cJDvO6n4a5kVW6bdvLMY
ZppZuwvcFZmGDCyX6Bd1xLV7IXJ6VmqHVZoV4m4dedXjQmcJOQUBUIh/klH0Q8rnvrUyK9vkLijS
CqGjn1uF4R/VBvYd33GuBvo4vggljJBTk4tr48LLbdx36Cztdu9rnjUWA2jwSBcwcMa8NjKu1oY+
G7nq8D5Ek4frMXbbCGZwa8DnkuM+O3ur3SbdrrHwkwrqrtO9+H6HTp7cUIExUCRI4ULDiyD8GrAb
20ubDJZQbx5ZXIcP9wedwwrP8RHpIdX4IOerTjyMtU0uUT2odZNe+1EfeqRx46AqYySDqWB27YNh
pVVDAtPznZm45aDPVX3KVp4pTtsh7V5skhkZ8bSmQcdlerYSGnu589g88Q8e7F5nwYupj9nweDxA
KdTigMssPXyHiNKqn4Z/HGdabpoVyphce2CeSBIO7dW2/cbX40O8EBB3S45uBFyDxWRnSkorMANd
A3nsrEpqgZGNLY7+soCnarYkfBmemIRLQq5MLcsZna8VqNxILmGBUeQJCOMo3bT1bXrFFZcO8/SD
ZMnSw7xSZnadtrsDWBEFRhLuQp1+EkPMHq1Q9JqYXg0adwU7Y9jYtBmKReLYbgbApUDz74TBIbk9
l/+Zy+Dwk0bp1HToilJnaSufBrTtEVInuMm+DKqGRIBGdyJquXI8g4otUWaqMZ88VfH7n+W4m+vb
wfImgPbszozY7x6M+fssLanz5xLZqlOHsXG7ILflRwSb3r8M1U72vhJvqhm+b0VPpRjwgbVu2wGd
3JXe2bcNRNzje8HDnuK9pBmfL40FhpBGO4rxHyrJ58k5RxxEP5GTzjm1GaChcVDAP1QS+bM0AUqg
OgnGbUib6cb+0bjvDgAXc/veqCwaSk+jLOFZS+SHbPxf/6B/d7A9hVdwOs8MBguPJEwO5O6cMUD6
csDU5N1enw9WDENElmlt4eBE4aAcf1hCrVoug92Kc4xj4rnqAuohSKcjIaJZT4zrDDbOX84Dgx5k
0JOc6Uyyrliie+GdUNaS3rv3jt7+9TG3/7BZsjlr6BiinL/QEHAltI7yXLWtQXKxuVYXSlBNnd97
BkZxH5454pOrwoP7+YjzWz8UatXvYxGk3BQ3VpVd+1GOC5UCS9ANlhVVw/cqzRZ8+UeVhFx2UjZp
3HQLFUkVXKwZ+TMKhRGFUEoSyxjIyOrQf9qJoZ21zoMRVqcVTcThmgLjau+wRZKrvGuUVjE5NDjE
y/Aavzho39iLRs7tSRMCwPFAj5yr2bjLCeS0C5D9GE8uy6n90zD1mg4XJM5Mon3S728SbhYDG3CI
ES91O27TuUmT2vwAdXjcVx+DecVKtAnmfy0/PE2pUg/dG3SR4XR1klZZqODbeHBV2+LdcoZMmTGQ
ezMGIXyMbcJzVkjhvq5xqzcjvkNkkDhEq5aeQmB13gSkwGdQj/owP5PoN43qLf8G3jCZNz24IMU/
7cSGZeaD6OmduYXGdzLCwuB/nTPD4WVnjiYJmUYaZkC9/gmSRLcdFrTT+9ppFCcKwIVGPrGMa8L7
L/lOSjuaal5yRdLC6S7trHmeHCeKQt6hncvnzDx5oNYgNOH7esE6B0L+IB8VOqdKY4CCXJR4qY51
aW8FQBg5jdyGEui0VZfZrs4j/Az0+kLLqAHCtutwXlE7rcQjD0hOGUDVjw6eO9wuaJnJNtEynLQl
KQc0KOHAi4muuBtm7o/ZejapB8Gp8WDBTptBhE+pIVeuxfGD4EurZl2N/R+8zbSjIQd3dO7yVtQ7
mLrFmJ7aHcPMwWddBr0h4KfIE2aevVzaXlEYy0OVqTSAmU3eaKYFdt0PAlDhg/nr1wRCIQOfMozL
foV9d9FRrPw7so66GjVt/zYg5TnUVLDDdYkTRZRwqKSihz1Ar+6CwvfMc1O9HLHETjnTlHGTLsmP
RP8cSGLiZn9sqC1gPZHEWrmPEAivMaJ6ceqmKwwbM6RzIm/uGOIq8lCGQpQHnFAjxuNQ0rU3eRhG
sVutcweUa52lKOZ8daDfSKV03yjDh6bAUs3GcH2VDvVyuG9hA8tQcdkyVnz9FBaL91Xo10ThUjeF
leTP4ms0cyJXgWGjQsSr415tlU/CVfsj7xgjg3cWFoNBCTyTwSejiDYNUUGW8d2Ct8NCbcdziy54
ZLxK85MlXRpGdRfcEL5Ofo5BYt88DAGMgVe60XavuSCoG6szkzOgKuCuvbTyOdXuWRn8eCFYoQVG
SLP91VPxJLuOtwqXQbH+GhceEY7J6Uy2oiVcytWqYH/P85Ji5AafLNElwMJuMAnCgbsfUs2ca61Y
x8P5fdxon9Lz9AyGmo5ajx0dnGjMz8SfU+OxQu0qQR6Rbw/T9m4Xj1O/kNdBuo12CgdcOph2PK/i
i9MPC8SfJBdrTKoq+g/4UU2rrHHaz4TyM1yqczuf1KU94CVLfaVEZPWOkIC4EgRD+nIQ9EqZrZhr
mLiH5TCDJqDhR6xs7z6ALLXK7jcE7pcUqSevOKx4W5HeMHak4lIKf5l+U3HB/Ic0VYg7B8/wfHzR
W0Cp3ssLLD3YmqBVyiquc5NkOlR6ZkDFtsyEXeyuPJohwTTNO81mpEk4phRKcIdSxiCesO6nHr8i
ArrkUkpJe/c3qXYuo7D5I7t99Y5fh9mmqMIaMKZ8xtsT3jo3imbLBvbBX7bf7cI4NW98tEFyxDQ6
vdwrBXGzyCuGOr0tqFak04ifQKAy7Ck5SuIdg7Aos5VQuFAssTOPSEcuttVvGvkQXtPu7Gx1STgj
UJc1MIRjiFgrGF8i3cjweJS1nM2ku3M5uxb31WRZNC7fAh/Eemua8g6DmHmJT+yeU5eqloab8BN0
xv9OyzAZ5EPARdzCYuYBIdg3YhMymJqRYSbPrvwDiS6LmYDPvYn5CUJsJL0hdLbD1MiJ/knNjQgy
mOBO8vqaQktz2dPuuDTfsAoSYhh7R1EIohOKs2KvtrN/MIv3ckTbzvi+IgBmcTR9hjiczLhldZPt
WSEEX7KluxcOsSz02+SSFXhm5gJUAMSZ4Slg436qJAt5GNZVxPng0cuJmpuM6FaBV941+nCmsqMf
18+c8PS6VOqc8243CTA9yQk5L2RSjm80bfxgYL8Db92c2NI+RiyeZEjdDVRwDuVDjUSuxrPgMIVZ
t8ObaqpRfNd/bCr44QOZ7y+FS6dPOaJBuHpmRbec7ER1pDbn3XPy4k6o3ny2hkVcJj9Veo6ltbbY
/eQV44sszX4cKbGNQe+bsId2OoGnmdMLapeR5Xs3Nhk1SvyGdNwJrFiPF7E2ujPezBSvYTmRBl9r
9y44ACSesVaTVb2cqdsdrukJre2Z0UGSqalG5p63ueDyCYLK50GnBerZiXUu2dsK820LqV9bpcNz
pOxhq4iFDlto5F23lh1EpONFO2v/QCvLCf26DGzuIT0ZVtaLhVJHFqtGmdYDTtTOoY8om323FNXP
fRGkYcSw6x+PQ1Ic0BBpR1U+Hhcb1WBn9Y3pHqxqHeJSr5MZcJ1XKzvKterx8WSAlt0WUhY2LxQW
CbRVQnQRJhDPKns7e+kYLcQMSkuopML0g0EKb/sxhgd3/fmgng2eooYsK44QI7Bnp3Byg+moB7bf
Ic/7S51DXGpoBHqeDJivdfftsSXjWtF8G4Mt0SWDXHcY0tF+wQTq1/AuMrhJCX8udaS+f+8uN27e
R6qnCW+gRrktJuORrhJt1Rwk5Izrkfy8Qr1fsXMDBj0aLUZOPmq6kq+4CcFwLryUGXHx1qta8ilj
/G1ZlnsbtNNZ+nIfN0of+aR6f1UZlZbmJt8PVw1j9RAIspxUal/MEbQ/Qf9fwWJ0ehQvLRfrFFqS
KA0Oc3AjiI4YOcT/SrI+EKaX/5hX2SdapTZcFIYAzIH/YwfaWXaUJ6SdQDW8VwA2RemkEcmINOyf
crLaFZFjFXTN+w8HpjhXU+HQAzlpd86Yf9ibN9W+InkipM7C2bqtfyNs+1jZCD8ARiEb16CQYSKG
Q/89eqnsaw9xm4Hc9P0p+0ebU5oMbD07SD/RVU05zzXwaouqxWJ7He3f2fEJ3BMNwM2ZRD/xAQiQ
xUeJJ2MPP+dwMcd2G1Y19UTowT4wVOehxEwF2k1bJWeyFwjol6xQk6Ln5kTWx2hZ3SSD5DsgZ+Yf
LVDV8SpcOEPEbsFdx87BcarXuaBJm2K7M1o8QlYFlYm0DPXxtpZHmsu96Udc1PtE7uzY4ih+p6n8
TdrrS9YiexUOctLIsYOqp620tsH71S0R2EtAdpUtWPHhlkZGvr1758SmGWiMdi5TkTE+waXwmHXP
a3SpSvpRqmgnZ+GCFz/AVrABh7gHf/zNXfXvLTZonChTmFCN1hfuP+RqHdLxTXoeRwxlKysbDYLa
x7V4wxleX2KrKuN2qFaO0tRRH2Osy6daznyOdIoCVFZjVOkP8zzEw4KN5z88+Jsw1GRciOU5f1M2
vImkfE96bR+hv8WJNoPRRLGzO5ZPrD1g5ueEm0VdnLQK7EcAr4GE1NvnXoIuTMp5R5h+M1bLFiLo
4a9xBta515+2ydqHgq6p2YDNbsFKS2mMgynEZMFsb0frxBaQkocsFKdjvaH6nXnmOKt0Fo634ZEc
LFVEEoLcSp61tM1LNsuf4p5NgUGW9q2OjOyrBkmOjUTDBUZRPYKIsfy/XcVOVAAbmr30rEBkICl8
jc+sHn+8mqwhqs9JrX6WWcCQmyGjp5MYR5yTXSNGzf9vBZS3PD1o2UAv5vazngh2VN6/u4aZ4zrj
b40WxdKq7GuFwx9CMzbx3JXQA9ci7tJOCGITHD7R5573Xn5qrkckO3u2/dZtYD02CbCZRCqF71NN
rMKV21spO9WQcdKZEVwQN+W9h07mlga/WrKc7tRFQoQ6k/vRqq+xUO9xCsh0FxY7IyO0MVOqI93+
wzBjDqdDyAChjCbLKDFKpkj5dj66nQqczdLgX9RrO54qYy+rMP7IwuCExb0Wvw0NyhRgKxbhX5CS
/IiHmTtcN3NVn2cCItiiFbDVONPItg2b8rKylEaA/DSlYgZYTIGOKH495xMnLZWVbjMaxc+uOhPa
epSCv3PdHejTo4H4e3iHdMG4aLeOCCHSISuuQODXeQnmuF+0v4pEw5ZgARJo/IpCZlZpHwJtUcnN
6O3T05m6TnnOAWdmHHs4iDNR0aL2dtt2aHDvF3Mkjqb2sWp9iJW53Tb6ASvyHuNvadlQH7RB8Dbo
eFMT+sTgJZAPSU4+62DueO0eeV21ZXam/Orna+Arflw6MtaidkPLdKx/z/VI92pVKa8RGOijEHy+
dYBSaaLo1hl7JtbY5rUdRXAt5v+dSip2xII3hOSTEsCFRs7V6esvKF40H7Dkz6pkj760IQQG2KtW
nVyuaN/T1Ma/QIfUeNOeeYdThSmfPbXufyeLTFEpMPCFbCTQlrUi/EtY296pqLNOjgdGcokEx3tg
vZgE8srZ0yeHzbyBKslqNCsfX4TAiUVRT/Yl9Z08oYga1sj3W+K9ZIU4WLuqTpUudz3SdLNdUAns
uMQnLQkzRI2UkR4ZWE/akSCPu7xnyt99eKHG1I7TVBTAiMu1G7FJu25qVhWse7Ao+zl2gVH/qs6n
55c/fF+wrwocTN5ceKg+r5pZFevytuknd5n5n1WZJMSPfTZ00H9et4KjNjZrzgpiE42vT1WSVRP4
UDCHpawKQRHaWQHdl2AqwhPkISx/XUxPk+2irVpY93sXHvGssSFb7e2L1P+/U5qKrdl1PvfMbjbe
TGV7C2UaNGnBHhxaLlB9JK1s0K7vQ+Nqplp9ihjKTUXX1hbPd/vh0s8j+nb6FLd3+TJp1wBBYLGZ
fwDVB8u35PUDAh/7vYt1661onTKdTJc+FRgwf4VVWecpN9JCZUvUhuhKugZiVSygIxqmhzzmGIfs
punJrkUvfjQYYUMNmETjd6fTVqGTBojU/awGkrXaG+VfaKMwNUnYQCwkQ+lxXrTjiiqTuf8ix79V
OoYlNC81bd3EzqW8COPE6wP6QahVdM0QZnSJf8V68pxaubJ2oTVPoXuzZNahFwjGvynD09o3iQFZ
X+UmaVCwt3vOmT2I8jMjeFefsvsMyHRev6GSE150JkGoa5w5tDvVoXVW0KpVZltV0WiflPSy8QKO
omCr5y2qJKLwS+vd0Os0N5THVGt+IcSsHCUzhdD8MAF3mDYkWtao/0g0mFgaGj+li+NZfIIl4YjN
JC/PmGUlOr5yNuaXIDH2MJNR+BtA8SXdGgwwwtDe5MAJEARrWYOKI96Nvt034wIIXExSbKQhvSPG
2vDq+7ljrb7JsRKXiml3HNElSWCfnM53RcaAdx+8Eu9tunaTMg1rQ5a7JSY+mZkET5AbrKXxtziz
IZHiNZugZS1M5OLl2aejIKoxxeIBuu3XuvZeP/jOB9V6wh1b7c0/9cEK8aDkb0inaugv8sJDcp9I
03p8ud69ikuB7m6+Jc9+EDeaImoPQcnSheCupYo3GdHhrNm9dkGEGjVOSnN/Qkl6hhsvOABvM70e
ui4rUPjRAhsUcZpoeiGlxoAF7Do1K9CDUG/W0U1kC+zaQFWOPjTQgBKNCv1EQcXKFNhaiMuYC9D9
YecyAzwRy6AFsuwYb+UB0t/lyGw+lyaKMQoomOHhjYitt4xeR/NvdPRuK7q/yk87rQ+8doHg4q46
mEc9osSkjjVm+My417pt3L+wXvwD4dx9orVbMq+kuwqmfFoMNr8jCdIVL51Mx/wgxd/Sc3H+g0rE
xTuQc4LENds3mpJUYEtUXfGx22SSKG4SIds43zMUk/1DviH5/T/xrlWdX3ggnIFGOZ4yz48GlBRu
i1ErFUsOhEAhrEuKWZYPUE8C+tyjx47MIRse27TYz6EEW6RqUmGmUm2v6v1LZ8BC9niNXoDqMyqt
2agf1mUUhlHsLmJqPW4D736jb9TZi22qB7//oNKaxQ/jAace1jYkd+q2wNZkdshetXgoy8LCl3dM
6qvamMhwYw7l3FA1WTOdQiOfPL6+X3wT6CVIdY0wnmThEfGBlgOcWLksT0rdS9qFs/e7K5vC00oL
+llHD2zj6Ny2jyqg+PDk40jT9EzMfuojBk+bH/lz2VtqPoqOJKi1bt1kgeC0eGFdAp+HQqXP9qDu
o5y3i/mNF2WQ5NCgzoj0yZUUydcQuvGlBZ5GXwQhM/heCqBU/YmxDHQAAoBSz8KBr3VHVYzjkmi7
f9xH6UXlylA0nyU96EwQMdBHkw5XDfcNG+4AWZfDigIA702Wo7f7FvQyBkBeijEqi/fest6kP0Pb
LLOhA22fIavQR6Tjd+L2RUkXoqQ4ITmXp0G7Fb6GUMnMIWmQ6Ik5NHkmqfysQyT6IDrsY0Is3500
sZkn9JHHACaLQlU+pe9pVC3O2B+6F4XNRk8jQ6NGdm4F0AxW4Fw3bjFNp0uYgohciq58YUP5Z2Bj
KP1XjjuMLW3YJLvyMSi3keDeEruig4LwMLgegrw08XVruGgE7q2+8ELqm8d9K+W5kjn1fuh97Q+T
cfimxOMeeR9zffKDw9J/5+QUbuE9OwN8F+e/jv9fQ9hzyfuQApVhC54s+x9jDrXR6mjUFJcCJunE
vxogiaxIgNQ9dfJwWWuEGl5FnLiSQ8CCsMXZc2bkxU00odyqXAYcTPj/eLVVHeeDNH90dDa7OwYe
w0h4uuuZDcQlpUO++zo7S38SglYoyqFXx5dB0GCVJ853kjQ97KLgAANaFnmTt/I1UBcyNi2HEfkl
61Y8WbkumytenFnR9eOtjS3E/aKlQfiRHILBoCaOraCYpO9u/a8i3MzXBIDDwStYYmm3zAY8XGH3
+1xfZOC3ixFrH5YTCzcSXVQy2dGBwHraXAdrfI82vWIYrqKBze7/DDF6/QD2VdSRFLjleWprm6+J
imzDQtjzusMhE5FYjuCc5EPOI6kpIonCEh9igf/L9mz2wPlEQEsWniZlODFcttbA25ZKZdAEn3hB
oC4CCvtXZyZsxAQRCzs994swuohNrqHuXOATam0bTbm4lBfGIUrSTlv8llL3LN+hV7NV4negsMbM
osjDKpNwu/0NApIHb6yqy3QUDczGdXcSwpUx2v9IEM0IlRXgeMeYxFbUk2hpdCRvGsISc4RAYapK
sTM/361FBT7vMTWnbeT/1sp+Xf1Y7Io3kXo0eUoZa5in54NdDKBndmHlEAuqjPFhi8TzF1P59hoq
UPa89iviz2vNzOXFVu+x36wQ7jOq6syEZQdJ2i8wQOUaANF29Qm4da9801X1BWhExAY8ef8ZFiiy
/Bl9OGlb6QQCNF24jxaFA+DkwbP+fRQfjut48CBeFvYvCAhrh6e35brwMzAwWS4tSjLTnwc22tso
yfm8TRI6KFhcI57WHssOftsW84ueu9ZIDsQFE/dT+DRqCNZ7SMdwh6uQR5GEwSNZF12cxYiikV6z
5yan3l9tf5jOnzBF463qPH11V6yj8aMaLO12Rw7KTZxQKOBaf9rVFgyfV/LClN2x/yjSeHMBCmLa
vi/W8s8b1fhpC+ghkaaYCrV/Cr7AJK6mlrpLycqafTYFDX642WZyHB/D3JSFmZLvibrL4AxJgNP/
YGLr08tMdnWjSSWna3pPwZVrgloFy0oeTu89jz6Rm0AU0F822lhpbeiLJDcyuk3Xek/4fuNLDy90
S2fJ7g8cY6YGuKspf12RMKVMYJwxWGhiYiVRRPQLY8rLqravuHNgF8tOi7mcdMvpmrgYgfMN6bOi
kUZ821UqWnUdMnHrNrvq45/o7h2cEQIxWCaYStVNFk6ZVkiCOZ+kbWJgobBQd1vj9Kkj+rESIeoc
zYnjacUrn30W5RFMRPxbC8g35IAiqmj5EDm5ZL2Y0BjgXaooQRVnUzu71BMicVjs1WuZ8rM/9RYo
pUj+3E55lyFl8MScFUlVyj8Wsi7C7UBGfd6O5h2rjXQebcPdmyQiRP1r0Dkn7ijTN9y1USWHtAKT
IkkLsaXG+Imp6to5Smcw5zzMNeAHprKoBr0piMHDvGAMIGmRI0VwFWWrjap2X7fa3f4jBg6MsxuC
HABdQpcw12gxzOYAWuBFWMlGw6BsxtiVillAfYmymdP/yiJcHF8DOTcPNjaonL2ghgx1GixDuT/k
83s2WT7ja1u79mtNFocjvE6QJf3toHwan8Ca4ewDLe43oPwxHCKKW/ilL2a4aucVB63SNI6VoXp3
nJ/YGBlk0/k+5dxgA4WRSV25M6M0cnIt8q1V8iYFVOXQoD3ePTKK0Ov/hb8Lnuzex8z+P8njFhpt
9vD5UII5mIkC2zZtVW0cHqsz888GVnMrVb0kRDxAq0kP35MFJ45ibw0tb8/vrQfc/hZ2l20STwi1
26R+BOj8B0wPWVebyOcsWsBI2Rb0EHhvSsF36hoxerdjUAkCxgOpNX+GttfOIt4L71i1NlQzCReg
pXnOd00gLMyv0rywCQi4aEj2HyZG6oSIne0VRrCbz6xpEqZaHJII7F2YozkWxlpA3AIPUm0G5Nhz
59cS+d8JBUzc7WGg+l4bQ0behHM1sGB67Av9eO03NAozfy+4LfSJeymppCSEYhKWVma6uZscyD2/
amGCoL1/hHA055hxMN3g3ofqKWwAvbG9ajZGoiVGYHZQO6YBndAiOEgOShdIa0Yzz5hDybc9/Xr/
DLpW2x+dnNEiaHQb7/PQEcT67UAG2aFoF2K0qfbGXk36MqsIRzzqW1UvW4AIrmolmM1CXPzMVICy
qS7d9zd0P6yN7Xk29eomNLYDbsQXzDp8o7meuFLo9PnkNYnLjWbvsbU6LCcSWlKITkJM7zOe10uN
GEkeFxRbhNMHdNj7V2R5osWqiUA2LTOmLyokD45JzpNQ+JGTZUeFDDR7swAMOstQTPSe74tjHQa/
kiMN5CGSAVnQdIxRb1CpH1j9mq0IiB4kRRMyYeCX7cFHqB2sbZWt8Nol09deN3A26P9chFRSVkZ4
t5S75McvyFm4yLWM5XJz5CO1LYxRSW5MTS7TMMRYx/J/QrujJLjrsJAYn7SV+7vVtDQxwjoshQO+
e7mO0AkG0CC1OiCI9dtT9+vRJn3djtpy+bWb/VPxWMCzyY7vWP00Rbai0coOlpf4bP2vuRkEWqwk
0n08EcgxCZY8Bow0QFuXXjZHbK41kq4r6CH/3QO615i12mRUIsGmg4+VnGSyTo0yM5zDVUAsTx7W
9n3Cd4zVzcd2lA6O9KkJHTdYUWJ7YZs/6a6cgLbdk1LUc6DAoCZpLktdFYcFQu8S9Dx45rQyvOhI
vda6w7iFH7NVGquxGv3tCTN/8afUY6kA12Mv9x1mnfAOL6v+GCmKcPRGs3nt075Ho7rYaupFl7Ie
8FFWlngaYrSvPsVEztX0DCJTeJszaUk4WWiZQZAhjKiUeQATWBsIkcrmrbkcMdd6DS/P/DhaH3qq
jMNl4Gx6c2B9VkFH8XX+Yat59yLzPvzcqspxWC9QJmY50acgYnnvBMAquQVGwSkl9wvpXwlFVMJl
3CjJtpDdU0IbgU5KZewtYRvEmLSvc68n2lwAc+Ffe4bUGv4Xps2ORiLQ9v6dxDOl8ss4QV7dwFCa
mHCHHxlrFizzXeIkR7Nurv530IFf02QdqaMFYV1MpZrWyDVmpE8RGsbaic/VNxdrgpMX6ruqI0+w
3y/FZUB1ybEyWYB11gEH12Z7i1piqOSQ6+AMbZ7jmLM+zHNlXdO5m8jbdM8jsfqXrk0sFPJmlf5W
UPuXeZKtJNj35zvIeiRKlHAm9gXn9khxWyfRz+50imaO0KTqu/k1KM14tNOtoqG+nVZlPWhawyIV
cJU5aRagUIIIc2akOsfsunJaBFBGh7laMKiKptk6Tk4jRqoT8CxpESEj1uQlkxJQDvLZYsC7HqCi
oRcelvJOBpS4MfBfSKMFzPAJonTkTyNlELCQnyHxJCxUEH8eK0AIwDWnr+Sbx52NnZonO4NeNy90
U0lBm8xLMMRjCVMOCVZqbPXswBjqzybod4896GsVs52ZKR4+XJt/wNfFiSPpWcACJchjpS9EYIZZ
ztKFQyEAna39AER0C6hqZB0RWCUdI+O5AIxnAcBhoa8HeHR2xKLHOCCqiRz86rNfPHTPGckhMj/T
0R/bljK0Pn/baTZX1GmAu1f1pMZY19pFXh6B1Dlu6VlAyNiRE1aAnNo14xCErw+gqXNge0kIIQ44
T3pI/HWYL9g+Eu9eCE3NlQ/w0byL+/Sa2qHqJ1YGUAnphBiHTYEbxtjT5OGq2VXG0NvMQAM2qRrT
9frVX8aIg6mygrQgrUqZAbqPq5mtPkVg9mzNdNeZel663NJ8GM8QfMLzTZXDLpDSPy1AF2e1SPcv
K6UJntAiwG3CDPQYEIhGAya5+Ctmj1xKlClABX95uiFwAGD7lvDQqu8plqZPN8xac+flTHC9kgD0
CmZajOsr3jzkSu/gOIKzZWOjjpfZ9d/7wbzBWGCgLQ5cx/iF4d4A9rhKCEOrjmwhg0pHat0MuwHv
GfmJO5yuuFV4Wq5uHZLr5KzJc36wM97qbH8DKL6HaRHojyDMLHgFT4ByDrluwrSBtVUK/XJMXm1Y
31gCr5KTHclYFuz6cdW2sa+LS0LdGvKUPRsltt+gPMNgCRk/3TF+W8PG4CYZULnJctOCseGnO0Bu
y6AUFXbkwW0nVodVAcdozB8gmWgY2kkZ1PRs5BIYK7Qy4GKE5yBNPodK/nBNDRIqDInKFQrBRBzQ
8X1MFu1b7ziU2GFfd1/rXEcmHbk+hZftHNGJF6+YwPU3TNHrxvAsepxs1x8f1BziTK1ygOjX5qSC
hif+pcclpnuxeF8LAr84K56sWORIIdGZSmPhfzqEdJMFk3ozhQCMB/yKnNHrNTxl59ZxhDvGC1qV
Ez1e2j54OBaryo/gh3OYOQmSikqflS4swoQaW1kydnCEImEAwKGz+ULrh72IPf9LQIePKKcu0e2P
85iG390ksNT46xJpzvv9/A0Ssc2vYRSEj2nsR5H3QY6MOXiLS3PsaqSfXiEfbmfiSNEWdVJHJ38u
1t9qHHx3QfM3DbJv0uc6NH64YGTr1kXTGGs+UNO5xvzbzbwHh1JGlyts9FFVd4vSyz+k2vyPqw+2
rzbBG7Taoq7lwGKCprZVkysz1UdFBiL7Bceg+jtlXR+bKZbEDjMMdx1QpJnDEWiASfk+tjDGG8x2
gUHuGuOU6cUzKuT/L+xvJBvpWh09TFNN3my/2HuNuaHFS+2+vmh3okeLjndMNlqDrh94bfUpGkKL
ktJEQ1fyBL1iZLSEZ5p8aTSQ1WI33fw11fjN/8B7PO/eghRe4e87qEfULetc8S11Ulh+nraHiGkh
CGvoqHs24Qi9Sch/cD/BZm14LnGRVd2f7hQkDowLlVrQ8uhXRa3MpSlF4KOngaYMRYUH+L8dslsg
AnsuspZPvajJmFI4rqXDeLsmhxYeuVl+HNXYQVm5MHz+yHXd3SmSTsAGpzGRipse1Z2mc/4+gSpT
q3vQskKfIOH33BwwVUDKQ4IhH+SahQ//zboXmhsc/zh+uiWKPdqaJ6yD/L8W/qartHcuk0/WN583
w1UdCOXQ4AXr7B8gWDs9BSvJObrzeq0rEBOQP9zTiPEwos7ZlxN1Lwubc0v5KZdVlhdSZG3PaSEm
s0vJXFGeK0dW9RUq9zYHGoRpTm1JK7irssbiclTqeCtdobAprhm6GayJCf7y8+EZkNLUBeJzVUqD
Gj1X+h8fXHnLjkaSo9ua/Rb+Rh1b20zdAYddtG0te9gEfXKMDVQS53ck2hm1Hp/hbbNcKuaPHUPC
oqEAiAoVV5bMV3EPWW0qrdaQ9tOZ2hK3bMKbLhgb3yI004HvQ0HA/2+pZlvoFQCauBTZtsz2WXdu
34bjgEKf3bD0GYfSFGpJ35c6U5pyo3shFliZdIUl6E5ezncwsqP64bSLFDn3klJG2+j618Vj1H+D
mFwTNBHjyJVS4W9H36jjtItgm7lrsxM4jmkjvuNtwnZhUqqImT5JLsHw8ORTgbq6U4nlNvYOaK3M
8T+4H6SJbGYhLlLvR+g8mKKdPox11M9pdQAvcvCoMgXHMCrEhqujTp1GCNpAgJ5EVfrfa74q/F4u
uoeWp0iP6+DP0cI6QaDtByB5I4/WszO/bEA8ZGPLYAZISeLp53gMoinKYIx1rHGtDeM7MdTIHSN2
8/8BcJqv5aqWRkN6g7i4DPGXmsa7TWZ66wGlG9gPF7p/fFfQmQprUGhZObZ0suXgRZvVY8nSxa1e
6srjdYcjzgo7lD8WKYKNPNfijAW5MsHEiZcw3UgcycBen+mOCgGI/ZGvmxJ+remTYItIHR922xJ6
APKWA0ICyPPlXPlMEuNYemsGpamDfsBXHrEsPZOzEs41hPKaWf7+lkvooITcCMyd4PKx8pUkCf/4
J1clkkaDVBi0CYD0yqlh3W+TS9qNYwxbwWr33QXrTnH3SSBANRPrAcafHxWU0jG4BLLCGLyKsOka
733efVWNpt5P/yQ2S1l8Ozauw3J7AIOOJBa5AiV6/eKuZ+p60iYmp4H2nO5Boa5F39NvGo75c8Ar
vCvdakT24PwVBMtZ1IeaD2yjlHD0Gd7FZ3IWnKAz2Y9ybaD/2ft8T0W+IwHdlBsUO1Hyunp0BaOm
D3IM8HckcLibbMYFnnQlCOVYQyH4xcdSSH4lUAHDlq7x+4Dq20klJuvo6yd+81NEZay6BDt+ITnL
0d4VI+qyE8Ipb2B9roTiBHPhuvd3oY6qnRrGstmvCNOd7KdziaOX0y9t557o8lgLbdLLECoVOwIu
pxCzUyOBOhX1Wp3E+kS2FtLNPOQ93yxeFoZ4Afj6Yl1OpCafwML9uXG/xGgz6uP9AyyhJCBbUycF
z2d4aj0fFhqugpkt8hmRq7nZlwhpfxxxXon1246dtYdrWCCt7HOnAawzGVAPON9ArWl0AwBFQ1Oh
TAxPWJen8KfxxRudPi6NpGaM64l52oOwjwj/LuEr4DcMkj4SRv6WRR1bi7b9KeEZzs5lqTXjDGkz
sqnYnsRAfwP32FOjD/ZIOIo3luKnDsVD6ZQehNS00h12Pfh7qYlC85WuBst6gx5w4TLnUjlhoABa
F2x28CGqtyR9tDtrUKdz/32zNGzccqUPALsvBxwAw5WDJcDzSDzTs1T+fj4YSnZ5FL7CUgVkNuMF
DsNPHagUHkI+16E4NSw2w4snxUevUkiHTkU30YDkI1DXH97Q4oF30ko7JrsEcPbC/71OASq/H6Rs
l6vh2/tvgFC/QekbgCPc/XHkgodO4HRrS06o/lZkBFRkCQb4RthrhxvEsltYWXk21vp3UCuwu0vL
wb86J5xQR4vO8MuRDTtG7miZdpHlRkXgGelV/NKp6/x/MMeWly6xnyG7jDMWxMTPESzhRTEE3T+7
eMl2o0PQOvNX17pJIZoWWQ+CWvBvCvsAZdlBa4MeCLdPpeyH/ZCNRKUF0Txef0qYCkZyPV2WGrZk
3183hp20V26DwWimzmKqpK+kdMEcNtMVVlYr31ecOgLxyVMccf/NLzIRnF+vk/R3VEzC+l8/dOqB
EnPemUxoJYqbmwmALxKKBeOu8RJnUdMUqN6fE0yDMIT8wQmlZcLLYM/LcYfNbN/M2Jn8u1q0Le7/
eaqdjeqiN3CF1YlCdbAbAlDUwd/KAbc31XBV0d2q5d1qV8j55piOSQZ2xTPHEcHdCmaorXoRuVZ8
BUK/fedTHG7DBkClhhlikIHPdTwfH05DK3FYiQ5ibUSyi+cGkU2927iOe7s5POKHr4AXxYASOyOC
kNVrnwIFOVBXaYfPTVShcxp1E1ox1Kf3kv2hUmluPZmdyJGONuIOai4D09jG3Qw1vyVBoF9iU/hb
gFghnDJu6pb5jL5Tb7naBm8ZuyS/ZvqMX/cjKpzwcI155ybaAJ4EAXuJnbfO5QoR1nX9c83QR7vS
y8h5j7jPwY/88b2340otIXHP2KG5JHw+f4STh5ekO5t0fklrNtiGEYrnOQpemfxLnMI/zdvRCc3o
XtR2+rHAAfpN7+mILpXMNseTJnJofWyUSDawvJZVhp+3Xuk1eGyTLB4HY8m/pZ+yDbiaTapjjgVK
jCZCVYwCh35x4VAYGpcftXHmYMZLmM/irDc3yPSDmsUMJXPDTj+avOflph6pmFuC2XQhbetk95F3
NU/yaVRtoPgaeVrBq3JNehUCHkXsZkkOMUGu5wrYl0QAFmePsarSyQjIjZeJ9VNraI6IAX1tQ6BB
zu5e9wR5x3KAhj/JrIEbibXuXItfh9qgaqn3S+4HsHdFrRwkmOaPgF2bU0VsFJEEBGehU9G9pPEj
mov22LAqHln0tZYwygj3TbC0ISo/twXqLnhd6Otvi2CS5xAa/U7RNeACTh28bjOoUG6RWllXZMvW
02f8Wcb+IeqbGKXiPcszL5SrfUJQNSTNmE1ku256aXJPDUmzELQFCfsVqQMVHcJRS/IcMDFW4Z9s
zUK7SpYygxWolJit6Kf8dGjshjx2HuwY4aMbNyyAcojfh3x6doQM77FhxoPhwrzLQMhWmV5cKeQn
SPui8mg17AKAmxpOdNdB59xPEp0SPM1M38IDEeMhsLI7uPJAjQj2UIlTg6g1Db426yvqccg55h0n
soPcvCRNnVxRTLakqPDGm5j6LLRJAoDoZfmAoMcaY1H0l1i7gvOTpMOVq8kEwdsIbmSLVUdo8xQg
NG3In4NL+CWYJYZtCrM3V3HmrYMydHg3CiHYIWawzMPjfHkAOlswrcuKZm7GZpoLpW89jButAhut
FeHDGwUqUvYKcdrx6lFgJTWK1kwPO8GuHurqNuG9Wf246gwoPM0lHrD1jY8+JJLv5i/g9ji/6APL
fxKLqeYhEAUE14/L13+N8/dm7l4CxRrCjfbcgF4QESfQgXj0v4Ofhs6SHQTbmhPEie24HRvjIesW
CtNWb2bD53bizKJ2bt7sG1qU/E0pnAVTsrRkl/NxJ3PgFcHrNzPTU/8ayIY44ExHsY79O9ASFxiS
RsLGEJ1anuXvLZuZUxKwWzg8rueQ7/huNY9cLqo+RURtk8iIA3Wv9YOEApFLI63EE6dkQ8gVTS58
6LDK5C3Ad7GgPfXXmcW3xFQjsky73dhYC4PRgV7aKjlk0CcJMBxS6vJcGLgn2wDqCcqf9tFDr5eI
vntml0MuqzcZdqgLa3S5CganEGR1PLKN7ZdaZjJ9iWulQbUkQ8biCzNqtdAR7roSJswP3koiD/Dg
+skAAf69x2DoBF3BgCuKMxSvxz0qbxkckwYKRRrCiYbBVjdJIRexYU/G3bY2Woyea9waHZ3PKV6G
IqY8Qz1g1Zcres22qHRxX95pVhnEafxti4J0zUt4EfGlSkOR0EfmuvxIIEgb/yYAFJye+LYXr+e1
ZttCiQKVu1JcGrj8izv+GqmLKjqxp+mosELU2iY0cYz6gn7m5UOxQLDfWEQ856YcEKLhc/UzF2hx
633qCEtqNe21zhFquD0MZYK3deFm0FDWJp/6nazsjFIdK1g6AeF6Dimfs76DDaxl5hcfAbEt6JcJ
9HEvFdycbwdi4JTYnxqWoI+AGBB6j4T84hP04E4XhEt6tuuJZcyZzqdwnA928g3+Ix/smxMleZTt
gRcGZA6YK+4wDX+/N4fSBtEG+4xMVwaeIducXeKmhJNKa9YaBwFkeM7FdSTJzdH6Czn3i+N8bvqH
vJyghU+8qCMl4ZowqUoaSSEpdY6rwDKuoP7cPV+AzB2R2rxM7qkOtixdW/+ratIQDs3IWBy7lfcY
N+6JqlAFKt/YIO3csThvh/LwCmVjYC+nq2teS0UMf++7EUsYIkakG13jHx7lg1ggpCmX8OE65fUI
D0pQJiP8EcSTMChWFgruHhM1yH3YUqFocZIeqFlz3IrzG5LkgWb/9wWqqWMA41PZIjP1rc9W+A7W
hZFXtQWgmSDQRHeKK0SPx0M7CA/CTGKknPOyauWixNhDutJRcoBMsYPGm3MJOxpGZMVLIkPl3UAf
vm1aCtZNv7gc6e78IxjMM4BYdsO1tgL2pPJ/Nf2m4jpzP8FJFMKgRWIiBVboXZj95d6qpS1DTpSN
WitPdM75XWGybgLoVLYlRYufge+wDERy1I71oAGzlWgHEpP1cvSk//syQ0sNIU+ntwOpctRWIOet
oMiFZHBFu6XfkCKQnoNog4+xLAd9uUrykZhekrgnQOM4UutZLOJri6wbd/hnncsn4lM70EqPe0C5
yMZ4941wYu4m5mtA6PV7EHmlqMJLpfpA5W71Ga0BK5G5QQiUqrQNW77HNl1tAsOGs+BQGgIv8kas
ziDiU9OPWwN7isA+w8vKNOEdd7tpj5EvE2u449J3DW8eRQuu+xaiee5J10sR94hI3sFjO1R9OsQ7
4yRNxxZq18DjWZWPId2uDZgwAQw8AQCvdMozckCXQIg91Vncuz3SBrucdkxHuXng+D7g5fTyJEOx
efkpwWdBLHZ4hce1TQr4ZGb5LjVem2aCNMVq2n+RPQ3GxA5wBD03BLVQVwuKdXAjvGBEMuj87vbn
O1hVeiEiGbeLC5+p/twvdQP1m8q0CCNlvqobeRPZqLvy70bWlEJzStfqocGtzSJ2npw03JqtfBAd
DoL+za5L0tu20vwFvcfBukSsMLEPYnaC3q0k3mOtctKvpUG+y00SD2ISyw9nvFWDAlBl2pxVbcOO
rUGOQmtCHdL1HyxX1wGsgVBy/Ea8FOSz0yPk+xKZ0584gAQL0UV5zfyxGkGiiLosuo8lAiigBiHW
SrjzFD+EtqFptYCxeNMmH/hr9ABBZPkKyhBOCmN4lxg9GLJyJy6HPiM2tTd3DKlV/vCp8YROEI16
sE9cJgTdUq57/NALujQFXTeQLjTECEZ6zEZwc3brb2WWf39RbWhl0g1jQcOC6S7xPY9GkHH1l+Te
Pk65VN0NSDrgYbKbBIpsQtTWkWNF5W/cJcy9QAgXGJyw/y7a820svMmGfSywrphNjnZPxHORckT0
L/NTaVMzH1Peu419SiFgoq3RKJGajLbbKViiif3bMsKzXdy8ABC9lp4soieI0SBZo4OAiuzqOA5p
OTxK6neFSMhSi1GmToVx4yMzfNr3vikAe9KjiewHEm1+Hz4ovkHKSuv1wU1HXccCIcpm0I9LJCDg
r36zVeLS2YPVAnD5VdT73LHkcv8HhM/2RxpyvtPFldOeHGldTEXDDo4gEH4omg4kkDTjqeIm+jlc
XTSG1Nme+pVraRN8MNOMXPH0NZ9Y3rmVRaThqiwJpX1+wQKxQb4IT5z/iUIzA7rQOllKbJeCWjPs
UeNmV4ReS00bWAERGPe4M52a6wJsq3Q3yUYE8VhiBvMq5LdpLgM87pJLgBEmb1/rWumuvbaafxKk
65alQn69unANNM77Bda40qxTcQ1I0BPQ3BhNYOVkkOn/9le7hbytYr7n9buAhBOhRJxjFgswWCjs
XbU0hc56J9O+DwCRG92r7+5J0Stsq1hRAEU9G9u47kBnrKgvLnbrvkJlsJHe/fu6MRt8R3yie4+x
ywOaD3aPakk3ZzViGzQ5LiZT4bizA08w0Pso0UTnkGgjTxSIPAPq2xkUrh9Eat/Wj37LLSnyaGCw
RyodYEcyDwR+LTnujk1aLIQTYNyVR0PTctTETfbDriezx4I0U2GCwFSc9e5WY3lw6hlPayY732+8
gqPT7kS3C8hEL0vguA+konb7ABDrzvK/ysKWQwNoQzVSh89zwg6zivuIDr65OFHluhIt3CksPkm7
WM+NtNsI0qfXjRxItIWrZnETghbatGjLUoJizv9sfLmSUlOIqydDxUj233aRxGnFXHQzzv2GxrLu
dhVvZuVNii30y082H3h1V2PTg/L94hoDwTM6k+y1Z10KDbptTih/CMJMIfgwi7nwwH8LJBTaQLvM
YsOr3v7YVfRWwX64b2IuDOjAAdIHrfXyFW/Sl3hNQ7urfRM15WWKag4UBjPHrrv0yQsNjtV71EBz
6U6n/7SL8Sqe63rVMIohJ8WZ0Oqda5pYBRInLsRCRbX071HI/14Lz6aTShmhUHQJ3TOvVOvbI3q8
uyvzWqYWoGqu0lQCbV524tX1KP4ctIiMNMcMMEZlFy2PrprjP0m7MrfLBrykq8ergkxsBtNRhic7
wqPFGJ66MZTaPHzQB2ZHi0AElnjbXANT/iwHI6zI/PlIO2wNC1As1J9KswgqY8t28rTrOR+DRGs3
6w3+qaSKrjEqs6cRQrR9je8WxeE+7PCUwkDQvrE8RnxvY+h/YfW5co+Xrwl7K9n9R14c8Bx+5sPP
HRdYFy55KWpE+EsgkXyl9k1e+XBI3VgffRPxKukifWbAtBEW4jjaQWoW/wBhvg/prFJl1HVGlgXw
4xUtASdbCSPTq3uXESDiBmd/kLtNi4mLF3amsGVUQHg0fCydAW2EbEMfPvzX8fGX5qxXnZ1KsSds
e8L3YcflsnNddwauSGAhlw8wZnHsfHBfs/N/prOLWMN0wDHOfRqJG/+2+jsA8AEXttVvQe6zuw4d
74HFFJIDsHpIJYc/F3YciW4gf6647F6lSWwgR1nBw0sDznetabS3gobjl7c3LeFSRuww7zGB4Vu2
pbfEAdCkJn8/a9AfAPMerHmeHang7yQCbfLiA/raxY8ZPVY+/5y2b9mbUPFYGAuat0nGluEkrnwu
r6McyRVxb5dITnzHrQ7OxgKv+NWR12DODabTSQSNeGHB6H50cAKba75U053ev6SxOCaF3RnuvdXO
kTy63ZIfbPnuWMpHme6TIHCjIvD3HHReMHlfB48rSVtYJGxSVqFamZugjvyTmGkWfjUQOJJ3qjyJ
aedYOI0J7jHuao043WaQf8TtBfXkJllTp1AM5Dc63gZD/tPx4JoBG4GY66loxKVVysThbVmd7+/3
mqmV2YYotjvQZCjJe/Nz8Q5YcfKMwRDRIN9j+YnZjLa4z+x/3Tphef9Wg4RJTlbMwgIeNJpQEgGl
ZgbNdIoD+TQHFI6ViXer3Nc03MLfAH6XknPmSB2t1M+bmjO+o+m/+2B0uDj9xlYRZl7S2bz18XS7
Xa7Fgz9OocXTuZ5esqD3hdkgESd+0dh8Ufpu9JmIq88IqnK1xDMzl4mQqlc8nPmtUTuA3EeWYVgj
JSab9VWz6otWB7f7sJvO4j/KyNEsA3ntL0por8iP6fYi+mkBDLhL3LEiU7BXegyFQGiDIJNtBHqb
yYtvHqSnAZybUGBA3CcupAn12MAVMk8eXNqSIDNyQu3PBqHT3t+FWAFo744dsoO2T6w2IvCo6zoI
2msFdMHikFwo4VeIH9uupiEoL18Bha75oxp6KrBJ5dVK/FUdCZigzaLWxxNHtuA3KN7o1o2lb5iF
ioayMrhPCEicnvtLeDvsjk5Ig3pmh2CdjtwWfjxTF2VFqgcyFubZ2012/7tPTifkg7eFKYFmHGzx
RJHxDSiK8CPbWTPLSrtJWeQx0tQsZ1ZA1loEjb2tTO8S9fp9i5rGjtM3SHJzmoi4wXiMaRJmyaA+
wNx/womvfBhyFeuEfISkItQ+UNQ/Fave5lj0BPjgHEsw/wygBvfiaEzcW9Edp/sKPTHWrZ7LF4GS
Nz2YujiCXcgoIj4BiFTs9jlrke0UUsonsu8frCF/BaCmC7qtkboqVreyYjvj06dWtR6cBEsY6Jhr
Eb2/rI9ouZBTXJMqxdZT0G2HiNIbi4tI+Gu25fYEEUMhwbBOAUHEvZzT8IJ1zG+mIuMUXVZINsEw
ioZdG1V4f4oL7hIu0YF2kUldeD4gMrYtyjNO+I/S8JFkEcmQJWfinHWrh/4XFRXKdYIe43IQ619c
jrIqzOzSDU/ci/+P9j+3762nERlaNPLvUeawpq/uLXAW4oOlQ2RpYXFBh0I3asB2BNy6pnmbJoxQ
I0APvmTCLgUpUF52urlsKSOOafBWtsEJk5kyM9Bgt8TONt24xcGvL+Am4YAh6QYCM4vKg6tCCT12
g0B3pGPamKhH8O6z21KeFGPCQyMO8ipKLwkE0VTXd23m7aMTrmus20RwOqRatm6tVTuvDCIOWcga
iIzwsWXWUCRbUHbhk8Xj4PaREB+RWtGpr3/Bp4u/cf0Ttxo0mmWjCwlqKERj3ngCqgxwdvlyKVcy
1WaQGwOHZmCwaBcaQ5gDZiZF6IWUTP23Fj2/GgTdPB99RWT9SVFtnF3bWWdeD90amFlmjvgv/dqy
c3qc6eJ5B5jcUpdEoCxUHT+drYhINRfrQ/4RnpCJOGbL96EyJc3t2k5CtPzp6UUpi8QN9Jhs9p5Z
DQMXSN3fAsZalHeDvZ4X3WUBszYWqq2429TuVTYI3qf4sUn8/oQEj6YT28GBnmdeejuHBdODr4O5
U2x95GfRPF0vKKsz870k19KU+a28pfDs4EBJsU9qBbRX0O+yAP9+k7+/ZSNzSXgf3LC8efmz24vt
NwV1hnaaG521H7EC+IVCIRDz1RMFTgCtnAcz8BhObPw5wpdveVmIew7Y93Bdtkb5j/TganIJF8q8
OqerHZGiGoIVo7EYS+qJarJBS+B2HJjuG7WgSEplS1c+RZp34+x5rcMcIoXLCU5v1/TSm04ZZYRN
aIvtBOhRzf7FiH9gnN+1KqlohemqRNsduxtpMMaiYI+UKtX+Nn5v/dzrp33xANZf8biaIAK9n1Re
Vy9O+bphWOxTjniNDpKE3uMOI+n5702K89q39+1YP/42CEBdzpI3eUeRYnA5N/3074IRwikuuBnN
RNmRp0hRxO5MYjJr7HxHIRqK5ZSH78Vwl0tYAfO+oLm5Pkv1u1EuMnLU5lngB7vk/t/L8KJmTW8W
ouRboCl6gAzf7huGx/kEf3NSMdF0fCoX6p5BZHaXHVi0vEhdw9aqUzlk7ANn1im9KRHqCizk7GsX
4WiUPwiGpgGrwTKfSbmqhKxCVM8fuSIUZQk9PgdMP4jdguIiNM4iS21CUShoYHFiZWQlbgnBabsU
QWaQbYXHr6QQGLeDmOnSjrNtpM+/x5Yj80PHEgY3FSXCT2fg+3+lTqGH2S13quPjMfP/psc0PkkU
hdlpA/OenSGHBo9IRZXqTcxSt4TMKM7wDtOsMZHYpLBF8DS7ERYre/AZHSGjDybkuQ/p2Dwd4/Xq
ha9haFrvXtukis5ig0fl5Y7k8QwfCpTdpmjUmi2zBJbRRfYfsR/yggeiGW9z2PRG8KzPE3HxM9TI
qbdreTJdXufpX7+p8JNq1SDizqg2Tm1po8JNA7f8wBMfvRKd1WzdQXIopwCJAGYNNATtA4e2iTet
h/I2T83QPZ09NFG9R2xrdbuxyXGmdKmVqxAscV15R/bJjGCF+vt100A5MeyvQfR2hBZbWv/QR7A+
PpBh6823uv0gRJWdx2JINV9oai0F/GWA06RnFLs/GEwzFDXX1HduGVR6h3hdvVh1BKG1NK8Jxhxg
rMRui0XAG26roQpD9vlpuHfmPbp9qQiW06UjnPRrl/Bo36kB5eydt9XRFy87bi4YvLeG7Blc8Ck5
3csgmDh38hDueCuEkZ4TteH0mgwFxxOG/Rn0HVvRyO9DWISmh1zAlooUtwzzawYL2tvNNi8eUkzN
+hyh+1HjlRdxjCpeNrIsBGHF7rNt1VWXRvOU5EWPP6tNhkB+gXrrELYuDzH0/kZ0pltC48p1ofVh
XnvwHX5gFsRBwhiYLF+P8MEIcXdKW16tw+i1mrtFBhwjUa7usV5rl3Z9EP8A/lNz4OYlDjvFfEPy
kGJ5lBtTjjIPR8aRmbB5DGoVWmUqXrP4n8vbh4AyxlUbF1hcqrQ77eUTYMQpdnfT2AEGYBRIiycv
nesbisvbnQhivYnIUMs/8NiJ6YdmzuMVcROTFx54Pd96TUP1CiLH/owic3kUvI6mG/Cmk3/1+Nox
DI3Nu1n33fwPyo2XslIbgEhkbmJNhbC8cCmiwGdriToP9uAtvphaIlq+23UAbfg3zq1IWlRTGljX
G7xqh1DBBI8NiwnpNafktsO1xF3rm0VaoJNeL9AbcFp/Wg12CdBIfTO6xBG3BIi80Dg+hyXA2Vub
6z94vbBhFSRLkLfgfKnNyNJooUXmhxcenclfU+oNWl4jQooaywWxdgLBV1SDcxJVMi/mpXrFRt5r
xD2PUhhXw6JkoG7WnOJEPxFVkf7o1XuE596IO8yeq7v7rEY3tR4AaLhbp/UoypdIm+1FWkAQTkhK
JNlE8bd4A02C6tkc2nMyhqjHBs0/kFLmMcJMZ1zoMECtZiYj68WZktrglEtbdXVdpmtsjIFA5WXt
4QHm3OIwMj821c3JLVNmL2gUNr51xmGwYICwgy+JvtWwcL+iL7gOTaVrTuPNyjwixigKL6yct+9w
ozFSa7on35FKNFhcKkGm9tMkSbbMPMJduapKAzpOJidIvPG5IXIVU4JFbnoA0Ot3KqjeEt+dbLN7
rISEoN3x5D4Bx7Oef8p7jqHsCEI82CAoIlN1UT6qTcgjox9og2OFpUmJ60rc3gvGhfTF3Rnjh22x
wPXbe4FvWZX9+4rSwRjcgedZv3rP5Ks6tXDAH+HXsTjf36sEfgbqAY4aXflzEfwM29ePdcYbY4I9
08qZhWeiTaW8Rdrcx2uqmoygQPEH+M1BG528M/q1h0p4vNmDj/SWSVHzwv0lwsx5fu9ILiqE4xuj
lFOVYCrYnGzqfuFOssN7urXrssJahf+II375JyPP0VkEQeiosl3AwiTdB4zu0BojDTze3iodPpXK
//KKkPQZxxLBBEFfAMd5YLraC6SJgJWKTwuOdNCTVr9YDNXrJY4H62tMYqPivC7I8XEI9jeP31OI
cAvy8gUEciuMLTWjyry+6d6R+Oq2VF0+CjhcZ+UsKbkNehUGr9rfdJWvJ2dHbFWwIcgppWWzgQ2M
6LbLHYdTvEZt+QJiPHim9h4C/SCo4JiG3ZnAW7jDmha6qcew47OEXEsOS6nKFYAIb8qL9NzJ27JJ
+rAgfo14l1R8Ho93xEh+JDt/9XBO9ARbRV/NwXFq7Ktn+HuAfrodgOYCTSEXJJAnwassJAdS5Rto
rCOqfVbWnauGA696fhf5r/vlqEDq1Wh/IX2Y7As7pQnC1SPT8dG9Y3VY8NzEcfsT7ZsEnhBfip5k
MOPsaR61O6zu9jbgbxy+ShCRI2ee6zC0CPFEiTjmf1bOQAS2zPdj3r3lMVs1tc6bkExa+ulf/Lrk
Mum42m970bVSAHBewISpCFnvc/jt0dKU7H7rc7ywj95Jpk6FBHYbSotUhHflTM3Z0tiMW0yj+hgQ
PIZHjkiY63DiSDPQn6S4Ne18oH63RRiGhB0hVV9ky1OvojDX/UZgJ0mgugpg4rYrIkZbalzGqO82
bPT2tMCjco3B+TBaKS6d7HnuFp+yPX7bCC6rdabxAtYkM05RL8rk7t4FAMkiCc7SlN8oN344ou2p
aiSE7q+XtaUK4mBpFH+0kIVAaFkfd3KwQ+YTWuzZm5Gz9y2VqZ+6387HE8uH2dar3bwJy8bs6yO+
7k2F8ccSCf0Mg/C9HZvFlKjM5n9G/zRCB6Rd7XWwr9JnY7pP9Hzr91cJV2hnzhJomEN05oSqRDhE
4za0WCCo8BSRwNKNlnwPgfYAEqr8HLnYlrkKpZkgGdAd9yjvevDrwMkz/U0f0X+DND1VosIeYZte
T0qyr571d2wu7o1bfBea62G+Y2BF2el1aAFRAkd0xgWWLzBHrcQSAQ3VtL0LYqkB5mWEx9WoK6Q9
Hya3GxPVztFcYA22z/2Mhvzy67xsEUbR2f61KwrxLkAZGsMR5Bu2r30raR71E4cjmPAnxoQ9kS5b
ZPa0zwn70d6gSUGHP6o4UT2wSbRVWru/aUzNcQaIUPIne2XlULjjje7hB+X+k8gos1y1icGLrkhR
6V1jOT8m/PnjO6cTWC7kIBI9H+6oqAJADsrnIMaK9oCFKxDs4H1Jp0fpMLy2okBp3asWsvv1j3le
E58jBChJvu9DZBwXt6SMIFbP/ACDJ9F2zWJjsSeDcSUMu2++EW0GOxMWrNIMRQRB+zYCUJZ8os//
zKmfgRUTYcVjB5/oNgssy7Tjf/gW2zf3orgM1/Ik7FRBpIAM/q4UVcAhwSk/Vtta2F9JEI8ggjQd
+WpoLHnX6bN+lSZgfa9V13K8rAZl1x7je2Tl9ERYiAuqd8CEYq3FHoFTuM8SKQKtE9TnvzlwL4Rs
34kow0Ig+vIMo4/lfXaCalX15aW85B5xBrA5NQRL+92Wq/QX9HO2naEFghnJe8QK1H2JSC1DraRD
XNBXJt/B6g2ZO4+Ay7LeMg3SNj8WD7EdcePelkD+QI36SifVGpjR7sQYUBUbw38tYQgAUDiIm6Vi
EXTPgVGVrvSIygIhV+rWHt+ZzmPTt4vEJRleGyKX3r2xfUQz9Ifs5ScJTULDc+OOgaz5TC1qvqGX
dj71ptM+enQ6Nv7pAotN1VL9zssZhrakTTHyTRe+pS0EuqawwAdqh+nfD//Uwry2+bmGyJjlvqd3
R8fPwAS9IS5BaCuqJCkbLiMyymQKiew3vtlaVzNHrk+K8tBNt02N+eJ/L9mwhZ13eBRJyWdjtjwb
B4vsYfguTxHPh4sqZcQ0y5c1gBleokihFQnsCPOIyDzVGmpprvx5j440mSTcxuI6i9LosWxq4pMI
6ePdoMaybeT8z34o3gf1GUK7cEyBCDvDajQAoVYZB9z4t2lp/vZlUPDspvRYlf0t7XHJ1oGdj9gS
nT0G/gw+AhAHENX8ifMtM0QdLtJgn99gv6wJdlWa4hWqWZvUeGCYXK55UEVLQ1MPuwdfyThjlo8H
QsTVIhyMgXVCl+DwrVTTZWsruPFyOhAlVdlHaRsFdFHV1Hl+KEF3isdsanYeccXqO37bE/0+yOHN
pQioaDuXmokyyZPbyaHN0ewYuNaYITCRJMn66Tfosr4b0DmYmNV2ngA89cmIXyArOBqvAwu7hpWb
BJ3L04wPuT+8C+Pefk9GS2Em9i+Lb1eQtf8K3kKlM50eRjz2r2ag1zCJaB7zqkhtDtUSYCht210U
eLzAKvAv/abDyR7ajNzdY3rftfimuk1BGiPB70jIEZkDINcIPRBZ5Yqzx7s1Ejhv7bxSeVZWGbbs
MukTrgh/nO5undCfYOTqyUW6MyyYricqMa2zbfJ3qqMsH/hqByc/Lx4/HLci8ay/4PnJtHb69+I0
8S8Vn99Ln0QwYW37UYJRs8tDk0Q0CFTdhkDGUsQkNlB2d7gmMYyJmcUFnyyjd9AkytsVIqI1rn/P
Dqc8jJr/j8ge/TaTDwE0ss+b71jb3WJSvrDUciaRZTqLbx9IXbZWUyng6JeWVSGDkoLfiESq7Nle
zcrJ0gFeONu9S6rCYW4SIWY/QlyGhm4JPdp7K1gHw8uX0nqn4IGUt10VKbjtXb77+P+3lWdnxmR7
nMqzvsAP+yGuilpb8JGYC59DGzKBzyh0Wq6Lb+tv+ttOucmnGtkGzuxzlFlPOLfLzgNn1jU8h0Vm
B7fq7OYBFF1ejtaGi9oYxpyxxAt5V5s1kVtxbq7noxtu8jyJbT5PW3MZDLe7x7f9hQejrsG4DTz9
YqZM8+Snm6r4ueJhwHr9sYARdCJLTsPBW2SiobBADj/KN/fHU5ZOhsyGYohko20Gc9po5da2cZu3
p7m+xu68w9YQ1UWXXNC+Na87xIasakE7848O6qS+Tzl3ZKZDhdyuCaa6SeXpmjQTSQQeTQMmJNkX
hVWFWpd761WpIqhPVVyx8ujQRxzHyRWKj/ZFqz2axVHt2Y+n10pYLt2D25bUeAJWomvE0ajLRfdc
Mxp54SHHpFXO3NyXoF90PE23MWoW2BXoIRAWECO6UOQEDqlhOyDbMuTxg53x1Fc7qVbcxd+46l2V
s9auJ2kKEMUh/jQTA4KxMEApEPuJOgBcUcaWVfIFaglr1FIPtblRVyohoJZ1iQDuMxZDc2WCQrhH
oQgQ+B2jgGkIGzQ4YEWQG4UADFawRhHN5LRSxtEr5TLCdZJsCczE8jdbVpZO3K1vck0JNwbDle/n
Wcrbky6OxpvOanOy+e4tjD+Sl74lPX/OZ5WPlwRy7dU3gwv5A44nR1xvZqGNNVqm+5qRo5eTXIGT
wEc+NRiHRXf2Zr5oUqqEsRcGExV0eZZ+7dqOvxDjqSLjZLWLqQM4FoDFLnqzLfhAg2zYFO9af1Ag
VanflWCsUBS5o//5Qq1js1e/ewtOb3Dcc69/XRN1PSw41YHHc+MggsFW44LvDPcdPnLZrJ9tWv22
AmrHQ4MwqCCnK5PDAijraeZNmEVf8snMCUCnvJUw/k3nyiEP4uzukd82Ni0V1A3F/t3OEidPaHXS
8HjXj3QEFMVhuNKhLjhkyaSoUy5xJuUZKDT6cycbW67y0XFSbid3OuDooL9cXaRK7yGwMp+vCGN/
mTF+vcBiAvvUntZIIlOXtd2/d0Dj3tlxhOAgtMvo08hd8BUYgewt196nlJ01GZGpNXF/vm89QTj7
6liB1cUMN5mO7EYMOQbGTgBrV5WoEC8onl2/EvMmLRcfsXjrJon3EE6B2FHVTFP+MndxaaqhjQh8
ThDejCtPYfV2f1uQ8lETY681Xxs5ZtPm24YGJZGUXf7tUIhsnRngdCypAVPI2HtfPzXLQjHhb2zz
buGLiQJckULGnrcPqPP4f8Bgu35UcyWGwDNRB/R5ybOJ4uNKXfqUbhtgVDRBQFmC008Su5WKUmZS
Jlq18xQyOaD6SXvMV0lpDK5CqwX8EkaDDqZDPFxZleaJAnb0CZqYzSqEZXUv0llDcQVVmjpv8m1N
l4UcegF5gMLOIzxmLNRZVyg1AugLpMGbp//eJyeFJxf9EzsBvn+4hYe5/CYYiwaCmgY6AiS242VD
+ciPBkoK1nAVh35h9A+0skeojVPPVIYRQAexQpgsI5f++u6JbXe4qDbrZ+llSGjHKXy8ffgPxtMf
eg3wnAwGPPUiCRP6vZxbwv0bmF4H98JH8sKqv2FA+o6TDOasWgsE3nxizcEZAVh02mrv7yPtCoFX
pdhaQLv+vkwsBNI5PQZvRi0lE1H+EOGYC3qD+AG5lip5wQVg0BT9IxLItCXQwkAqEjKl01fS576j
NOKdVIEyTyXyYeroV8ZkQA799HOGaMCyfjPMEIkKQNlHtJGxDljzIvq5bzS2uFzCqTJLRT+GJodl
+48GUsWh/iR25knxPKv0d54ivznU9omABglnddWXtkgofUpNr0zGThN75dU9q6ZItvlrn8nhhsfG
y+TBpG7cpkqZj22xi3Vl69PA7GaqRsEPIxJye6/ZkAzQEebHARU1Y+hl6QzRaaKisV4oeIUEQ3NK
1vc9tsFuOOoBv7yIx41gglcjVMRyKGCNgjh4yUdg3N1o6INdMofMnyx/voYEw8IHUoQSfPzzeQUN
zdTVPl0aJpYiKpFvehQvdsMTkPXiotfyJw5wQyNy9EMHcxcZ24Gp+DEFa6U8J1MT/F88dFoQL0Ex
WxQ0Yl12C1uQwIATgduBHEbJMySEMMvI3pf/1jJhCg2PbMKmEJsiZRQJib3wn8UxUmox8D/6/gkN
uFiLv4dE5dx2LJSyWZm/LGeK7gCe6XUWH/DL+Mgxu/sqnqspZE6NEs/YTsqyiP65B78qGEHMXe/d
n1G+AO1HKWEEEYHvP+jqABR90IOAh53IDjKS7/51oyqBDSEkxHt4zvVd5iIBUZ0JF0Esj13C0NPS
pTgw40Qs0mmdZAe/QMhY4zilormdPRZJy+yiL/+1PMpw2k9FsjLZ5gimD2cb3nu2jXoEKg8/AFzn
1sNoLCZmVBygV9WFtItwRoJjde8o/uXruo/+Adc8CXl2+X5CWwOJQ/NxUD/P53xVOzjcqeYi/Kbg
+FgTqzIPHw1lhgYwSs3xChvQ73CKEsqvrl3zBppujWxsCm0OjCB504AhucGMth2rRpKpSk0nz5FX
ti35J52liFRTtEb6INnDuWyZNcAPisgpIRGqrmcY128vVaj62c6LjdOoAyrpc8iBGnIaVYJS3Mn0
iWF0TEMz01cQ4M5L1oVHoj6GFGKuWDDBtYVMdipgiRDkM2TZQRIil2eUQFikRaNDr+F56meOQkqh
e5uGva5aOp7Dh6Bc1nUhSG77/v2GH+G5V8cBxSxofAXaeD/EB10WDDcdN1LdTLTwMfhKtFqXu0uS
Dd5h/UwyZaJvWMT/zGqOMVt4TUjIdmkVU/6wVUBITzLX50s06gTojete48Oubpr2SViZeR2X5734
2fDGVFriTjPdPHwhOsr5dlZlkKtJATCzC8lTC/DH8W0tDbtzsEWZkQ+2c5sJdkc4YuKYJwu2a00+
2F8mro8KjjdFOX1Ylfd1g+DuLEcaFofIQnHegMI0uYo02VjmSmNvUPMBETClmLRJgQMl5NeNZg8k
r9ay4upCuM/9iWwtzHbcKpnNf74J6KKbY8tYFGLosphRyAcKFbSSXFtswQNKy7Xsmw82SOONMWqC
Q0WBN48DZHJld6WoYqi6LjIaDWvigli97VAvBv3pacxT9+jUtcx0w6cwRjPTk+3fIHvZwqjEdVbP
ghgcygM3NYhvUheZre+OgNCtvHv1EtRc9IeIVecpHrH1sYhCkqTeSQLo4iivkG8fUI+c2OnMwuAh
hNZ3LLYLvbZlzTHZKlAsA+afCNMHKAsdU5oMMKCE63XumUfpZC4FPmdzUDYzjFYkLX+pf2uL8Lvl
8bgdlX9SQGBxhAm5771wBvJxh6cYHQP4pQPKP0xZFruyas5uF457r6ek0RSfY6Xv1gtPs1TaOUKV
DgE/wibY/n5rBjlt/azXHcGJX2IjPsZgGVhWO7SN8X0rUcKZZawhfYTjprbiXfzytOx2HkKF6c+P
h+kTtQeQHB4+g8A+8elwlOtCQlToGdRj0ypioT4QjncRyP1GpUFoja4GZomLkc6QtGLaVtebKFJI
CgOzB5Tl7Vx2YVs0XJ6z7y4jKWn+vark7Q9oHJdFLwQUwB4lrZvrvTsPh3vbnqG/j1os7PED5krD
bKM7Hs70dMop6sA8y8bS343dqx7zqOvn28eems7FdkbriSRjyZXUAOc10wfl5TPluEYxnYdvhg94
WMJyXL/SDoo07jz50yRuMVaeTEb8DLeNskhy6jSj83yTR+p03+tH+mF05VzTWYOb26usliDZlvDG
WCOV/UGESDZ8AboOaGJ6TwdRfV9bShgNZo3CHPDlCHawF5S0v+y1uABlhEs5bpHUzJqjd5UqEMTm
64G1NeT1csogF1NOsN346w+23spiatFmvLXWHy8TrmGRE/THFyd/0/geHjo2ZKTQujb4lPlf7Btx
ekL09suvZIwaBKCFj/U5zhd3xeDOP+x9PYpbpWLx/9SpnpvM2AGBQHrD2Kob1XPG9CVz6Y6PkDOv
Bu9LqdLN+61q+KtfmlbssDpsvN+v1ZirPoEJ8XxfgW+d7aLbNVl3t0bdtX427L/3Vxyr0S5p9uVC
hgIK++d175Gupu/7bllc6absXmwxZLrv/raqtPbDFFGMyF3LGLmgfcqJPCsBw70qlpe8uMJMQ+Wc
+a+YGmgE8U4htsmxrV33johy+O//6Xs9nHSFphLXJWNFt2k3+EIghyto0uYiLxg2BrBjrZNZv5o7
sKJRZzzAYpsjSiPn/2Pxvpm9qMjTpqnFv35V7Ub30quIzgSQFZwPFwxuQKs4OG9QwZSezNBuI2UB
ImnDYPfU00NHePqwL2SI3DRs+8QwxdGd0VqvsJcr4XZSVK7fcCYucDLtI8RkXb2HDr02KP1iS4KA
9xby50tjwnkQxEbgyIHsz+mO2kLcvzgc7OyWzI48prI3GRa2YSy7JzRSiCVcmSZm0+Nnavp4AwfL
vFuO65rmgLJlN1p3juNnRVQnSVGanGO6V2alWA6xGtDvfbD2BvKqvduoT6EGntfO+lI/sPCMoO/m
29TgWbkUPSXZtdppTVD6gtpSqS27gYlcXJdMNIGAt9n4MIYck8TJzpw+RENxpG3mKGCXh0jBkaFy
FofWyEBYN87xc7X8ozGr7CrxDsL0Xswi9rKxcE5K2Ov0ip9gIGod1noWkCh9U8EM4rt7s9XXB9wg
kg3CE+bo2YF8k23xJcZRcZgwoU1m3ipOQ2blh2BNHMdBRweV/wEXowj/Z2HoW0yh6+M4THFYjtl6
ZRbiGDERrxGNygS5oQDnu/4wV3zJbpaPTCMejMf9kcUUXnGkbU8A4w2sWaLVp7Aok+Q3kuoIY/+B
T5bAnGa8o+SF31/X7iIchNubY0D3i1SJNqE21PUCDYq6e+3zh2FKNtNhNjbTQxHhWsp58TyROxzt
Yh+xS+RaMuJYEYDVZfa5UPpOKXT16xGKoj1YYRujoFt2S/h3n2URE2gUk1mYBnrfUSP/1cpvls6A
/ia5C1NCAmyxiM+pVpfdIjRuSwFLnltT7TD7QwQHRrXxi5e1caRf73k0u1aHsLti/vmYsGbVD7/t
GXZlvnyZfAONdSWeKuXhO4yFgka+KSdG+kTiFeCdMxoAVsKQvCQgk/+5LSYMEYPPsY2FJc157CaG
zkjkBD/GGe7FgWpJ/33VCC045GntSARXayUAOXdB37548oZLLlfsvM4zor8CJvAwkurWt3FeDtLZ
Tk6koslFKPKWIGn3RXb09Sk5jM2imZe8+nTUUl8mQt+7BBy4Z7ylrYNigX2BKaHP2zoT0DUWBpip
wlygawmqE8SWB8GAXyK38KYnlVclt7P44nlA0N4iQf+oegfDWIQmy8V4upn5bjsZWYNSzddPkZc6
didgMOe15ONuxcA1mK/Vb8cUNRpJFKMP1jS5RPkxXai6VqRP4x/7q4HQXGA8rOSYq91D79StnaGJ
r1CgvO4ULCqy/rw7hiBvHPGw4G3PBRwDwNub0yy3QJ9OpuGFxaNuklppsb1ZVJf3EC3CV2iDStb2
a7+wC6Pd3b37dQdU0njtsMkp7nqsHxj3maYjmi4s3IKqCNOA59QM+DnB9xo3EdQ85QUuo8VMGVMF
EHBiHe18XLhmjhntj/q1duKfbBzz3ALJXJ3lpts1pWnh4V2KhhMx1TCWVK8Uhh73eG9bY09Y0VxX
xpzh2HUM+fOZ01F4Dfj53s6JhwEeaH8lGfPuWp7+rtwstnwiCiU4HmGBvHcYtG9gF47+GFYaxjTt
1D+UL9Zbeem7VXyPYRio1yFQo6fg4Q4fwddswW16dwd/CvRIDOyArsQZgLfIfobgKRV2VXs4Gc8g
3JD4sFIsI3RQVnA3qGuHbWGp0GMK+BeuYakIm2seoQtkPFl4RfOG4dGPD7bHwegqckgIDdw72mVY
XVYUWJ76X5OfK19ysX3o/3BZm/vwbkD3EEy+eeUy/NpRIKBXZLOkO6FGDP/fTd50dEf7cO7QkNrS
vvDJw3RqBkEtHe+S/pdMndes6W8o7rjJYZ/OeRdF0FqZaxNJ7oBeJRbQPOCJtGXbFSPj1K2lci4g
RYTSBCCd4jMjdwFcXasKATFSkRuqxgQxcm3EctnAT/QrDP5ted9sTb96gkuWMHgUnZvzxacFwC5g
K3ZwUYRPPLQ8xSID9EstUHQbkMZ8TwxJxSHOo+QObqIovxhNUPw/VlJrr/HQVm5b1vGT2Ao3DLqD
at0PDuSb6rHwDqWQ14qiQQGn1ezgdmsR8MfzH0jvEn6HAWvs1Vu/3rTJHRmNv8reSIKas4FQc71p
Hz7DLbv6kgWp+onPjYfauuZH7RBJuXSDq9wSQVxnknwC56AmqvzNnyjYrpJ0IYcWEBDZEsWVQB+h
83nhnDsAw/yysfnNmxfEIEjGx023g4CSsf8bN3fyS0V/QvKjoeXHORYRzpijyi7Z9mRSi+XOMbyO
ae0gYxegu9HbDoD9kzD8J5y1wkGFGctHw5teak0SMt4W08BygRv9Cy/Lf/SHMkmGA1Oa4Hb2KdQQ
gm4r7nPwUqgEOusX6/BObsDT+Xntzj3ZMtUQAAILufmRoeCz3DENTmvmCBaWvU4wMLz9i0oB4ZHS
NmqiN27xlVN/jgmcXmDil/eo15r7T1kNUwfA+jJaS2NHxfsIIroLABbji4DgbyMx+BbQc7vyk/50
caO7ckl2D9IHs84/+u5l7ZyMb/jVjA3FZgUXf8qhZiu6WN8l0khsxXrF5ZU6BD+jgGz62FBk+LXN
TirmNWzLycqIrMXLP8CxCc899a8sVWuA7C0jv938bOLAoFoF8mpsGkLjNPOIe/JK5ZSuwMO659EY
h+koBMEX00JSAnlNO7WsZF+HC5YS7ofspJYVr9DDsZcXm3e1+vek0SwWEHuE3VhEhRDrmKEnQhC1
a3J4d0V+yYWtpm2h7oKxxFBaJ0QOVxoZ/9z64qwQws5T5VX871rymH8pj1If+vnuJL2faf3hA+ue
g3MTWt+31IDKfg+nKjEegExIFPa57c2438yjpKeDlXaqzCV3iLkN+vm1nfbYrUoA6nh4R8kHe91I
mfIjs+917y4g5E1oBH9nTQzc9IP+AivGZoQcNBDEkYdf/ElRqu6zwFqC2+nEO2DHxH1ZjnBKKCif
CGkrFfVBRFTL+oupzq4pGS+mbx4iT3VEKd8oXsEnXPwYXVyWbedYew024pKQZa3uUYD/4bYc2O8x
WGbbsviZLocAoOT03UgBBS4kWrbLFoVqBvqIqpdF62oApDiioC+ySdRS6s1coUBR00OV/X1QDwtu
tzjXoj9AmElqsgIeXCFoskM5EfriXQ98Cxu2uX/RmmiwvBQ9zuxBZhOZq6naxtowckXcvd+m7SVw
lcThs5rHZhpvG4PqLwqmteECXduqbl8yiAm/WN6hSBwIQLiwZ/6gzfUdnOMbu9lmd4SbFH7PKqxx
0SewFnPAQqMs3cncUW7jB2jS9GUMj3RqugeztbkavAaJGDblkkH5UXPlNancMRMFEDsqTP296YSv
EtWurU+3mSHWwJwvkBfJuG4ZdkYV07E3u6x5ZLXQM7Y6uUik8EFEEb2Kdr6ogqRxVAO0577XtJq1
Rkn4UIDasCPPeR7hmj3HmMtDqVarYYTvN7p1tBKKoMsTGHMVu32rgFIzSJ7zGqj1K+6WDQWJXgH0
IfXjosfDvUVUdAcprc8/4IPj5UsG4Kb4WYjQS+BCYc7nQBiNGFoqC5dqW7d6kc4omQu+u1may50I
F0gtvW4XZ8ZU8ziS58DrWf7nivFa0Fe6U2XBsJC9zYedhcvq1XkPmsCuo69u4x/rxQqPjxcCEPo3
aFXzfOJVpXUuLbghzPyDbEbPWvbUs3dJRCx1ESQGJP+99Tg/4Uh1pQnJYb1RRR08f2fEEDjsaxcf
hXSvZJsXZmlyqV4QCPDePcYo8srB4PVumb6uqjx8ZYUdydrWeNyKDzmjUx3AUSl0iD8uVCpsovSq
ENf7CZCru7jjHl/W+L/RpypDVxUoMrgRBve40NbG+ZNwxeDiPq3kG0JT+g9os974g3kyskja45i4
Uh7I5AsCmMfZjeDmParKekJVC23JAB9YSHU2ZsiGUwUG403OiLrgBdpB4gMGX+RZn3FfXt7ruasN
JkCKf0tSdkQlhZIuhsPuhIcNSQBCde+Dn2YnXiFDHnNVVNsfCowk+bigUCeXPG7AvWj6gL4ztbSH
VNmNHyrCBGWfEI8kl+mO/0lMeZA26YZOLdyvTtVACFBwsu2Ug4qM+HpNtg+5+6SY6/gRXX0mMHX+
5HQb4lUwyd0iFiq0LKk3kOsVpnTyyS80Yip1W5/7LTD5phNH+Ey7pxeO1CWMAjU6jtecrAE1kI/c
Hky4ATf6MXVZ36beyovqnYVtPxOAMmaUigqZtl+NcaJdfg/9AGkM2IhJZ8TwuYs+QiuiiWs/V4B3
aTV+4cs87rmW4S0zYK4gSTyTdm5S+ygk2aALcY2paD3msAApuJkWQ/5rrP1LDjwZCOWryfv+V7eO
ZROzsR0xGJVAVz73VHB0JW8BG913T3tp3CrKl/zEhSZZT5ygwZwN5dyXZp4xUKphj9RiXGAqgUnH
HoYSpVFnxGeQjsYjyVMDTtcReo/XG0CIjwgUhbaNI7155CotEFQpiW3WQn35IW2KHWjLNZAYkmbM
SJssjB+9NkbkeQaP7sBW8KtZOe/Cq0LXhGPX24qyegbsqyvH8S3MztKlUkUEserRvzySxFIkKXDe
ye3GhoREEuXNSj8Rg4CX3smEl/wI+QOPBFW+2xBfsD5tZy6vIaJtztp7ZgM/lqs0S3huCcBr0TFa
6x3PStPfxwioeqoP0OemZhmwcyNvED1/KrOZGqu3KY0VeyXJcePwS7+bqc0Y/+sYMqxW91vO2yDO
b6YtPYz6W/WVbbhUVd8Tdai8EsOoHl+G3BR70TtkiYm9TaQLbQz2ONL0Xn1tEMgCZzXtEtQZGHpY
pf9R4cJXN/Z5UJpX/Sgnd593JHhJP4Uu0yKQRHMAFUf0dXYkJoUuF0ECFXzcOQhtGsPBqjMhVPX6
6KHWqUALPKXhIn3HeNfgVYihFHHDn6rUlSpy6/EmTDY/OJd1R3dhbBE5TIuwS0aaqr63ufq8PEbD
2VYNuog7FF6tx1BogUi0iQ/HSVQ7i4ZEVZMQuVl1qLfKgxaftnSwFvxJV+ywQ6uTuYAYxPZSrlOw
I398OOGvzj0bQst/fP6Wg7jwpFebMApIGH26fO+ugiePLunZyZ/7T/N0yEL3p/kR0hPmJ5jLC4vi
l/voYsIhw6zZTudogEBAxzuu3bwuuRznworMEdIY6Miei5HcArtBRcX32MwfrhBCc8zufX9h3bpM
9MwzL71gcAyoBy3R7moVS1jQSZWadn1EwcQSDxHNjSM0MMMKrIu0pPR69Fny9VOg+apRgnyEaPVI
OA5m1YsCjk1movqF8D74i7CmSie4ZSP9lbIeux+O+KqURvjolRzATZf7/TShym6+cLhXaR5wfXV5
WTtKIIgmsMmjBywWx7SPyjSDoCp+qbkL039u6FegWTEISLLCtPIGpZxjUvRciPy138POwIoYm68i
bQIYuczJOnTDNrDiC5NtgDIVThmU6fQuXZ6YqZkSeeWopZ8UBfVtYKWQ93+WsDIiciYaIi7rdP3N
ONsN7NU5c8leL4PQUf9Ygem49nVVv+FKD91JU6o0ZDCOCdszc9xYVz9bykSWsF8z8xQG5XSNZzCS
JsuZqGGswlFsitipf9GiG/LR/KgrBrrTCObAXifedpKerA161FW6IycfKtdjiacao9eZ9ftedlct
AnJNS9Upl5MQtUq6e+CBxGrrMWNlSpV4HOTIcIWBRMGRGZcjl+pVburhxJNqwja/5fmSOTB4uh7U
XL4GgyvRmKJ5J2+2uPK9X/GzC7NiVKIMTyqwYV+p3Bg61UchNhuwWwF3LPFeZa8aNxl6mOSl1+fa
dU1kUyQlH+ExPnjI6xOYTa8erzOfIqw7zHfJ0pVt7eEry80jFkqYNdV3rJuVb8J50EyAcvmb5y63
oEGWIC11iAZ1J9YDfAcMMv/Y1HuTBWu7a0mpi3JRd5dY+TTB6vzBzh54Al2K96BRumWB6MCbYs9o
uqwDp1GxGghxxVGcvhFE4gg2ZD+UdpBPUTkn86e00T0FOFutOTkKgHrZdwIXTAs1TM+L3i/21HBu
4lO5n7mcaBvK+M8HoFZVf5B09JqcYDcvY03ugS0rFyfBaGOeHq4nuAJEPz2JZgFQZ05ALZsSZdVC
yRdtJ0lHc6oUblUUDouCi212ssE9aafsbgsxCeX0ZZkjJOTQ8tLGMB5JtoHYEr5XvabFSzZW4Qnv
Oxpy1ZHnxGYyJiQTo/knBLTo8gNtjs7cpeU6mmmn9TvvX+kU5Efy7CEujCDxFozA3KhE/hG7q7I9
/iPP9M/RY9F9jLYXpWkraeqfncQvG+5vuyeXgggGlveZOhB9zCziuuGY3z/qSUx/51kK0TNSIVjD
LSBzLi2hGIlriI+gD5mfLOnuY1pZueoMuUj1dA0tzZQydQEFcteGKH57WyFrgtHXNPBJZskNDC3K
s3wYOgA+CVmyMDa+2wWII0cZNK/CWoKmB8s8uRwGTXIiTgUdL37fhyj3Sn937qxDnvs5wyknv/58
Wx+RKNRXkSVHh9x6/rJH8ydj3mJkvOsHRP1YKt8oBKiCSMTRL2SUN0sEtIpMaQhAJDE8BVoTeiOC
rZQAMymXx1S1xQAqZqRTkvlcem59ToKGkhlUy+TTpPFdqF5LReZc9YJfQIalkpIIperRjZdBaO2k
JKOq3C2Q4Gh4PZkgWf6gT9yMI13zZaWh6OadWFEYbWT5Kf1BFShH7/P1navDWUPArcT69FJlm9u+
Y/sXegCFydoffdaGS+ZjXy/Edi0j0+VNv5I7pdYdcg9GyXMxids17/oZt+juRUHkkB80J+EKYCLS
zsn92P9g2iyYNoVp7BLDsmrDXjosCyk8woH6h5BeoE2ENyYu8S1RwiFtWFGe4a5qXTtfg7WSF515
poQJhXbT0IoWTW2Jq9KkW/uFHUyv2eQs7fY1AFWrKloZpCtV4nhd+3YbHU8qZV3Hk/mC9/gBf0sK
hHQ8RqPFVy3fn8l8pRXNP5xhvz2xDGMLX76UqQKoxpKVydyVl2tcfKMTUm2lywLaIvAo8ictQ05Y
lVINPScxT/LrGUs47kW4Rarl9wXOtRkzwB7+yR2VjmDWaxY/KPjjGjKGP3u3wQLysJbV8dlBc6F7
T24rEcIvdqWOjf/wKVHc7wlL+GViaDX9X17xZKA7M48xjrdCKieAix8OqevQfm4GCyCMRlDMEU7d
lmbV1gFHrswhmkfah76vGeGgo12+UpEicYpnMk+wP76fNLSZv1AyfNBIMtw9zip7VYkFylvHyorl
vqanfJFMvExd+16WI6grLii1hW8xrnxoWHlqSIDhpowkAQmXLhvPj1ogwQzxUqdWkQCqkUGiSOMZ
6uygXi7sqWJiG6SQzrsc90fznq5s9FLGcqDMKIzIYfV/Az26tlGVMonfQp28mks2miU5fDJ1p0NE
BvkMarOrjwLUfVNY/A+SId9TvQ32K4FiBQplSji0wSB3kyfmgojBNDKa2edBSxf/M2yw43fGcy0I
JbR9fdzXA4qZOOVDuelawbfPZzSJIHUSPqLY3l89/nbWBmZtuM2fKxo1KwWYdIrJGdw9nb5fzsEk
CdRAtEuphpYiXLc2Jfccvc1RiHvyzTrzNXFejwzY339vdiPMblWTtYXKrfQSb+hGtFBrWIDNkMXA
Q5PkA3WsmJ2m+8RF7lzP8zo8P9pPAG2MEi1Ltg++0huKcT/KrU6lSTofSvbAKKG0kyDQHxbJEnAw
jXg/Aulb391Xt3KXqmhNydG2gdVH+aJi5hzaKIweg6wQLffCBdJ7324Af8FAps0qw/eaocosXYWK
+19F6plGFVBH82WHMzU3OU49APHEvtW3XfwLsHt9eEI2KMkTXwfHzvsz+ERlkOw30YJg9xHYy+TY
3UsmOHobk6BRQ7+RoIEhAEQclVPi7lQ3qiyrtwLqE8mfwxFNeiSAO/mXrscsWk+lPJ6z5/XNp+b5
9TNqnPTwn/p8AWJzS2tCEpooKLXV3oXpFlv5//kn8KogxIZg1lF8HiycdkPiDjZlzZTKheyFUVK1
2Pw7pSuceAwL6HG9FWxoSwjjI9eB/AJJCBm3Xc0HzZxVKoEhpmIKIRiUOQdzCyG6GcgoqDHj3ROS
LwwzNfcpOwsCsh5FsMtaIC6DG/KrBNzZ0JbCQxXSepjoHv38til41mUnYSqUyZkMaVEEHZcmBNDm
dv1jShtpF22DXuz0En8kl1O2Uw1GrIFjhdB8AaBeW+Ki40NLYXMCyxUuuskTZoUkNJ0hEjkO3H2E
06vKNOOT4LtYXyyzdnrIbVushRsVdgp6mCpSco5UnVNju5fPMGj8oMHuvaYpofkOt2uZc8jFU+oI
p5DVPxBqoenxStXPUAo/M08H1afqZGn5Nz5gHJ6XZowDOrR2LyRUrFtX+Szdnrzm/XJPkwuURJAu
e5y8qi8H+FX18Xsdki9WfqnI/cZkOA7leUVfo/JZfFgBaAVdnLiGrFQTLi31/Sl6KcatA4tJiUFJ
bNUi3sdj5aDKuBQxYgblZ70G61/uxh5dxdhcZw8+iYGcXU6nAb4GpkNzKEt6cly5wWQMd6A6uMda
yv0XpwOJZBfYL4M4LFft12ge3nG5/7bIOTRUQWMhC3BVEcUnxeI4Zw4BhESigytf0WlZ/u+JXceB
98YErovgfrcvL4XiRx6ZkimokHOioiRkA3H5O7RXaDrCh7JQdlt+hnAant3tRnC6GPBaDx2VddsD
6waa23cM94Va0ZN9pCWrFBQDhvRys4acVmG4tXnagz5Ttm7DUR3Bj8QnzuJecdQ/VhKTJkxcMWo+
F9CdUPgR5N9O8uiA8yb5fLizHQLZqubvh86PCJvQy6qHA9x4ZQ4xts7EldAZSz/kZuUY35SEnkmn
pm7XFMMuFXLKAZPGrRI/NDZ4N2y35tn3EFbsJtFUXTmZzbS0/yQDJlQ1j0fK7IbUhmx8Dxb6R1KT
b0AnpszfW28wIIr4/0eyfi+4J22I4A4hkJWLSOh5/zPG5ZsSH8WYQgcW8yLChvFKOoTLY/AY7sj+
hdyV0t79sThPYfrVTd75RRej3KBs8c+VMsZ0l9Bnb2Lj2IT6fyAHFb8iSXNa9REEgAJ8C3A640oM
eufjUBn3RlMpj5JsumkVsrNfe7bwtWKQXu+2GqVyrI9iWGHPox1r0O3n7SLg93SqU4MIkd7p6S/L
/RLyWp6skMs0M29cJvEzcf1NpTjyI4SXg+d4G3jEwd8YXkaAcL+EZOxYkXDykZl44lyFnSjGBrke
0tUukSlajKs0c9JQd81Q6z6HUXPY7Yz79bjGIdZQj4lKNsD6CXPaFmVLxMkFSxlgWYVhhyuW7X2H
ig3w10tYD89+oBFJWvCXYLbMZ5+tly4umd681XEzNbN0nLv4svxbI4uc8nUAWvLa3zSyIiTKS6iI
2gs6ko02+M1E+RmKDH9KDwrAZjr4dF9jcP45hIKUYHxbsjks38Jc0xI947RpfOcaBdJASrTSpKtv
ypUKriEYpT4Cg9WUEdgU64HOOvYqTgOJ+sokT2Axzs8nAOe47brQ5pU8vsnrfmcgivDy3Zz5Sufn
t/App+kHRAC6OThbORKfXiKa17Z4iVPi58oaUsO7iWikndJLUIFmrq1TsNNQIOO3IUhStEaXSnLx
6WooHZukJoJ9AR4zn+TRRXMymqH8gO/6/sTzEY8AEPVoYWjDZv1JdQhICXoJok8q8h9Uhze3c/Gn
QSfNDd5RZej0ZQYfrhTXBg0nutG4iaPW+DgnHIREmZUUBH7LEVQZIFmN1biCifwZ7drayKzi4ITm
ycN6MChYFQYqbE0dXBaZduuoe/lK7rPlRyhVlSqePEQjClC9gkLqSn6vIGMJJbcp6JBevSpxb9UT
5M7Cgc97LsS8+s7qswbJ7Lv5YKYR3fYuy9/7LwWjGRJqFvhrUXrb+Z6iRtLZlpkFzINIEW+wFIL/
+0JNfOt4ZPhIK5fjrQaIZu28YUhHAB0GZtI+fNQyIXSxGES/vTiYdiDKquYep3gaT5VGvO5E9ylH
8lIU6aVlMIb2444cLnqiYZb1JEG2z/M/XmM54Esyna8F0n5ufnBqUy0/bAkmSU8ZCW/JPBC3SCqN
kYU3ftKNVXktoEEZcB6iVFDlDJ6tW3fWsXvhFYUIvOy6MOAMesImEgkNkewqDdTn67wpzl+X7Tnn
TD/zOrEVWYNvqbtKVdHV2/dvByneHAOn/sv1h4SGptqKWV+OEgGffnHAv5JEcHmtD9o/eUHkQu+2
9Tmgma4RToKqmfEIqvz6cH1tsdvcPgN9deivOgmQaGgc0QdpkB0S7i1tOtCPytQe3Sm5jJC+aw6D
LSZDuNksgC3dZBgIcnw7vcW5CGVBwTnp9oXGRE/u7rjodFLGrCMGJUHagIyI6KbIjuArF7io/8BX
f37yi3Lv7AnKP6B9EKx33n5yRREpegcFUY4loz+gd3SJdccvSD5HmZwUlUdKFJFv9Gu7l9MhR8rf
odSd4tuFFUPyEU2Ddcp17z7DpB658nVt4En1rIWJIdPRMb2xfMdIAqO/OnKxYw3IJJNHMaCqoHgj
8yRd/wEYz2MAd5jENNERwHYoMgYUXIyGo444/kq5/y+UoB5IpXb2DEU0CDlwlkx9yPZA8s6N4Z6Q
i1ZfXieqW5QFv9IttiYh+3Z0QhC5BghwYr03OXbbkIdBtZ19535tgubc+YxOLa5INF3KJz+IHrAA
5Mywn/tFCIIBDYje5055wKq3yd1HQrc3QSNYaUyAR2t6fr8tYJm5ffiXPrr9fgMwPuBQNDqnOi8e
FK+KmaOZCDhgBOSuLrJqNG/swg4b0eI9gxTZR01XOTse+HeHgE9NEZWENJOlwF2qfQRe36pslRyV
daW/XIP8k04t0YslYFNrOixFjA2Dq8Y8+NKz5TsiB2W/xny0HIiV+htJKSibdfoqILgFJUga7GLD
vKcBYejugFYZw/Ir0r0OeloVuk1Jf3T2QRoKETmfuPslRubQrhtzu+2ZyDGo2om7Q13xTN0q2PYa
k5OzLAYpkZM09JYloE/iDes1c3AOY8E4B8lYRWIeEcSj3SpczMe0wdS+5HsLJ0FQ6Qfqy4MTsZy7
S/7mxHyj9G58XooEUWryhyECWj09WkB1JA1zXwW6OLW8xa4WzYV2iy904ro8cc1vwtCnUuBvVcM3
jHrUDu71oT9aQtw8RK/gUMIi/P6jU+82J3OGVpT4pVRpnv2FTLAm6r1UXWQ7IQs4Wm4H6ShPJM4F
P04gwOX7BwqBY2toEskqvwMzoaSh46RaqvDQs1aajHy7VJ3+CerlxSC56bK8/zY5JLXapm6ryIT9
eoHGx/4mhwKVPtt+8HcyfZTRzme+fPtuYRwL/znTN7gQUUO1E1oRGbhrSTG01OGQP76MYijM/UIY
8u4glPGMA1SDIsMcVv0auHmWOh57sJqcIRMnQ0cczYJ2T0dC0tvXd13Zxm69lKlyQuqoFTDaJ1cf
CamxAWhMtGUv4SuNOWh+r4yfLM8h5R9w06fxTD4JQ0qwO9vAWPfl9b0wVET9Tni+CX5agibkCjy2
AGOAxaHswXhk4HKj3Z2Jkj4/oYKiyE/tfjmoih643mfAEXDtz9qXSxjLVqr8uTW3Od1mJHILPVs4
3sKQ/IYKkTp1sP2hKqjiGuoI1kkV9t8kXA1+ljYpjW+XGfj/yoOhdRT3XlwgwNGyi1HVYgWiKMbl
aQgagTKa6XsyIKWevIjh0FYE9fP9MYJsdIt6tjLTB9ftovGyFGvdnElx2FZFegxpONXe74iACq7D
rNAeQisq6c8VBYoXeSa6VIE2P8+nwktvwfL71J4fkfHrK920WHfI+wErrspy+JIyKYbfjjdpXchw
70WRhAgifhJzZuPp8ApX5+l3gfJPu+CdQss0pbQj5GSaiWKYHQaR0IxswIx0Vko38z577o+5M2NL
dkpwHbhwC8WMf+bAGrZP+GSVligrrP1H7k/zSp1q7iG/tgxjPf39DOY8ZGKZnDcDjX5/qaYbixq8
QYtBj+tGlwNBzHNuyU8kUSV9+zXKb0USiMB9JYZZVvNE0YOd3RsysIpeDIK7PPqHrP+I6ngi7QT6
NfZSneu1zif12eBy5KnB8cWPR8SAaKM0ao2fg6BGLoFs1Ou3koYkIlIylSjd6V8vwLt/8dMTkb3B
QVKrIRNz4N7cJpS57MbDO1vGHaszUDj+8CRTi2PhfWdP7t44ZrVMSlnsk6XbxCAWV4C3xaD3T98o
bdUEmEyEOnpedJBxfG/R7684DDPD7e5TyeqoQ1ppg6C0R1SCrLRnDXocyyOxNo45lc8DwDkpADAg
D3iFIGkXqYo+gBziatrlQOlXztAutiSoxm/sNDOGI3BC3OOh/d5osDNXNYQCdC7qOnQ0wFDN3L99
4kFIexcVl8WYkO9HKTvGy+yL1JRRvs42/hz1k1crz0eIG3Qa/LSnnZgWUDIrhg/xYMDKZzm8SpZw
awGkvgYn0IT1WOhcgyuzF09U5CPWJVtfCw1CAaZXx+iaC+3SYXSO3v1+smnsRqnHT5sebti2Aqo7
y6kLpLC8gLTywIyQwSXG0Cn+RZvoShZpZ5k7SsVPdRBuC100Lbi6Dhmz+iZ5R1BPDn9SNCb+YAld
82vi7B/QwpCo6nz/WFMlhIQdKqMINCCzeuWI1ok9O3LlV3rJbOFnbUgrNumDNEJTA7HCo7eA+Gl9
6YPKhY8AOPIXg+M+rG2tWCZ01fUXWDcTEEfFpFW1t7/hG+/elDmpb4JiCQySrvZurkS6ZKEoqnVQ
o7u2hB+9Qa6VxfomF0vxo7Nx5cqy5gOKWHGOevKkyMJvnfc+T4/pNKGRso/QSKunZCjBz+5xMrrG
dJJUFPeRXbp0v1X9Ye4Jm8ZzaXCotiybfQqJF/xCUKwcmxJg5XRiCfftVn3JsmqtEes7L6NO6vo7
FLDODrLC+lJPQYUDwIHr55LHuKFcaG56XUzsR0ALfC1esCnGDiX9UASo8r953HTOgtnQpJHJmC18
dUl4LBpC2FULbQ6JxF2biNC1CEtb27r/5eDciXEdDOdZL0rqFgsDgkKnzBBP4uE3neoeh6lPhYP2
b4bUbMHOGcs3jH0LHmuzhgWIlt8kHWaRkWLXRo9RScTjENVXcj4aqYEFYdtWPIAX7jhmKOHIy3np
1w7+094KUMTWlEpSw83lNkvFeAQB/SGtK1XK/kPlYaj6yMn539421PjWukPp3Ob6oMssI/JGTk2c
XvzukMIXEmUG5a19vIwRGogh9Rgi3GWp4zMJ0TPoHx9gMUwsSQaO18YC642TZUmLB0Jb6UaMm1cT
uys/BwbCwIXt7hJQiGvwrMv4aAAb91a1opyh+QkIHrr2VI5CK9kkBcLLlqsUFgfMIefS8t5rmHph
nD31+a9oOpCLNe8k6m6l4GopZqK+sShy4yulmuTEL2QYhhKNOYE8TBX8rQMMdykldx1Q6gvLluru
5sKqOQnnmkToHrLL2c+U0B31o9D483oYBuncD641xjKF6zEU8K1mFIBPAR4/a/g0AXO5EtWhUGDE
3iReadJe+bD0k/ao6fcCDjlycEYFkrNyY71qxKCnXmvyzDhN+qt8J/C6Kg3RAwTFZ9Za17TQbr4x
mxfF8SCYi2tp6ksQnvwDy80lALF9t/43FEWxK9xzhLkpVVPx0Se0rh+nzC6NIVd3jcUna44wLwrJ
VJWjH2mMzft0HLU8MXbiqb4vaUGKG2L46dYXq+Uwx/uKEV+u9TWp6T9PsXca+bxI1idOoSrWz7tr
XI6YkJx8+IrSYLJv1LtHf7vOQqsKzIhtFl4bRVa/psABFGb8+2UHP1LGnThp6/WpuI/isiqMGEVV
qoDT1fPTaaJVsFt8nR/KosW/gTL/Bh2q1PRo6Ce9ZU/P/ikOTV0aj9rPqXbaiatcCCocx8uw45jn
++1ruhBsjRHW0wRIxJivn7vnMhwMGoyMViiI9+JTOlAPgfbOGUaZrn7Gtcc1xTKKYMPaagU6/nQP
fA3VCqOh4KwzhqNCMczsN1COHZCY87YoQG4HAWmVL+gTtiTBqwMcmhTkbyINpmihW/Z7UP6q6nEe
PaJVwVIwmgqF5iOLjsuJ1fH1qb48uTAUrEMrkgLnz0dGQdSPvVAYJR7JnWlNsdjTr1wHhH8+p02G
9ql7v/8G2K+2IE1C36fpIqmSYW2ROg/PF185pzf0wGAs7YNytw58E0wgz1mMrNLQrFSD453Smi2G
41vB02pw7ciFq+f7UOP3fc/gU/CVfe0rnycQLSjMsYoJwhd0xFTpIeaFwqrdxZyf7xPuW/DHnnkD
aVPo9MMg8AE7cJwAtfymzTeF5n6ttyGmAEcrz6WO3whpO1IUCXJPWiKvbITrwu/GLUt2rdZQ91bX
vJ2jzMU4VUyS7/mOWCnwHYncJt//Mf8gB9DxBN6sBc6BFUQ+y6wTzjdKg/D/SxlZxEjlhPinLnS7
SDEpJQTS61nmuaRupaBBrVOZ2wCLAznQXF14zDjXUBi4WVzT2wBGwiT7PhnFxBBI8jUeJWcKFl8C
REspXatpEbtye1YIsj1gZ0YyI7kqQ7wtuPX8zts6K0zrbK7igMlrdPcC0UWLWGO9Rt5YmuhU3F7/
rWBf4VEVlo0oLAtQv39xSDlkG86yq4ryclaLzOcFY7sTm4RWR7jVA9n4yRjMdrOIQGXnsKp227bR
9dkInC3A2nQMDYQuB3UgLxhERGAA52BmZzPA8thCtJW7lULRV3bZYH3gzKdmhddAAcwM2g7IAkd7
zJidUgBaySuuC9WEZsgoc+a765FhhQ/bljpVsjB0fU15A4IEHWApAInU5hkhHZo7GDWle+10CxRA
0b6pEFV7hVTTRlt9079iFHGF7GAugI7UgxOCQxrFx85KCmXWOdsgqTDs8NLS6RaMsDG7IhsVnW+p
0V6FTZLCtTx6i74XRxR9VESNaY1GtS3miUQYLXpyIwbGONhV9+iJYmUJ4LfeKAioQpKJp6bR+je3
/l1uBUhXyMbEEgrA81j7HnYwx8j/L+Dv+loPytXGS9IDJvfxOkGnMDmNc9b9LdjZpzlpv7UXXwBy
0U/K8t/a7FlvIyVRFs5gNVPAJY30RZLHrsuiGdDte7Bp1P0vbTfN+bbctgxoP9X9v/7T31WGRPsi
G62Jy372FZ77BXl6mLs2n3+gYP3nN3uG8fBuE+7TyIzjDHr2jX5QKPliPzsWxYagTj6/YOEhUbH/
TgBWcTi2Am2DkSQzBSmsabK5slktnuhw60VX2IdsZz389KKS/eKxs4ct+P3bhwteb9CjEbkE8jxV
PHGgYWlWUQi2lxViep00prgRqGCK5Qa07jrC0dCpVr5OwYQNOWCUV9Ug1/Kui6HJ08xCzlBn4r/D
H3zEKFTUd4AORfjyyIpwbHcb35sFxit0H1kADopf2ZkxgQc1JY2m/inkAKS+marCZvSEuuKeqmHw
zk+PfR4UAqSn+YUz4LwLvvkz+EtjWlC8knfw+6/V3Z8Gp+isNZ6f+RiP9Ys+XpVAG5KVk5u3uxf5
0QEezD6nqNXNzAn9PqwB6hV49CEgYvJvU+FlG+z5ebl6ZONfrvy0Tjk3VsFwgeDnai6lxh6J5te7
M4uBnlpRRYsQkA9iuFR1XltsBtTYGpUCcpk5Oiu2oGWAIQQrJOuWnGFjqeWFBg5BXbll1Z2jodTa
Y5RXrg/gZPn/ADckGoDzxS+o7obUFKu8EI5MM10JyCiT0vZ+ixIqav6FFcHTCUXGK8XHnw8ZGhD+
7Wanu+exJp0zk2z3zRMhBLO5texGabG/UXmYt1CP6DPiTs6FDQb0iuzUwdpFaRX/CzCCNVDYUVea
oa+R2lqqI5QsCoe/vt8vYGFguWQkXaZ3E+0YxtB9+w7x6/tbLT/OeebjAHxADKG57FQ3rrK5G0fk
WAtWT3UArOjcWGz9CRr+kAF2dvOiYWFT89gfKSq2Se7EF/Sh2KaK0n9O4zO8CsV9LgcGCsubxuoe
ClrLxYAqPYGlepi7w2RZ48tLIsd2GNzLh1Vza8oEiYhrTiyP+pv4627bGYED0HsX8FmUEQGeT3pV
vUPzPs1eYifuHDzYoCkcTxLgfGeHnBwxs8QSa+eOiFjWj3nQw7jM2dWDxchH4cchjbMT08H8KIvd
Hfm33ZCe95I4XIuWzw9w7ACklNQzDDatQZHawDkJFk8iitgF363BK+S2ur3ipBbeLBP4QXpBRRnX
ZymyxKY4HRg1s/uKLDg6KbwflHAt9ei2PJl8kPWLJ5YVrWoANgZaEvIllN/Uya1mRHXrqmA8OkFq
Jf3pAg7iilvUVEXZYPoaJgtxpUu/1McZsEZSdKyBitXBPAxhh+nFSEWl1FgF1l8PhrcPb6jO1JSe
aQE7EORlZCAy/ZpgQR8FEsMrnqM4CEZvS1qNlZpLfaXkAfH37HAi8iFeOYbf173z3n8W2djXEYE3
giE1YXyo7GWUDkVa8D/aTRTjxSqA8vp+W/BTVrh8Oaaagx3fbXLpsNuAlC/049TcCHUA6Xefacw7
M9lZfA+GMduHBSq1MPqTUz1ZFI1RsWVu3JZoF2qw4MdYtOe+9fxg+DucJW9GHDhlaGhfSFg3m1/G
J2T07gqwH52tLs5RFifqr/kF8aerrIdeF/amDojevGLMd0+qSldqwmX4ijJzzq8yELhSmoBfa7Dt
OaMx6ahAxwgkIh45XdRy/kT1JdJ47wzhCmlbyi0xJtl5sXFi4xwJwG+2eIMxywVoOyNYCJamy98Z
eAlcReAu22O7sf558c/orVx62qafytmoqnCL1x23CHinbTSqM6IMqG2OGC4ktZNPP2M8qv5YPFuY
c1bWpsGeivNAQIjmJjwOmFPp++2mKTJwR8Ix22IHa5XNNVlT33YEQh/hUIEE5aKurNDXwRU7gLHt
pVY5iONvmmCC2ahI6k8AM8PtBEFI9XX8qcsYqrnTvzWMIv6KsclJZVVFjeJD1UPpJO0fo8nQA7uw
ju38cW/ITwSZ5wFYZN2Nm7no2Yk8glhMQQx02AgDXd7rsWCdU24bVwpQ358UwRDArirN3/qB0730
ZtIgWOqwhHYO0FNlK7USdcOk2FghhFtzkGWIYMUrPTfMqdvk5a52C33GpW8jdG0Fsycb4pXzDy3D
SLXJs4nzJ/zxtHKdcjq5nvlOMuNI06UN9jfYE9CY68E4t/lpRNno3t8XbLyON6TmEXEP1kAQr2lO
6mGSOfanLLsZEIwZmQmEg9HCaTIr/QuAkJbhGgTGePpMENrrUOLKsVN7XB52uYDx1mBT41Rr4+QL
tg4hyaCExcFW12htFfFjTqYTxaukllPQ/o9GUKCFB1CPEKIYypkw7jA4l4NLnDj6iDXF5EqzI4r3
whfAD2ESoCpJKqkxJeyeuc93mJqohYOKPj5VV4l/7cDR5A7rZwzSe1kTXzZoM5GOysnRR4ORqbfj
ko++NZhoCvJXOmLeJ4keqWGIRLylG3z5sylsvc02DzL7kbCL66ncZDrmY6ePXPPsrRq7vNRhnsFP
Db7FnrTSriTmHRtQ/bwLRfRU9dVd0YfzOeYjDxeXWR/FW2SXXDA+wSIk2GgBZvLsHWWZ3fW6MKdy
Va3TtuOJAOsoLWhKGitg0kOIOXzcbDmlJhlWPkXlg5ovWY4uSZqer9BMO3AltXRHzEMbz5N/PcB/
/QSN7A267ic+ZUG+gf49YMboVVAHLvo5Y1EgnPuTX3MBXcVok8K04dqDe4SuaDgj1Su0C4C0h+yq
zuVz/w028WuQc9ef6JfwQjjbmJ62RhjzIXDXRKiuePvKMT7ZTtsSXKNsk8gmjtowTxq8RVy1Fu4W
7fM/Na2oOaAIOGfHCngKu4bTkLsJuzeNOKLI7vbQbyqwhgnpobBOnMla3wqnc44AZvRtK3B0tPYv
gvx5Z+Yz/Eiv1g5xbvdz71AsXS3RCPAZrw0ca2Vx7cowFYZ8evzkXKxUJj4dGuWehVbeo0zjZ6Dl
sPgqCU5b5JH1RUqY1uHLSGCevAVY3fnadsj6iCgMr97WTvj7CMOP8codmuAuNMeNQwyrF9XuPV1U
C+2g4hx9vKW+2aZ4+r4pIj1bhBr8RDLK6Z95gcEhsyARHNsCnetXP8Nk/rPGd6iZg96361EZCv9Y
IjVvfPYuXiM3z+/HBYmukMBzBGTIbyHPnvy4zvvWBfzf87qmrGYoPmEwOvFd7HA3F4zA5KC+C4Ej
xm5wRkuZEp0Fjzgio7Vv54leruf4mdrhXzdnp582mo6XY1mV91Y2d1xRXAHb6F0zJCTm+EduFf9v
EewX20F666h1aGts7QSfw4tKWqyT1xA36GkHx7AaMsy+vha/Sz7YZJ8ttE4P2AL0aGQXsefMet9Q
Ea4gjLzak186heKlKWsaTsDdgat9smHILcnTKzy8XYNLlj7zVjda1LLYBuzmNjkst4mSXxl8+TR4
RNInbIA3zliVX4piK5OtLuui6BFalkheaYKDvC967ilGy7xWF2Ff/dSI4l/5K6tCBqvcOEPBSP/E
buHG6Ml9zPRuD68gvZtvrsSEb2II2iRWlFDJZ3l8/2DmdYwQH4I4Q8P6E0wV2D2x/0kmenDA5S3R
ZAmqzUEPJusiPrty9/uQpCH/KJWVwqxbB85osETRRI3kzCYAegmXaf4XLZVgEX4Rr90tODtennSP
dDe/f3pzIPXuibRJLmZFMZEd0X/w0wVuJa27WAHxyH4hfs8xMQlCCdtEcz9qSWBQnQkdekQW0MY3
2r/Xu+FUa73TKlocM7G9Vx3pAfy3V/vYSSD96maXUg61Ne6QHUUHSBmhvKCALEoQRLRN3xmP9kWf
M/SunXi7daYriSfTowxfcajea9cyZKwQbJl/mSbFkxpV/krkH4zyK/cR5GUqtpjdUHa8UAtgcBk3
sUMBHep0RA7Ex/tNzUERor2zFiQxyiMaJwuKdZW0wmmQIAD6VZfXM5i5N0UwJEB3GGBMHEzFE8Mi
2/BCi8Jky8TxPmUn5K8MDabrJyXagvJkbJBEp9nzO0KBBfrdq4VQCwvxlldP7oP53m9ldDKoCbFL
LytfPLSJ1tbo3CjTcgP5qyxTQPzSNH5tzMZ/4rZMSHG1MtKZiOSO6lTwIrf3R15ZznSyISdlwiz/
oHvax3JnjrkAWL0jJVcggBKU8g2EVUKtChD5qqfbFEqq4TrxwWX9X85h8hLLP0K+T8GnBVLyTr2t
zP0JhP+1b7C+fQKeF6qXlwiO1Y/g/RvqvMNdu6p7q7LtpPBVrdLDj0C8WuEAoWn67xo+GhhpY9Rz
YDoTihDJLlQudE7y1ucV2BbxgqCc6reDBiQtbo2HTuq/Z9dTpVRxKOfob2OT9/dPY/et6gqYeEYT
qWXWmoDcgOjcnFnvsABOQ4ABoQNn10b8xyWKr4V6n6gnVVzy7iNgvRlv78UhFkKZL4gj5Z5lJCij
sEGHND7f/Cc8SL2LM5SuVYYTe+TyyosQ+COGlTue/KatSmPfy8U3pH4x1uBDxZz4TG/vvO84NwQR
nC0ma6Z882iPPZzTWchKOWwn0xfuKv3MluO9aaikjDIC/1IU3Ki+TiJiTz5XaO8Z9zWKToJnzJoS
Qu2THd+9sSIziN4qTBaUoUjbqha4Q+cFKHuD8H3WUk9dmB/JmX3GHl2fcknwQ3uRRA+M08c2xNS5
tocYUk6fykyzEOuV30no2fiTDLw+Fr/KBmDnIm1Z/dX9zkiWUukompKcF6edX96f1VcxqJaAIban
yfMuXiFMUvOl9aqUGjo/zOjpzcWJmYF5KAcMpUUofgu1wdps2y7+KpQtm9kho4SktJr9A2bbYN5b
V2cGOS1miR42LovS9zLv43gAYm3yXUO6dJrnvWdEJtkmM+pV0KWLliUWdrzwZOOQUh2NXshbHDgE
SrvAXuf+zVQOmRGQA3w8V6uVjvakvrlx1UZUaKE3TYILsmVAEBYHoDjMaB7tCH7MRznf1dpJcMx7
UbDntz0b+S0xW2ICxbY8MfGCdl5v6THrrQZH+Sxb/WFBXMRaNmVcgPzB842zES2CuMnNRdHuHfa2
hspuCbunbPQi4Sd20KhDl7OqdC69bC33K6iFt2cu6WX+B+nKjq8ApDfQDRObf2Syqwk0oZWxQk9N
oTv0GIM3ixZL2i3CoDqzmdy0kkzkGg2JaXmWgkGjqnI7w5kqUGaaKgPL48ybRa7kA6pq+ZV8lQSt
HDe3ZGb18J6iWcW6b097RWzU3+N968PBkqOOV4GyQWQ+YeOXgz2OjOZRzQeBtBZJQIWYBLf/t16O
IUkvEMKbgXqMmmDGJ16mMuAGDEKKvKr+zw1ZNy+oXstTD8QuWJZoWHAqzjlW/EZMPTTM9S1HZOMH
l13y9kxv/Z0WvmUxubWpaSY4/0KXBrk515bEUNJTRHnsxDlU9SgP4w3/gaxyPD0g8UU/5fVGfYNp
6moqpBmmXgEoZid6CmSaOPMqz9DSbaEjaBjEdODNbodjaIgZ90zo50XZ9k3f7NpRdH7RqwcmFene
Ga2M6ae7P4hVIp6ztwb8dlC6Ymhp9R34SGxXHlEeu2MubCLQga87J0nxjTENqvtyQghwgDEpRJrp
ua5Q5XjjYfJ/3zrqoRiZXUs4Bw4zo0hnx/lgC1KUoZCEk2z9dK9rcymM8jQODIGLAwN4vhpiVpIn
Tm+9TdH4OcxX38FRFwL9CTCP+vfoIzaQnvLFwkLskD1Ovq0cCBLUQVU98LUvBCXQK0jeE4kilKOR
fzrjEyjYMUh9PaXTNR0aflvjDqgSoQV9NIXYumu1M/LDadccKFvNS+HCgU8exQynamuU/ZuDOiGu
AJNzzY9N9Hy/5snMTdSXj9Mwt8oZtlnnkOU2YD5E6N8Rp9ra67p3aAWLjMXvA9YBROAG/hULVYZu
E2Y90NlycZKFjqmrgyP9rF1atWVdLF98i2uFFj9KknGiXReNNfIEiQqBWxjkwByO1tfoU3GWsoH+
wzkc39QXCdxOAdX5FnsObb58X0OufEjwP4ttL2u+9mXiQnW0965pyFi/n/PLx2/x/wa8tbBAucwN
DI56pNrzZr2VZLViqZLEAZylGIy+jAW+Io9k+Lko6CMLfnS940sxwIHuDhGl7/J+wsBJaDEubUcz
2NT5lui/5RNAODQ7RCwTrL0Wp/AlAQyiMPeNcQUPXg+xmvJOAaqrO+WAluIZudJLIbCEqT9NIch3
GKuK+hQimYkk0zk8+hL78pSNF4gwvgJ7rUTurpW22/ttiHrFZHyfe+LW9Qz42fS1iVAnHNiPEP5b
xCoHMw5pWUsD6szYaKXAcnzmHrRRsFjcRfYDazsqXfdxfbBvNbtMeOU04KTgYDS5VnsH2OuFUCgp
iPDcbC+i872sqIwxDSwz2l8RCCI+r4D+EnBnyWfqqZ1sxfuR9RyeXr8m9sByfoqGTSJa0A1l9L6C
sgfn1G2U1xdDsCkB4/Q37fiNFp9vXhUbV960yzPmeztAn3ngkId91bpaz9sadE0DLp3Eobggoe16
UuoNXCJv/bw0nKGH9KgE5e4LIAxdxXigtqLEuWmH7XLcUmj/Rbj/MShwhKS37uH8PvGldDu17zsc
e6qkNFTH1Ywq6fTI9oD8oJ+nS2l8aAi3951SJcs6+B3lYJpQubssXA7Uf4O06ObPL71w68pFz1l5
LU6Y5YQ2in/jeU7cKRDxYa95fWkjkc7LbTC0NzTpg6BjGFvaXzfNATLkLq/pRmT38YHKQ0Q6BUEO
YnWMl3iax8ilMJYbUcFRXWpajNG1MwlHGMwPeDUoqOp5juq7hiqIniAePf6SOC/9vJue9mdunFNc
hDNNLMezRrfLIvXXHR4t/teQVjyiThy7XUMmQhqkkNOlMjJED/tjUPTc7kOs1SAEmBqQah+bEMhZ
pADYFKWyvvS2n9xwt6N4hOPdt7rUMNYvycD4EfVR815wPKW9OkNH9/UJM8x3tsQcYvj4g7gW9hTs
8aNPjSHs83hpQn5SSH3HUu6JMMZDiC9V/3mygzLIT9sst02Uba8fqGFGMZjJA/s3mPjY1a/AU9Ho
Hi5tDMSwvnAB3fiNyY2uMGkzqy5hWOpMON12IhZKehqLuSyn6rkcd0uYuB6yzroV4V520Pj6LVjs
le9yuKnvY8rhjkrX7tOrk218vOnKzHJk8R56oAQBt4e/5U5xPgM/GKvOm2QHeZZbbytUWr86wSIM
1CB4/lmvkGOld7IAH0VecwuxRRseb35eW375r9B0n7eKWdeBmykqtb3eM5jXRQQzQDVOEYfhROi7
PulObRN/fya1i7snc9lnGxRE6vjDbIrRimynBav9KH/HlzuknwAoPGUoflYG8lhtX755zSMves91
YpyEcWBzc1G9MGIjPmfC3rGuXXXaN81rQR+C/iJeeWimAi6cRQruHNfd2UFeS+/POMaCJ7VfyoQN
qu4w/xLidT8AMPgzvG8gaayhxe5KUNRx+jF1Xq9XtJrnaZ8qmByUWbcVJXgibvJQTjWW3zuOiZk7
xSmTdmruMoYBot76+LJFnJnhZl3QXPi1qlu7JNX9K5iZhd7AR/ERy6f1rOm1i4Hc9bj99J6RXMyr
G9HSoMhRGA8D/UXT0i2Oum572TY+S+4/xHoL9wMMyHqzCVVQ/vJabfYloaKcP6jsJOXN+ijPoE29
byuHogqXxjSa/4YaQTfD0mMI/Y+ymbr9KBX/OBetLsE4Y6onLLoGhflMfRzeXNSJqE74kXKBPULf
APA3O9cnmzWY8cpsxEC8Q5V+Wp4gwRmkJfwUK7QTrRYXmcfQ0dSUSuInbwRVcCHhznRequNBvsAq
cOS2qwDyz8HgkvD5ga2LisofHKzAZTmXexA6dC8mLXKnx8vn8mkP+l4D75kVEvbMHJeiX4DpnOa5
dglUwhg/my5lSdJ+mR6bbLwLUaBzWQwDitxWgoVsDuq+kRhKmCje5HbEFjt9dYk+8y3bhue/e1pX
KQd3zqeNN4YTLzGtxeixRPSWbzF9oQfdIvL9N/9+Osfa8a1dnvhYEBWoNZfIt7xsOhtdt2kmAITa
095iv81VisDwx+WycnGYqypL1tQUfpj6KXtyUMrCu78vMOQzQi93ZILw28P6cbnVtXmhsn/pguMD
ceMHpybkSL4GXDaN9QxVRaKe3mhNBlN+TlIBU9O76WDl9JLm+r/8pqG8IbPUPZcfdSa5ZUBXL5bt
Y2+oCUcWZyw+oi5c6vCISpXQoeoMncEiTVB386fzwcY75HKKLd7nKRy2Z9WVK34bruOBZkvJ2Ybv
5B2IJNKMN1IRJ6W1RZXVUnxvpTIZ6x25eF6A/mxeKI/GdwWLCBbhBjddVzNnE5B4u6GujDjXMvFs
VDaKLMiQZ05Z+L2i8l6MAp4KYZ/BJgNoscHzJ/Ep4e266RG/pF+5DBtJT/NNJSOJoRRLmrdT+Stq
A4/rDXfgGJO4OrSIWwy7xFXwIoVjMKK1M7xOF6qdZXrmycNscjV1QAVIaofbvRvWlgC+04zW8rub
rRApqIiEJGmoVQuEiNmCnU+VjV4Rpuzk545cv+Ty17dljgGnQbuZUJq6sSn7aLX9bFyRglooq1sO
wtbtdWx6Q1WXtFIL0NiR3hX7OKzN1KgFKStys+6YCFC6OCco+5ag5SySPIzDOdmmrhiPr6rz74gh
S86QtQ4Cc1t17cKX9ZtlzAkM0sk6zESUN0M1FlrdRQ4GK2sc5PV/t21Q0hJvEsXLBNCUdCbIpdMT
PjDt1uOilvd1+NToDo1OF+VEI7ghCisRBlDqOtjLPARa3/EFNtsD4uJfewT2hXcxYcQDJEHgGxGh
0YIFJiXszZVXSMefb1uBX+HJNFl1VZIU0esyjlZf0B2BZ21cCmanGn0DieQbermpja4psS5fviI6
UPr0/HcNANG4qj7pIGC2rAgFyRLQqXEjWOxYP+ygmIvzHzdf1Mlc9u5cugMpiCL2mqLFhKNIytQr
DNpIswNA4rpM6Ce38LZxjDaE+EPZ7kDGSTHLA2JPiviI5BxkhDf/igdTWQc9b9q5sNzJnSBn7ZMv
9U9rBvsASOzbmXWCHmHiBIFclJBULxpt0S14fyFZenMh1L/OATsW9ChIODSUqvMmGvAdlFl7kCR1
JQPkaiFCvrfWqj8ARLqCZkPJS0kirJHXZWEOk0VHPmMLry+U1GGyS1PdP9Q3t0Zn9bLmstw50gxE
hPiua6kPIXT6GSVygx6vXanBgvt+PLG+YKWNqEUXxXB2LXp4cBwhRy2KQbq4NNzLU1t9BFOl/1ui
Qf1H46O/ZGZ3TNzE+uqXtJ3BdhhZDey03lbDgIQbTV+Rm2xS7ZeE8ueognhUKnSUaiSXvWTEDLaQ
FK1gJHGHsoeeqZpFfxhxap5zXJ9mgVnHBFHy88r4IS+gNb+8xTBoNV3DKGwhqUZzGVP9Mo2sNmey
3nZLGYooltdMNpmdbZWu8VgIm65yuULA5VoHzXxwCJ95QFTL1APoOehVppsvks2XYvY85UhBsr4t
JeIjGIhwTQUod3M3qhEUSMHvBrDzBw2DT89ILFaIivVqr6Tkqx8O+9scR7lqIoccEmJSxmwx7abH
FP/o/6kD1YVlJM/9a3/lrkOQ4mBd/gQmhs2xAbPV5a9e/aUZR8UCbmE/hHe1W0GZPOsRDvuDQ75N
k7dg1rY3bAEFMAC/Z4DECVxcZ0+Pebo7jddsr031NL9jngL0PavLaL+UogiJDlopmsYmTjUIkuht
4IU1rZOb8oV7QSwou0YKLbEPm5gNaljVTiyy0JSK6CSekFzdaQQ5CZVYoeUxT6DB7eH8FUm+zruL
DzseUkDEKrGRd/xjCV24zH+hYOOhbexLSeod3UZLeINuAo805/FNPl08F1zumPIMfS5ap6kdxRdq
C9D1KlKFM3ylMQnao7NWXX4gG5NuUjC5a2uVO8/nnb57ldD0027ZW+3JhblpF0fX8V5ZEVND/sPF
8iZCSQy9yLh+u9qOGunhD6xTXkENsIqgUi8U9BxL/dT0ei2wop69SNalJog2hcLGqPDc6M7tLCXT
GVYqRLOHOZdcIP2Zkq330YewLYKhPlPNcUC+rpHRj+0omHWRG8KSdA5xuLsvZ4XawHdHrQtzWgJa
eyVVEQJdYU/liDDfYwC+RrVSzpnhOKSvhanXGVVl1SNYQ55MbXmGwkosJQ4BieZ5zWVWjhETeQeM
qyUXWqfgyj+TUkn/9i12zupbf0aI4LdEFP25xwnSKpOxBh9DsXL//ut8oB0X4RP9HYOvhlhcGFSi
xdsGuppEpav+t4oLWxJtLnt/v/E9UV8g4ZmTb8Ag/6hoxSk7VOejO34uiaQTOZFPBBPkSWPWpeXA
ECjNeeGmoGfwMljGmXv6QzINptkqqxScKn/18FZjrVkq9Xdc+/Evrdd8ymvKwnKsNeoSmIEG0SoY
xuMrCsO9qadEXd3vKMRL9o8jGAwdNJ/eNzAUQdetiy1Iu9z707sbpXm7ZgbfgAe6vGhwvaBYHJkp
fou3Z7kvQFu/GLK8e2r6ipol8jWImRi3I6X4qzhmsfLXH5SMIPYkGxOQ0yavCgnzZST4FqJgNsM+
fdjf9FI4JWF6q4kXJqzuJOPVULI5sU3uh8UprgtFHaAF7Ey4orUlrVdNwpkvzuObwESpM2cpO4ia
RFjoTXl2OTM7vPKraI41PASWI+L3J/G1kSq9pEIgX1wgylpn0fgDWIeAOsmagNibjleoj9r2ZMPN
kzm5G+tNEk/Vw3qPkig2ADImdUU+g3sDNITs0hYEocthZmXlnqL2/hiW3xfK0ppYIv/3bUCN3BXm
GdIJ/meBgHIzqP6hmzM9y+AF4kb2EMMUO3ot4KIAJWgTy5aayiUQc/PstJg3slescXSc2718pw60
5AFaKcfqYXofPTE6L1ce9yOiG9jNcxKYeSqdYhv7QlOSYaYHjy9XCpGYHGwr7+J7jU4tkITjUSbk
Nbwa90tuqjzvvfkCa/gLKr0EGrO1TAzKAwsFFN/N8bGCtRUuXWvQnnbhXTrW4Y+pEKXAU1N7ileX
7i3eBesPnN93k5ywOuZ8BeobRdNC/dGwzB+8o9MnCwWMpnVS+Gltr0Ab/Lmx83omuLEkI2oOAIaX
TnP1PxUtfh+0S4GD+YiqrhG7bDmNjWexP5DlQCtibQDOyPT67x2IzK2ZjOF65uYOy53z/fOUxtJa
t3e5jRbDmGTV9Tvf1+nayX4GPcD9D76q8NVtafoQMTPNeL2TS4i/KgWV4f2H0SiNEMSF2rRob4cs
fhcr8cW8VAImF4TPXCWvMiEAy7Tl3AflOTTyqoN3pWkOoRlifYnWf8MhXGDXdXQOUvFqNTA3kLnH
g7yd5Atn50q2bETKl0Led/LebQPWSIUp4rultAZ888XvxCaOYVdcTDV0ZsXpag6ybIylRbJ6Jfdy
dD4neebx24a7OtHSUk9HseoEANOwHIc/z+DQV9kEw3TUQrArO9lYwZi/z2uQtVqreK2CUzOH8Nod
cZAZQkYGMC//eIdlpiAWJasDlIGadLaO7z7VlqRMvbmAyI70s/Zr1+AtBXbksfkpaFGiZemquCcS
dFe7xzzE+Eiayx21aO6phjSx/UUoVFNSfSA0r9JEy3g+JQVwQQZ3XgtPFXOz1siHG3tLv6uK8c+d
uWCOmmZXWPdCuetfPMqeVJJ5cUTLsIlAF7ADv0o7Fmy/93+Bui+ISWYWX0uBPkIAQXcPWAl98o8g
ShfFWKWqCKzjM6HqjHVWZyOCtbp7XlXvFDn8zRaMDkYmV6rm/DT1FzYg9E40NzfmavdaYuZItTSL
OEWG36N5Z2sbqIOYuNRY8Fjz+NAR2bCZud9ufFIoshhTyC4/HiB8i2ikdzvIDWcc0jkvfPVWBYbZ
oJ+CwT6a1i5qaCaASvWRDULjbdNq3eWQWKxKQk8XQN2zLUDOq3e8b1QbU8oFMSxj2riPwOApDz2g
Sru1iyhXwDkdrqiLS9n74EcJPxP3tJBIvYn8P2tULx4L5gOSN6/6cfKZfKqvJkVuG/Oqy8+cjGUt
YGYWqjW8ViaY05w754OFYb9tC6BMjfNEs9B5w6m1QjM7EULei01/AK4j9RnlPeW8Lu2Dg7HdMhLW
712S1GV6qmZo+DCAGcB+yJBiyxwa3LGVXxvatLXnAWV1+/w8xWb0zsQKERUE5ChRzW57BdPPqJIM
LzhB6uFMyfdyk5jH3EolchlWVzaXdyvyL3y5Tkr9RWuQkIcr0fHtofc16b0Geg0DUM1ueNB+9So1
zaTG94UOUBwIhGr+z2QpZK4LRhwouT6C1WPELmzgN+zZQoCeHbn6tKLolUy4v02rfThB0YvPd4Hc
VowajCTDWJV1ry+51P3OrVk5pZtCOjp9Sdvm2eZjCR/GLfQya/3Ce0Dt7JQDIzKsRtifi+L7K8vX
uWNpf/NvdUmo6M/Yb4aOX5tY/PBrIQJgkbygcymqwoz5C+3a8Z6lsOs71kKg85FTjTUI0OC8dMcC
pXDtrNfMW/WnJtpHLrFCeIeJeQCmYTmRqwgUZKGXUMsGBEaa9OpjfQ69Mk5V1B6YqA0EJlj6l/FL
IB7E7tqi5bkjhUUdFLBKUQBGlXNQqs2LWrAIBsSGkm2B/oiFKOBEu1bbqGDS9vB8QrIgjAV5vGc9
l0WDUHMXQwS814NB2Yre4pG9ZEndwF0mHJNCYxmjYLgp+b2el1ZhtrI3+u8dbzs0s8UxaQG+IAzj
2PSguaWYpPKotkl+5M2CuNl1pjvaoh989MWqGWOpwYs0uyO3tftG7Dn5P7iAof+MyJArQUki6frk
cshI28qsmLU2rGfj6/VbsAJWMKsqPXxJ6KpJegK0HIEcodsGMgx5bBi4VLcj9+ZtP7FlaunqkRj0
T2MGZF5Q2AzMIu1SDoIFlaQvBeVUeEwvea/TGIqWRuXW2rpipv1E3HMBKWviXuvVwiqJREkim6Xa
cLgerqyhjhLmmnULD4jqxgMMuOO1VyVicSbs1KyM432n0DU0/u1ztybVOoKC7dQqYuI0wkUNhNVc
sARIN9idAZrknDPPqWKy8j0K5FcV3evM/Nb7US64Xji9NMv9fx6jll3P7OmkjyYqLGnbHvB8tPy3
jQQegDyTsV6QZ8jlgjOZwyeE86XSTPWUyz8NZKc40tzKKMczeNJe66BCxVmB8pyu+qqEir90BOEw
/cCrnQL1ksGhqdsUWY92WOA2G2qlp0lmvgNYmWwjQmhZ1aJgxTjBGBXmPPp/OIE/vBvBcTJQPKQU
g1P8bOOCNWbtv0l+NrUA+p1doX94+X6oLV3LiJTv+f204zq6tQed9T119zv3eb2vxpY6EYl7KQyn
vuUQgEmqTZu+8J7XlN2jMRy7lQtARDUg/9koZ6XkpVReS6LMpLBC/jetVyO9xeTlFXI+U4iqhmsO
LayG755r4ffM3Nid+HnRCQFf6zcJQH1BcIpdcp4pago3Mf3QwJQbAkAIrPLLw+LISPl4xzyokgnb
xj0GzxF0tF7MqAijj77mg9Hz7Ta4XlLzOPxNvgrqWzKv/Y22kxDBlPEsBRqPf23700X+BHvzYmTD
H07YRcMVaQaS59vVsu/4W60ZNyLSfyzW3XkOxw5148wwlVXarsGbHygnKZFo1sg+uxqjPS9Y5clW
as1KnkF0RT2Pyz0q/Tsh6OK1iZ6oS4FOXE4Q40Kkdmm6WqAQpP5P7BdUF066ocZ+hZiVDXuhxiTi
OTNVeUhfKXksS4JHXS+z+2RVPCmy0h4vujp5I5wkpp/psCC0w8c3BvROBZfyYGFhKB0V6+yBjIex
Qup3l8+znKQL4O4OLavrb1jB59BO3Q7kWw+f88s5GjPo6Kq3TgW1Ng6G/R05PN3FX+/OTQIgMtH1
mpkUUju3szDlU8TVu/U1GeH2MAgA1mAUOJdJhWlyUF6uNETcGr6M+wFfqKHjr+vicRtvueRjrLI0
uPkYSyR1jmcS3/cqPs7xPjRdxy5eEXC2iMxpvsbINtDlVSHEiBo8vYFUaKivTXCmfI6UI1eIlZXE
NDLlDigiBE05roOAaM7JQBl7G5EDCJ1QRsJ8uMOG9DN/m2ErMkA2yMNpQ7+y4P0TkcPLJc5K0vPl
qcUYkmu8l+2YB8wtCsKNdS8hoX7IS+LTvPFk6l58SL4zlOeNsgVmRMqBa2e4ZImUGMi4SmkFR5Vm
T84vShtlXivD9RhrU9T5whjnGgaNnSiPFRrXXOByF9NFMeQWhmfHsIIxBRYJub/bUtBLnRoQQffr
hr8aK1zPWmXVT48H/ykFQlq2jTrFk9+d6HL/uA4/U31DJlbHdgVJuCUS8OPl2BXtkxQXe8SMxAvu
juMA1CW/Lcxo9/hmhZjus72VxluaMKrkgX/E2x2DLOymR3+AdcAJ15WlMihD80lhzx2zJIXjdYrn
8UMeLB7wNVgUCUwQH3gvldck7y+QlUmjMhe7A6EnqtJq7WH8USBSgtpawOwLd9TDUMHjY83uDofr
oonNiw9DeKAizW2icPuS9iTBLUP8I/6a8NSE2dY3t3538rigAaPOvxPfJiw4/ec9ojW6p5JfOc57
32JNaJxiVDbWBE1CaM32Y/s0KgIutIRw8Um0yUE3BFmHDUi4eDjZAg/+thXiSTcXgFQmm2GoVEWd
iATV80aHq4vzxzLvlzkf8uq3fo9GWj97r/OHBQp/DMkpepr9rAhrp6UPn+Q4DUnFkhCSYCrF2gRJ
u1VAfW7PAnxhMisOMFuP1ZbN7r55bIHJjpmB/3TC6OG3y2bMAmHmxgfw0ZWtxCeAEH+LRSDocMHt
X9b3FlvVZxlQ+uNAyEItCYtZqmuN/7chh3F6gf4RzVO0k6eVgnLQD+AiaBRCjTltly0sV1vqY+5u
SetcP6Q7dSnwamLEpPnN+hSZD6tOdlSlpvPRB0z5hrJe5Va2NA6EWvMT6UO4LFPXILiG4RWMc+Hk
pIXJwbhmeghWH+sadEyNyBIob//KoAT1nkezTcJYBfGNzxRq29QRDh43MwL1rPs6ZbJ8WJTPvNiL
nkG+8iQqzJGtAwCvL+jENoCxOhTrJuQcpeBGJqOFeXEkJ2K+NqmSCCTs+MGjC1Y0PsC4urTvH1q+
2KsvA74BXeCzigqswQe7VKOpoHqA8lQFSJd8NyBmCuaYXNWL04kkcjrcYMA4gvo4Gse1x9AJx1kK
qHtLY6G7INiQUVG0eStVfZxSNGtXSGfpMnLwcQgQbuZ6veJGrR6RRrUY7/e0/hpw7cqLR4piXcUe
a8+Lj7apQWDlXo0AcL3fW0eX/gkiLItOEWraLg46PKh6viL0eunwtppksE22Jphd8nQY5znA/x84
mln2lU9kVgKjB8rHSj+1dzbbdxcnDdCLuXgYgbylQJpw1qEsGKsmTOUGh4vy1/elH4MQZ/HALh1Q
schecRI9HhNcFMAGSlI9lTtK7zdNTNPV78hllT/0YB33+rb3US5M0KZKXpWeQ0oX9I1+5+letocr
qNW1/GPnyZrLHmqoGLeSJhCM9h3IFJaUurzOYhrXoUvZxejvovA/D1Vstk278srzD0FitOsovBJN
hYVphws4JIkivawR4fzcEhLlHOfH5IpOsxLMM1RHW3+nA0v467AgVSsVAIm6aN2+3neEnS0y3mL2
/JqfK2jTErF2zwDIfixi+RQ8Tl8EOE4eCHyvE8GRLnByXx5C/irYsBiw1pJT/3czPo6dRqgSN0N9
sFM+ya2hFV0Qzey1F4jNkhqVY+V4qMyD0SiOCi2U6xp5t3ZgErJXqQq/DbStAsPDbOK14VRQDC/R
C3gmY+aSC8MTqLoNsNV7aC0Et3qpCnpC+HYWGjZzmJMQWN1EX8nn+f37ap8ggUhGiziybRAZlKN+
e+I1xsR3qNh2CRqxi7yLxODyrpJq3HJogc4DrEAPvYfUV/rJOardIigsaRVDyp8YCQTPZwnqVWEA
FR+tMwAPuQVy45L5kxUp946ZAQPVR609aWSmGnCbe/JJBenkT8WbHDYSXpeVKHR8uvhVltEaefjY
cF+rCbOkIhtozA4dd+oZ7b5Xn+p0xP3fuA2zg08eUUcE/6TD1wW6kGfTF7H85lUetzwKt08AOHr6
q8GMNhTSS6UAvokkjPSn/FhAB2m2pN5sKkglCjONjK5cjDcywofl4rQLCKCSQus8uCbRN4A8qBTi
N4gC6EfCGQxJVqPMYi5CpqEearJ1i+8AX+6x7R2cXKrWuaXIX1+I6oLhBWnBdJ4oy0L0PiiR6vx+
tJP4x5sBejAT6xS5gUmZUxh0zTrFrv7j4NrEEx2C9JmNx9a4uEO1K+HaLUOloeFCJScSZadKrgWY
IatuQlJcSZhn3Ns2Sj3y+VdMAbKUzdLGII47FjpBXw4kQs4MaY9uTNCTmztstYX+LcaW6G9DG2Rc
sIzy7keNrQGif0TH3J0Ky7a1geCIn6NJ5mHSjmbW4zFq2Bivpmgg/h78HrkSdrZBk4t/eAm2wezk
/OAG0i2pHRtda0jLYoPTQdULv5ySrLB/vBAyXnqjcQdG4i1Lu1qj++9louObmuJMfP2p8J9zqMtx
7dljvAe6bIfw/HQliGLst4rXd9xa5wcrEG2O0cFVkyhmbik/z4A30wNOEMNG5xXlC9P7I1I53lbT
gTQnFCAFazK2ov847tUnDoTfI0/KyIceJfM7ARCo6zSJ5H/ePgGX9co3lo7LbvGzhnvICRdTKlc1
BOM+TtiCKXSsjZ+fTUSTIanpJFj6ybI7gTUWHD6XLqPym9QiTZfWUqZYS19DqrYyI8D8i3U9fzhf
+qFhRwJCTnJdkwKhze8OvIsDp0nBNSvoolZE3TTbHj+dSWIkjmdz5Jvu77Ocw7noOhtxHBhHm5lo
ozwv7yL25Hv0gVQprdt/FnxP+mtnhQyJkjTILo1ZVEHAQThfEQE5JrwmjMC2tXtpSqIT6YsWTt8I
Pz6+Ce8PtSUmgMPBUmV1koMGE6tQQ04saKCyB1GzNHsYCHptQDbPDHdB7/tjsqbRw8riXBf0bsfB
APXf1RDsW/2NYvQU9TKMOMP5+rwXSLa4Ndkh0ef119We5VgjkvLY617NcB24iPALisgNcoeYRgwY
7ddTvRy6sAEwjYAQYKa0qlFuUAvRECSBfb0mL8cz1QV/lvj9kJ5vBz5hp5DT0UnT9hA9EMTxeXy3
2ATEckWxRmc5uV4+2OMjfgBIxG8Bs+NzgpZZTyAm3MzpH47nfQx5AOX6YYdwEjGDAAHDXTSe1VX5
qkpraSDokpKWR65Ka56lobSr0kDvUxuPQewKU/kW8yHM1g37yl8sGIWXhBXa/Cf5wX5no/we4i/x
gdavrTofT5DBBoFGxwSwwEgG4CNE/jfwtVtaKqZjiVPzBYSfoQBvkrPCI7IcRLDyKUeAN1NSwg4C
hoLwBA487WmyieGqfp/PzKd3jd3x1gjB+FMaRwV0JpYZFLRjmM0eqzFgW0vowwRQZlGv237eSSTr
pSWHtnsjcKYvcQDGu6zwq6UK3x7dMN1tK5kOkspYyyuhltNWbGAUdPg0gAxoobx7ZC7+HY04e+7g
M5jDGHNUnDIV9KUb13t6p2h6bt2hd6fI7ha5FdiHQfvLa+HJ97vyV0B4p+6kVNsFB8IgyZSvOdHm
UmWkmyi6ABywI9Yj4b7YU0uzYxv9gt3LDxFBZl/exHdwo8LoxRZfho/jpr8Ite6wEQAiyXfwj2rf
UX0mkstaGFW/rVJuI3BvAY5hFj83NMBb0ChWpkSsba3HW8MXDwAarJBFAK0SF52AkztShhL6Lkjh
S8Udxgn2iaJJqoLPGpkGtTp/PMw2vWg/A3p3kTgrjhjACQR3++egBc4vA8i8b89hRV7zpAlvARDU
YnUtfRqV3/cnTCMqqJZZ0fP4MMqMMlomOjPtw7RJHtXJihkzvrG1a/Y5TnLicd43v7LThnHoQh6N
PXUzCvsYzjkfSwm5e+tijuyH4Lletd9N61UobrGO8jJhyqUUtFVqpu4Ze7Z7CCT7an6t2lths0f0
jHOPUyng2Kr0wAw/NeMKrEoYeybzsa+BmurxNHZb3a/rA+rw2p282ywb29pqm1rNpCQDFNdMxcv8
kyVvAZtuVc8Yq6gkIeuf+vQ4blk+kMZS1YTPjeo63eG4Qpkp2OhpO9jSgkYv0bd3kOhQ9NWRWnbh
eK31kag4+jOpUvY0V+zRvFmO0ARhqu5jtX2t5mcXuXcIHREYMsrIfcJ2PZPT5qpvmeAB0kRfAlXV
lbFd9sDdk0TX7q4ej+M7Z+5CoHX/I56rAsZuFr1c/TdJ715rrmpD+qhyxZz9OJSnZJacDIqFjceT
ggncp0k1naOMHugBRnJXexjoHIuzakUEShr09xvLYdBmvGtW2gO1jhy+l4TlPswAVHS7oZDoK5NF
KZvdbx0xen5hentQpgusBvf70AA0ppz/Kmo9AUQZwhrCXo91zDBV/TLkczVLF4K6Wvr64kkZrMvq
1mQYL1GheZQWPArp2sfQQBIzQ9apR75RYVV2tHc7pxtQ13EWZ5noibAk8qX6e/iPwN4+udKVMdAE
Vt0nc0jF9OpRhIIAE+lF20AVXicxMlpawdIwOC6NcCfPPJrtMeO11zEgamrSxWXp1hRorPhZpr9l
kCUF9o79HlZsdo1r5FqBBiRtu4N8iy20QxRtzisBqAIWA15yQ/fEnKTWS8ESGvdhikmyrZBnaJHm
alpdxo2ZJ5EENVrSSYHI9yCe5pMBVwPGogbXQnpwIMQiIjrKZ34fh5czcTWtclYuC60BAZfPU5j/
YZvJVI7KDS9GCOxqwNnBqAGbkGOS/9DiQUNNZ6dSsUBx3DSZuFr/S31BLVdjru0E/nNjqf5+7iwT
DLYZtQwn/xoSe5KeHKweRcmXq7iuhGXy8NoTSxTnDEVTyikA3GOPasv1sFhOsQrFYOO+zR/5wjyJ
i2bi7GYNJC4YLpDkRxG9WU7x232zH5lNbBcSV3HOpntmUSPmmBCllmDdrAGUbmB0+12NbUHFsGai
Xx7DN23SB8UKnnQ+Pd4YmAs47vq4drts4eCqpQ4GNSESDPh8EiK+1tG8Pr7RqAxXiIfwmLSCvSG1
Rh5mJi8CNB5W8NeZOm8jiyJiBtx7mi7CUegcO1ENRGU9+mx24ufTtMma4/Fw58ARubtR+dwunHe9
3pUR3K7E8RKPbHxJJ3R6ooGxtP+wQ5fDU88sBIAqCHUx28ZKDzmuWrjyJ0mgDr7yz2IY0LB+4ax5
mjknPToubW4V8NCVrUceDWGeaGnPxbyzzfq//hTWGuA/P+Nh+Aw63wxNAWJGz6UL5J9bfkbQKONb
ypqG7cgUL2Xwo//5Pz63QbuBGLcUEoNxcnTOG9tfxn8SMr2+7TBBTUfTMImIspUuhHVu3nir9IKh
sGrHGLuvR/1IujePTDE51ihF/0FcvCr0wqCMEAeMOJo10cAOnk6Fx9lCjaLhpO/araX4k8Y+L1JZ
s01ePk/2ssODiHYSEQwym1TP1B0OJgmfEoAsGlrVQ4ItpUdxqyQQXn84bQLhHRkaToqOGJOU5FJY
zIyzGj8Hir3+hVO/fWTR12BG5SX5pHKIM7SZNvobWv1k7kAd5WWi9nDapiw3qRJX2laT2mLybYlY
J3eCNTzfCva63VrESCrWKwVFAWzb6rj1Ltdf2lILAEi/fOJ0BUrwwyOsJ5CPxv8/oT02mJPLLlpz
QYELdUdovOWjHzbUhLwILrJtIgK6xYHHAzsmRf0JVFSffbZtr/KGrunljXcxxbQcuyx/WMWxIrIO
tasyuuz/EHMwyCtYk4b1UPI3XUSlLEhXTK6ZyP6NOlHjcHeRcJka4g5gopLnRprUVPXLgWN0SSwE
yIyExXrULKvYFG8KM0Nt3D+qlJWuoEpplSSHu85M/trYROiKk4P6jJqNEq8nJDNGHpnmgK1at8sY
JEacjaHk9/cOYOAeKDBAmK62zps2sVecwHbNeYWDNmZ7pJ6JKEgfl4nO0AxdPNIr8AGgVAy2u+a3
zMjMySjO8r5NoTmGpnK6vVEJaJ/W32FzsDQQH9fe3SxOXvWYk+LSL/7qtu+JML4TYRqkfu1J/a9F
HYlJ07QW+D4dOkHfBx7MQya9j2TDr0Q0Ftnt34aL/gVebAVXsMRuET4S+qCKRUruf64311ORAV5o
VWgceaXhKCSr4TXPs9JGrhM8FRSCK5ImuYuyXGdWNcW2ht6+qtZ6kLEfKjUnUKCnZQD/f3+W9Zlj
G3Inbjj6VRlUb9n40tH5FD5KwHCcAQ1LH+BTX2eMcWCw3M3HVl76c8kxZ2CIDn5dgzxy2ycBFGpE
ZWOvKzhGEcilZcY/7zUQlYo28qVIQyvSJ23+6GpFnblPaa3GyvLXP+TDk1C0Ly/KFX6ka1i7dNgA
dS6Y3hv+p6wzJNVyDf50VtVPhdiGBOb+oM/PdyvWmaa3IgpupeyebNG1t1J+73hoAa0q7FKSToal
fAjz19KoOnq86CZMSj+7tMU6C/NdUsyoIkg6aCDi9CAaKq2Od8ejlAMdUkuJctoYdRnKoUsTDYF+
+5P3i4LgayFze9jOxNqyWzfLJg1eQG0BqqpFArNXMknlp4ZZia2lU144Fc4gmLbp9LXEeiHLMY7/
83r6QTLseS8bydBlUZvLOg0gaqEfZWkyNZlrokT3yph9YPLOKFHyqhv6/b9DEvcA954gRLuqoPTw
1i2bxYYD5TxH+8tsReIuYPI7U7G2cJwo4OM/bvRpTK9VkbtSs/1gQmlcs6P+bIjChVE5q2M1kld6
x7zmIJhMaPFJYyffLn/akRll4RB/u6SoCcEbX8RCw9YqYx9FIWa5KIjsQvUiIK/UqXPWW2BJfyMO
AGE9c71pa4k99AMGdQpJp6y9KffIPmnrpZzj7OQNO0F5sfJZbhV9OzyxGQzm9gDZ0F1emb57UIIK
nCSb0c2ZHg7sCUMO+G9F3UCWquVxnpvlAqcNot+6oGCnPHPutlgk2RqbB1h1UKTvhPLEfGT2FdkO
3EHK6GSt7KdqEW1fTEEqipconOGNbk8lcVAXuMssH2DA6jrpJsgu+PDUuHHcLKyS9uB4DR7hlrB+
tSjO3E5zocmVwoxmBXwpHxTVjZ7xnYtE+SZi7Jf5D9gEywPqrJEzN2QFFQfTSbsjYnycbD8h8bKr
Mdc+md73AsrAz2e3zDn6vf2k4+mZ2PnTEN1mRWjjaDat9J8pMdBh+FhULtA4/hyKzqIbrEe274HX
sn4GAxcaN8gH1Cjady+vYlEOTswyQtN6lUL3u16I99l2oIKXm/60tSjl7L9BK70gfsGgurNs4aBX
mh3MRpQwrlkIwhlNMp+n4J4AT9vLhPEB8A0bPfGK4HCShkRDGjvUfofAMv7w6zkTxpjiUJkJu/wB
MmOevYgmhxqm/58oYIuVqiKBYV+aip4HNZ4S//lJYa9deDBf4/KuWwbVGFrulALNEU4Jr+VApe16
0Jt3TMemJquzqumNMfxLNPeyw6DuGwSSJa9TNKlRTvQXzvCTsi7qP9BCk/ZmYWErj5Lx6QG7ee7i
wm3tlNzOcyZ5snnxQP72vzBZtJiMrPR2r/0g4WddGr13psYX74FrSkQbW6471ClrjSS5/i6zcwG1
C4885SbtGLcpotQ20ZvJh9BXSxSSS+h3wQmMFB9Z4Rwmc/+OOf3TwXY5S31Q/0TFV5fhcKfa5XCl
LiU8JTq+AydoFKuTOsqjqqWGs15QvhiXTS2scs/7FPvW0UMJquYNwOePm/tLcslK7a9xw6qjOo7n
Rp74mZAPH+6xlbv9ksx+4jd/KOt86WYrOd90zB0RrBYoZxNGe1NevLPh4S2BUk/FG1+aKstqAdiG
4JqGRMdGBGzt/b3MTYg4ZBjHIj1GRHY+KlqWGnZ4FoCJZ9iJUayKDiNHzz5zV1oNGviaZVHsSHaa
dFuGF/SP+2Q1bTT4LVb5aMqTNHYMT0YlORomxwkNdb6WVv0FasY/8IQyUBQrWacWZA4wzgLDnLUt
/B+lmi//Vm34twvQN/nPo5wj2x2ozs4YTCYku3JOv/1By7/j6LfqlLKhV1ZRE1T8O5CXRQTQseS4
8RpytNW0r00fjeRlky+T4HDRMlQdICwXX77Cdg2cF9ozz1TBkt1/2TtMvCa3z/Wr9QHOx24icrQC
3cB+n3w2+AJiFdZzXOcGVcsWb/3qlp42hg+L8F+h16YXB1AmUQ0t2DjbIc7K22iG6xSGR5o3csSl
cUV6foT8XyedcW73LS+xDgRvDRauhbj5VQ3uXjDNKthKsJsJnB39wyKLiHbWT4ZRUTIyMhTEQ/Ms
5gqTWfKvjcYNMHQL+qRr6SLYVANovT+tLclo83O+xZZ236tMUeqKyFexTMXvHnBGT6al1aAgdNBY
MmGnNKj9Lqa8yt98TlmPlwjhl7uzsnCmuni2nd4Bk/LTw7qNrxt5ENNMaWqHW5keoIsqCF5t+NX/
5n8HN8SfHcy+9x+A79YRD9/L7+dIPaH0qNCDu87W7ruiV3wdu/lgBAbDxy1exi6ruiOK4iVqCZfw
dojzDfImyhopITJ4qPNqNILj6SWRmoaiIHG4Exl7xaYNQJCFMe+tKJ315QF2RMp9QzV+rNo2PvjG
wEgWg6Bnf8+uvmEPBQ/tRVEOzRtsZ6faQVYMaKIhE5yYtslgC6D3MZqxiKWw/3ln5pCOxK+VSwlq
K7EvNPtQ7wiY8DB7Cf8b/YP6S8t+8zPGxpdbJ5snmHF+d2c/R62eMM7y/KzbV2e+px7En50oejBP
6T8WC2e9O2qTuWHVlHoHBl0Vr3hsvlKGGA2OWXwOt7GbXEHNYMOq1Jf07fs1x2l1QltGSd3DYTWV
95i3Te2x4dWc3WtvNXNCe+HXzV2UQOHnh6u0fRsfb86PLHMr22k+nk/wm5IvYTsO0RPVWU+//Sml
/MKRLDPVZppecLAZAo76se4Hzw+x76wLZY+K+IqxmqZGiZqStrBO46NTk7yf2KBXuTEW1TKiN7Wf
jWZoFx4qky/q6+D0/C++F6udEJIFS06KUERt9gP9wVL3iwH9Q9lsKQlVrcdfU+XH8R218R7Hd3k6
S+Q5rTCkBdxReJcT5zGPnM6XP1Dw05qGy9l9YpzEfKDVelOrNvF/Xm0tmxuNgz6MNQwqeOO3OErj
FKIgOhaDc/pGSxuAEjnxxUiPAPCdgNAxxM3aD94EEEQsZC3SQmwV7k06AFdnOKrVt1jPXViR/94l
Oiy7/AEjgsjUXqvo7u7am7B23Fq/qh+2E+bWxIoEwpz/wUyeUmrKb7eLcRHxTFVpPf246KNGV3TT
XEyhEFHj3XFY/FHqFygiNhvLV9NKHelgFNV3nl2vliS9CWtGmz6h92WAdz2QFr8yojv3Snpwretb
iioEdECUelUPfDzGF2EAlU220LXcwPsAH2L9QgwbH2owdI1cTbZTr8VNX5R4BvI+cprseCo8/YDZ
clI9W/6MtqlkA0RBUfLdL732gWUqhN35jfQoDJMBCwwTyAnDlj1qFlVtEEPL6PWbJVPBgKWQUYAG
oWXuu6cEKq99xA2juJ9dgIm0CbAZgBSBi8L7fBvYoESEqBH8wb1JeyLDUTdsNQs8dBf7BO8bzPo/
1RM0RGFqhs56AswPXOlCSVx09W0rhD6Dwq2htS+AqHP8nccGPHDOrWzBMQx1d3QxxD8nUNleYLC6
Zdqzu0eLirb6d1/0zAMyWVpHQL83L3h2b6EEQu0dTsjYBskkpD9oanYQbYYSXK/tb+JjabM6231a
LO9Fe8tRued/WKDxJQ1l8qmi77HNJfE1YB/2vUlB0QVNPwr3lfvq0aVD3bcMHhBjG1i1Jz4/5d24
FJQb8K+ZCTRmbo0JJTMfQhGyz/ZOoME3ZzGKM15fBO2aGgoN5TIV99CB4JnN6UBhmPAhuVTGTL+z
b4HiTGDBUorxQBf2dG5t7YYBxmI8IeHZMej0j7vtdSoqb++fwlfxvrOtdzVfBJTEmC8PushGID+X
xIZ6lIHa6MDXLc8MZ1ev4N/TNVvRuADVh88zHJEYcKD8aF2JU6G0Jl7OwU3A2R5AMt9Io1K90unL
AGyc5zEoRZbTbmFZ5IT2XIWQ/11pVYhptWiPi7/CUnAzqxc1JxbWhoSVPGbwVXoy6qN0g2AhR5kM
b7WGckJlBgmzUJhv9NvyY9XqutXRHw5NUH6bp4BdNabOgYSOMZWPLM7nXBTc4LSYkWbgz5XbE4Qp
9UME7w15X28X8L/tgkFQlkoxvZ2T6YAmwJwKZaeFIRsj5IxNSjhKUamNUkSL02QPY27EWsCvmbev
is/6dVB9ysebAs03WeqpFIi4nCCNm6QWAGkfapQEedLfmF4k8gfTB+8IlDuZFqFYlwtVDLgLHEkM
rmei4zXrITZkQVbkF3GrlBEZZqnoT2lNqtNZh8bcPrOXBKYC0Nm9GHys32ZaVogKICWhJ4V+nIh1
x8jzdHaM6lrDFDx+SYOgwDli8ya68XHZG/X/8vRG7NAokSazMYlGqlWWMiA4HB79blvxNSPbejmv
2UR8hASA9h+osiWklnsBSgI6Xxr6uXz6CrJgfpH7RSKnMZYaqZeB7VGBCDayXS3OlOtE0/2P6dWU
QZcEx/OdTv1xzlr0TdJV0A0mxAIsskkmeGeDn9dWfXrkJ78mcrPpQMg2NsXUqgRqmWYI5Z2rkGFO
tz1TMmBxSb3WKPzfaA/btDYWnKEse7b42qhkVRhGw8iYTWF8RUf+j654THoHRW3NHDJOErE0rY0X
fjb0KSdDdu0lcsJhWHBTK+/Z6ZSMEQfFNJlEzOMZenaO7QmBzxobnR2NB1qeFkc6N/TyX45ukjPT
JI632+X/pVfZ6s76rXboLpLJKZcRSUUoglDR32+urb1M3KZu4t7vf2rXjY05q6iKecUqKBeN4C0d
QeBvsrv1QEQDq3ivzZW6uGT0ulXwPoeOdihsTR/n/nB6DxX8VqtOKS5yaIw3p8CtA2kvyXeU1mnS
2lURXKiZh02VXMT4H3pYUO2o4VCen44iL/h8b2Im3yEajj9pV7mf/rGVrmiYkxLgrmuuypYF8+sj
yCv+jFo12Wz8DBSeWrxEJZXucNkaQ2AKBiO0Huex1zkd4XNJMcwvFV3JzBHtz2R16lRv5GnF0FEo
H+W+tto7421rmhN2mlos0w3OZy6rvzi4ZO7u55VfDDWfnGKPy1QEt6WoFPEmpTUfWCyVrNmEwYKm
8nWVHl0btGbzmIDGJGUb9Xrc+GbeAl/caCfhfnCB86ggcBUExDCKstYOvlBhbigEWSE0KBSTSEVq
YOmeW3nYPJod7rfAFkfWwIZYuHLmw4eiuHzreh5TX9syyLVMvq41GElDiitjXPXZhM7Tv7AcUpmp
3VfYOc1+s763zzwMFBKMg77fDAOAUh2hkTIGf9KPDUfYLfzle0UtjGeQ096dyUFpyEQlFpxpLYmc
JSXQKDne5OMP3wCgDsRBfOAQmE75NnnOe+P17HlkLqYfMr3UpoPqiUEXplKjLIzeWyuKQzh5zSAn
H4FUARxpV5XKYozNaC91M0P9+h0h4e9r5d8PjTiLGTWzdENJkjbBuWy0UNRiBBfugb9jwaj1lTJw
YDk9QV3vaSqT/23sMhYtJAdHOYwZg0CSLFfjJXWMsTP/CtPDtYo9NCA90/lqkKykOZ4pH1h/sHpn
nFWom+4BehDFWsBA+ytr8oqwCpiCv1Rd1lplf2WAN21QohJhKdATXnSlsieDuu1oNVrtgxQT3DoZ
ObaQpd2sP1f28meE+1AEDmYU8XbewJXpu1vD3p4mrQEjXqveUflPYwYWyFYaJZgEoUoEX7vEwXfU
stUtB/486J7zrT0UL4+jibd91BYDToZeYlAzO6kNfJSUqOZWLeKfYr8YZX3OSXAKHiPMUeht2aaU
wGz6FBLR7bY5/HQAT3GoLi/8J4pIdOs5DMzEhizBgzvmoeDdR3jUzbTt/AaZbQKOwJp2UmS0CxqR
uk1Ef7Uox4a6cWskLrKqvZryEbjezEz66UlZDBcjoIBCoGoEqw+xG7GQL1ZGHCdOi1nHKuk4bSf1
iha4e3aSPYsMzrhbyQggDc2u1YNbTSVoDRJDk+dw8u/3y6ISwQ8XmYg6iloAtBaIV1EK13vj+vpe
sMY8BM/rW8J6guFeEgvQOFg+NlySAF5EEmiB06dY5BHYKxkVsgIHgpqH/xlmG/Jl3Zp15p/of9Og
hu3kFEYIGyQDiovz67Ii+EO1zLi8OhlOhpAjxdZ7bisF0R+3BU7HnaW4ryMGjqoyHM8fexnCgROs
kTa0/mwPySApEaj0ERXYxoyrb39t9k+QREM98cm2lVUhQmcEteOPy9VuAQfbmQg2kWrkj2HfmtW0
o8zXKNMXDPphfOZmdnnj04nPnQHBh92FiSa7efdAcOWrX2eJq5oR6nEbArGZgIA5DVlZ48ooM4j3
FkXXzJ/2pHwJo8RYtdOd/zpeosrIYaPpCxAXCNJemO3e8v/t8lMDsrv7EkxoaEjw20lEMpiwTjVv
hDKTdJSrgctiI5KOpHZIybauNNL44vNr1oUuKwhMJuVjtFkA9MflPA8kaX+5I4lugts5O8VvHzDE
3d7aSZsMrutQKS/e3u4dd0WH0WtoYeRMYRRPTrOZz+0kZy23QGKsO6JYz2TQql1BR/xBxuSvzgWL
nXbODPr2bMq3Cx27CpXpQLOmwM/PZZ7Z808oHpzb7kcZ4jcslYlPwTSoBGjBTJ4gYmY8hOKmQCZB
FqReLI2WntkGVK9BdEkIgBvoqL8v/gUwPCaAjdB/ybqXq/cBH3pxu38yY/IEEVuGawEWpqwhfFrv
3kPw+yI3e0mw+YLUonhCKOC5Jx4BMdI7yhMKV1NysVg+45ENNQUToICXJBNrBcQQNQ0Mw9udIpCV
ByDgzAF5/PKAUontYJPVtUZgxTN0NTMBKEa7E6alUnkFsPTLJrOeMIlnP2E8uICsBdBULgps07e1
z9TahYh6rU9s64EoY5/HKzWUaG4VU87h+3DdSmZ3ppKoXGiNZEqrVUIvHx0AVO/llqHuF25UwgPD
vaXmGxnx2AlIc9dijTIiMYB887kK+Q+W6wN+QVecoqTNebG8C0bNqaCPRI3syH+4KgpeGMpQ+E29
8qTWcIqDZz3omTOvJxnGTGFgAB0gBim21FPFpcmSfG6mpqYDWhGFSjtHeUP/LJXWae6RbXq0g4xA
AkM5FtrhOlwTuBevdoUBzslGxtrQB3IRWlZNIb7o7Cy8ouzQJf5baa5py/vPlY6WfBCYCZ3z3QZc
3tgvWM4JuLui4YULtsbeps8eORcnzevV0n8tFzQg9mXc2efleGZ1I2f7OUWQ7o+IgTAW5kIjsqLU
ch6tqAn+RcMNCVupsyDPm+Go9Bnusv10LDkb8sLLzmVNx8HaZmVpyH68XhCJlvCKuKQOSaCzbIcH
HO5Tk1/MHlT5LKEMnOzVRQDlzRVlGDgnv9z4z2Lek+J6bwJ6XFOqqUiE4F952QR6AlNfPnLAHeyF
kKy3S0DVAXu/5BqMYs/IRn1/gi8enLOg8ExZo5Nj1I9flgtsKQXzaD8yhNAPP/BrkVM3OMj/CA5u
QMx9BJ46E/dRtZZwFQmzQ7+HwIxkKxCQGvkbevr1pwEVpqMOBZ5PHlJXsC5FRbAiMjATadrPAVm8
9pqNJK/oOoQI2LLfC80FLo5gN8/Kf+biUotzBhun6WNb10lxWDFmH6IBdmJFASGuUttaYtyqJCNz
fPuYu/81hG1EpcdqG+gGwQUO2q+e83JjjA98bXsANxEf35nmE9i8Gk5ndB7GJC8O88940Lyet0JX
LbGtJeCC6p/OkyJtck01x5APNCxL//xXqTRHD05+lEuG6TJn3wIKzVqtmU3j5Di1VH52Ornq+h/f
cbeaSK/OPjMJY3T9VsmGjSy1M54viqL0A+HAMVFIAGHsSRF450c5eYHmVI6SpYDs6x6c3fZ9IixZ
1KrSzffFbpgNkjbwnf3J+K+RdK0ZBdcrMh0aRloV2NeItZsXG/7FSKuHzlgXXm1m1PChf7wdOSOM
In5KhJvr8lxlG7v205RW3aKxtCjpsmYoO7/Yc4xG/RdWC7QrkIKxHc5dhqT5bZcDj+L6U2Y/adB9
KrF1pbmPj06M1Scy3lCp5hv70jMB3YtpPVNa5MlNWOAahmfV0MWmw/UWT+TrRt4ozvfGInlqBbfR
HbbZQc0poTY/Isf1ivb3wmSmZYwnCd1Iol6hTvOJgp5gF9gycUQRxes5ZwfRa8nSXVrkOnnQcBYx
K+jHjHsrz4kUuzbs3Rz4ffeyOC2w00xPd6YqgtH6RGiM5t98Xc2MCAg+0ZY1Mj3UJzTgNP2g08V+
BECs/UnbW/nX+XJIoDzQalHjhfZTUE308pPcdqM1G0fb4uQYc/dzsAZTjxbC+935BrmpOMttJKW2
yHJ0jMzP7BOj8sAw+xcB4jnx/09THimjEebOaF7XVeEsZ3yH5czHYCOSZJ+Lj8DDogyBr9/llmLB
P+ebj3uGn3heiAeT6NrJ+6dqr8qGP2TMkCRNX3dEz2q2ePqB+cPKEp+q7mbwlCmw8SiuWjarlUel
z2slZr3cWJduelndpS6T/Ni5DLYV0DpreVYWfhNjKMflVKlduxr9TzDJZD77IpR+F0fLcwxHR7zp
IFGtsKta50xpd6S41OTSSg1oXpBDowA17oURThYZyxWAWT55v6GIUl2EirhdpRAeZfm9pNCrMAgu
DB2bq6rCkM/1qXan68AK984saXg0I72Ag1GfsBAlnybelJhtCLwn3ZHrOlW6tG6zEOV/wsH99vbL
5/9Qzu/WdR4DHuh56kMqI5rncTIV7QOFdlcLVBKs9HRCw+Xk+IBX4np1l1gPgSWcSPjG9IOeGuIZ
8rtnejm6rAYi9Q0tvE6hvze0RzhQR6BXcfhNvrCY0FWfs7WXa8NSIKlWerISvwIonovnT+65DRo4
usc8pgRgCGADqNPdirVyHYwNgBZvk+jC2EC+p1MBGQd7mkzvn26LsXmmz0uoQ2Vjc91+dLeU8YFs
yKKX7po5o1ooUfmLR1VByJle/ktB+5+x6Ubr9jxW/pdXB/i4z4rAUoZNqN9sZiZsjc32NiawjY4u
VvN0YLE8zTGyEk0AJ8LVRTkLt4Omx6+zsVwhz67+9xK0E/x597cObHQTY3ia3NYJgf23NLPBYwab
q1/k1obzIKE9ndqJMzvaF2fP+CZtpmmIZc+xsaisWA3E/yWUfkbYYUVJImGJmTmyEBoEqrMhqN+B
mTP75owDGyPOJFM7dAUm1PFeV/rCkEU7hTGiWCx8pSg9sRKZIJLiNOQnWEEQl89wCM2yWqjZM8We
kkouHyVVos0je/pTpTvTv+sMygy7bUo9P8PWj7aWoI+WPLORnJrtvNXj23Up3ap1Sbl5oQaYliU+
kwmR7sJ8CZcV5ciIlhaPxdjNH3IDne11qhoOXRTA7+39wOHAlRxEBF5sh4m9bfNRlZaszrdJuyP6
VCsU4DNcOJ6BbF8PJsBF6wVGWpl57ipSFtR12NJpvX1JLJFx2fuWLOa2z276E/nwmXsfBCjkjPA2
lR3DWuHJyCh/VP+3y39t5SGhM53CvxWs42Pi9A9QJ20j/8a6ZyD/S+VLH6ea7Tml0zgny7LPyqgK
B0mEdt1ABNVfUrcpjGkvsFkxdA8NtFlaUmniamQ0qcPqSm8YrgJHGJ/xxTY+3bThuAZN+SJXSM70
6R/IvXhKEWbG/R8/0+VYp2FBPxTyjcouQx8+Iq3Cgv44h6td/iwZF/qafIgQvsLJVA0zu+yMl0Mk
Q0ajMYhmWn3/shYEHUxCGdigxj1SxR816KLBZlMEJB6s9fLVIIqWdun94DPgYXZWdsNynmj5wqut
iFrLnbacFIMa6CXYtUYTdwoPeyeULmeANJ0StfbuOSPPFG/X1c9zN3cGWw0/p+041wQE3OdmHRqI
wH7qYfu+edPmi0QdwSG25EpMP6KE0WXfKCxkIg+Q1N7Pfh/pXbD6QCJ3iV+7BzWohQLq+m0hHHRR
cDslbiwyrUwMkI2bJ3CgoYCN3p0wis8jo/zTZuWAFp2etlp6gDdoJv+BoAs3cQeh+AENLsBfa1VI
4MUCeOKF+3XT3FcEFgN/BCJ2At8g0tM/bKbaDKLUfS9hFV6PDaE1oRwc3vb+RxLt7SoiL4gfMS4x
F7Sjtn/d0wIsTKo48zlnOkuKPyjbICYpJQJwjuTSDTDrL6A7EPKltapLdEGsjFk+FOh2I75CKwAF
Ri3zT24S3v4bLdT5zsp1psxtQOpW/w9sUddIYJryNWsiCe4kqN6tsVfdvCvxPEHKfmbmfBh5jXBn
BArct94iGjuJM3Es9y+OUe98d22Vh9izyWl1xyAruvAGVAGvOCB5V1dwJTxEzxwJDV5XAIuh0Exp
lQSukFmRj3gOBIbRtbxS7VWBqW99pcX31EjhpA03tC7NK2L19CfOLdT/FWvrlHyktqUfuL0lZcg3
8itn43mAodveeW+8XQAs0pjfUapzyqbvEqF5CnV9yfhhlInJF2ZxKOXGFzjae+gGxiFR/AUwFtMf
N4ux6+K14L8Rge1vUWs+FKoKIAZJ1JhxwGpyOMPHhDHwhCi8SeJcZuqYksij96ywxTnxkUO1IJy4
CvCAzLW9NO8S730y1vpv96b7N3smPDbAqpHeBg7gBK6nQM6w9fpF4DiaSaTZX8s6/teHNRrObbFu
AEl7XI/sl6k5BKTKpIoP9Cw0YJ3YM7lBzNhQn8Bopd2bcTKA9DNqClYrkxzUD3ZzxO9qESFo17uB
95ZkPkiZ1c8finceFm+QGNJeMNFPeYekoRgWe/HGewrLfgcVmYCfS7G74ICrkShbcRmB30Rqf+QX
qMTklImALmiXGvviQR7TlFhwx2cmOjnz3iO9VHIHmZwgKTuZDAp0Q4sUDm0kb5WcMp7Kfq8jYMd0
niwF67l2UIuqI3y6/WjBHSsCoT78vDRrbQGKplZOZKflqXYc05xSMPisSFVYCYS5kXWRiyxzH2Tk
3ufQEd2QE6SWdnQPyrka6446zR9bLxZZOYpmD2EkvxYJl4XHu66q7bfS0xDgkoz30nQDqJW7OeNh
fpfGXK4N+cpvRmGbr5mE0ccZALUWDhIzQ2Bu/QiQejdFT3AfAr0epI5WuqUA3XE/9k7rrnMp7qEt
6WL0NS4qEiq8IAuIHR9hgOYDw4gja0387f07uAGxFx7yoO7+1HqQEQm6Gp08fhPgFEBk3sS7EEeW
2zy3/UfLIOaYrhtHKrghhd+XO9+azxEVBwng0BYtOGEsoRelW8mGbFqGSj8cG5ucn1sCDZF1XOER
OA06MuCthwNVqppuJte1JN5vcI4SFAmpt4GqgLhjO0pendfW4EG2DlG+HjrzrYi4bMDu/oVM7MZK
4oL6t9IsHFCpJUOO21m0kSvdqs0U7fkIWDb/YRQY1ukaE3NoChtQLLNGwh0954wC4MxuHY/Vvjyx
2k01FKfdZvMNLDnd67eINDD1DUx51HLWdA1/9nBjXJ0hznNE5RR9nDB2POu46yf/6kPvpe3yTJhN
qWjzE2RFMQ4hb6AFjrs5CnJrkH7yguTQf5+1HbC6vy1R1U0oJDGhac052Oak9COGEYLVJ+ic/Alc
GZnCMjnCZOHnPB5qtGzWFxrZ57xhrnwxIoKb14ESe1/yUt4y0l0UloF50AEJpBtsod5hq+SnFK+C
ud96h6g9i5f8xB2zPZVY+NNZPnlaZ0fC58p9sc3pPuIzINDVXbs+bGwWJIFdbnj+RDyblARAgpBG
UVcHATAGpBEiRj2qyyJiEWns+QR+R2vly+DgeIcLPU3cV+gF9CDIEMkJAN2hFpWR7A2HT+KrGDUK
G86XJppjT+8uTZjsExvEgHabkOB5ij75jBK8wpaG/3IQ0+/RGUX7qBWtEWt8c1nlm1q0eXHW9mSo
eCYWnZKU5MzI0fL5n5yA1v/tbMKqmVplWcRNhI0X19q86RacwTKCK/Kamz+J07Bcic1XPGCGsXC8
hijHzlWW7kVWGkCbLMu+oDH/t+5fY1B4REGSngp1kHLLVHfSTVSywbkgKAv1iPycncCDbf6L7TIU
i4OvYuq8H42x9Aibzxkmqcvzly97AZ9K05VWIQrYdxQvdujxp3DA4ZdDn9aREbi6FbQwjAocFsZC
zv1hFLLfohPtubBgaxzsgBPrVCnOKiV3eGDTTTlgMCwRei+z3/AWnswnhkIxn1R0p9zuUd7MiRik
Zhnr5W2iWKhd+M38L0AUj4ZtKSlx694k6xM/YDWS7l9UCIcQdF7k7uUUcgBICvdlkQf73cKpiI3z
w6D4DM6T3JmXVQyDlG5VwFw8ly4ORNKV2MRJ0PS0t2OBmHF+EAyGAjMHddegMC1t1gtbSHhIltsy
Gm8s9uwWkiQl+CZgCFtt0gACJnqRMigmFItvOUBuSeJAxK6a5TD5qZP+vxEfK7R4IfVDLIEUY9qC
Y6uqLwU4iqtHTELFmKveQ9LtobwRz8/5vHVxbkHA9hkPreNYiobO1pCjwcsSA4R3uz34ei1SKBwU
IsB2KlRhkaMcuLu5UfoBG6BEJaNTKtsDYucV9H03P4aXBc73nnS3fdlhJIJFvX0nNlLqQIOQtkET
1GsM7pEpxW2zcq1rn6JwDj1JqW3xDjwruQ1o9PwGVkdZjIXdDzsRaE/4jApcDM2cz+/Ykbn+dtVm
/ouG2Mlkk6ZOkzOyet3sEKp1IiJb0ycBc8LdGo8l/MQ5UtF027n38NrUM11lc2c3C6TIr03+d9lO
BzCl77TmpzVoOKlwpK3/GTl/xwueC5dnYdIiYvEM9mi5ekkTxMxhWHWkdV2zvAclrXrSiJ947oOL
lCzCbRCCIvz96811bOBWYmV0v0YKDo1Mh6ZYKupps1s2cVNwnlgtWOOMyXs0cArE2oBwD4reQQ1x
9if6Kh5pnbP5uW7ItXzaxToWnkxKVWQUg2mv5cmIwMVD4JfaYsZ+VLXJFKLU2zSW4JZjv+DpwBIN
Sg8Xvsgd/VVoqfz4Tx7CBH4hoUr+PE7b5xjhEhCKei736Crp5+LUscb05qQVzp2ER3xJB/pE0qvL
fhZt0QZ1PyMnH1QO/+W3gf1zGdyO93tjkGNV/rEImamEt/V9exIVa7UafYiKp+eEKMDCBYjWvdE7
OHqyi1AcR37NYo6jrSfsU8uDU09H0bdp0qrUiqs+jHf/SwtQiFlDD1lUGNUfMFSxTd6nv9HpzG40
wyrD/v6hSTQvj9S/BSbta+AGF0JNVigI/+tE1vObpQrAN17ij4xsQ3fSJRoB+EYmrtFe8iyQRqNB
jCZYuWtRyWbBgOqD6ZW5ir3LlPUItnYREXsYxldueoBMFQ6s+0YC3EIeQoNU+ZA5PZ0gsYNOrRUL
WOI24Ui595Sc0cJqf2ozqE9gr39VWv+Z2OSWrBZcCvoi/B1sHNMrGbJCR7drELknfwA5uR7Xun+n
s/0ToJgWETG7xhaUI8IrhaPPOOjAZ6lcYLD67d1rYt9LCEq9I06IgcmrKTHftFv2I2Gyb7L0MYGs
RLhLbSD+yHnplASlh7ecCRTF70rzOb91pf3OEssteg3hqq2nsM39YU5Emt/oAslZaQet1Orhvrpm
qNlk0J91vWO8yJmItmwCu2dI4iAZDBOHTTf1xNQEfJY3/J3i0ly/eN/UmoRxXbnI8LC+R3MgcdP3
Wsauut0//iG5SSPVCSUsA8VVGwFwp6I5bD7mdSY7rY2nCkTbxeP/RHnUo6uZLnQzFvXQpy+UX0Pp
9j216at2r+Pejg/D9rzWP450SbQTtUUD0wmSzVDIlcSQVey0RXpIJEQTB5AFlnaV/Rn75mljzrk0
gQOhaj5lMDnBtUjgKdiBRBeDOyN1aHbxCCpV1RGSn9N+ljMLQ/AV/i3aRCJDAsEuIjFbBuYPgzVa
xtdOWx+F+YGypEJNQ3bKXt6MBsEXzn7UJ7Nl0GykgqX1Rfl0wD9yx4sDyJyB2K56jKmTTcUXYjkQ
UKOmEMy0Rj8y/+o+0R9z0UX03EdAquuIHrMOoQorGF4Fa0cLRd3T4DaraUP21gQXaTagKdR3CXFC
PLgFBgP50PMhndJandZeYkRzP3G+08Bp+mrJztv3+JSIjjTaoKUphFiG8oYvpmOrXLeRA+CWzew0
PjCKpO6/XSPlUZHvPFG+etX008+KdO+5wlHXuTn8kIzk4AILmGr+hHbacTAWxC/7bDgKSwJWYEMc
8I+4DUOR65SmHLpL+LfJPQ8lG67bBwuSZPOaF4SzfXe3lSJA1Pi075XRfy2Cy5hcYJzoVwsgWH9c
GXK+m3xyEuVMGQ631U36G9kahc/Kd8xwufLIjn5ZnM5jR2FZgX28/uWYXoGkklTjsL7eCdFxYsLZ
ImHAnxYM0StA/ASdiUVaOi0SsXp0wfSJPW6zlhnAyPhXzFlxQxC3mh/wHLFfSf+LZzwfopvS3xvJ
l9TTKB/iyxoDQOqawlICm+JDya6ZXI+Naxrhy/2c+CAAKJWvFb/Cz9EtiPhpKBnXQIRsbrR8rLLq
gHolzPe9a6YKsDD0V2QQcyZG2rhAda4o0k8N90nRyrksRUDJzsZh4oJ92yT8lw5gBmmJ5myj8XdS
hHgmiX/MErKHMRcPfssYEZQiqp59nXDuK0gBFNpao5KtV0t6v8hmeLk8xBpK3XuR3Po5lmBcXPHi
M2Fd69esR3YIEu5bbTebVrkfOBuJ6DBh0oWAgu+5fKeDm/gWlMSYPQxKqmLvV5xpLZBMLnjT93Ax
LU/L60atKvbuW5+RAqCUTXnaLHzNqQsXKGBrhZbLPAnVFptZ4za4WU3LPR8oNY/WCClkc42j2b7f
10LY1+Y8Vw4b4L/cHlKL93uylb4uC/RA0mPE2DgpJPAvoRVwCSIyo45LKx8Nj9G1x77dPDtq3PAz
VziaByNjURCUNLqpIYLQXDvwo89w5upXYWWth65BnHweJNoagNgIyzg8IFyVeY4dZLYljqnpDQj/
IwaKLfsholjW3Ea4D1W0wGQrR3MYVx4FxZ/CT+bO9DbE03RGK3sW2k/CT0MAyWzpiwe0BEspFIi+
El448PFcUhkU0dXNGovKyit7SqLnyKpJyeK9YUtmk4stUhWQTZF8MaiQUA+btqYGbLOaV4LI9N3X
U6UqHZL9zgqNFREAw8IdCjKHxwNFA0gR4yKBAlG7Fm9cDMvAzs7jiqivXNo7Q5bDkQ3YAhbDiAh4
htTrBnSf/oKDI8U5mQs3x7j9ZpPljw2yG0k5kUx5dUoApon8DlMo0+0JqGnuldsVItUfk9G/rvIt
SfCohibUghp9JZBoCJyxZjANLlYNpVV5uCWMApjgFNu21Unf0ZeUDYQu1UAd0TUL9yITsiK4tQai
O4rKCjQxfzgqnpklhUtA77NzzvsutqqlH4dGVzvB+7cIzLy4MhFEIGhi0rFde9R3uWlmiwCvZOm/
F+GdQh/FRxIMkjGZORpU++NndzbH9X/eeRp9FiU5x3cJGU6pQILq7gtlgb1GKHhkxqilGSolH75x
D1f8YQHHht7JuVR6Xo4mbZXOy/XjfYcAGbVYFI4Nn4b1s2kQrTYYhKjriVoLFIcjLTEV7Mh4XqUz
ieB+zsMbGPCP/NBEkxD2p4jzbYtMy1/TFt2DCYOsGqEKzqKlKpA8TLPfHgTHfeRIPAfVsVHG+f5b
h9Toqxb9UU6FcSw0tKF6EBybgVbVqDjOBmO4qu3wU5arARE9S04nn0UwUDXaHBrRApnTHE8Zd51E
izs9/KecG/pfFNbcjg9vTTTmYWp+EmxKFl/7BupAkac16/lGN9TSfiB2qk5P5c/N8lyxd5yJWqa+
itkNrTfkwLNPwriK3MYri0H4KhceXdExW279G1uGJZfF7tBoKvftxBqqHr4tfw3cy6J83PWL9e8B
298mAr7gFMfvImPdSgXzsTJz6BXXR2JfjRus1w2JBobBxoXGukj/ygDtCB0hIB0bHyJD+7nWkXCa
mxhdq+n8XR8RrYRHd186igk+BnPsnYrgdhOjbfkqEFF7ELzOSuTW9zV84QE2F7pRw3UUH/sYyIng
/V5zLGhiPdWPR599A90I38F8EPTtCklbenbNCuDiLTEGOoQEQ6Asd8rczdZcA5ci63AWnjiuAyTl
VpH+NEU0lSV+c2PwNO2YM56vq6WRYE3KwlQ5ttBu983iiY6Ib4KPuFQw3efaQ43mTqgUInNbrMZt
zpDM8WXnfv7P1VFxDNDwOGf9mGyxWnxoLpQBsTwDHDUG6h1tdsUeBvZaEFd5qP0lnRpmwKm4GdIF
w1G/UqnQG7JLh0ao/OEf+8SGb4SQVKRdUQFGMB5G1vFwcpRAHE5bwN7ZNbQ/IERwC37ODJQYp5mv
eODi3XAoskzgdNIhkVdWnSh1EPsE1ZRMNr6EXOgGpd58rHWx17waJb8htSII/x+Q2aPLk3xIDCSg
M82lMvWhGUVPa0S45zGRITL1BDTIhsL8yk8+OOfVF2oqNZl/pY1HoN4DFMqenmxo6E9x2ADIhL1w
qzsmiLE2mJGB4grvdAhGi+2MVKZIXfmjhlQXEosa8yJyQGO1liuD3XjEZXETVEJYAKsN2XdxnevF
uvr+o0L3Gsia32I0VI0LpdddMTrKz59ML/gTfmRl385MV4584JnEGGFajtJBYDuTLE4FxDkd4nCx
/Tzd2wr7arimKfzkVZxkhxc6BjojW+hpMziE0v9Co0yVfSC6Db+rnoE5vG2jQTPeEwPe/cBf8ghh
rnFXpheaTNSspbCe1h9eu49fhP4oOuJou+4UkS23UE8T/BG5pfinJ0BGOnteXmPel/L7R5fVjIgx
IFjO/okFeeAKEU0QBLvrFEZr3byXb4J9DjSSE8n5OOOdRvGYC4T8rYoPgxZDkuBsQC/T34Ap+mfK
e144cBb4gTWreaI5TAJn5C83zwbtEXHP8BlfwGJVS/Dr8NuFZi68pmBWQt6T7NurwUnH0ynqQXGS
PYw7XEl5zA0IjqPZbQKSP4HS4LJJTHTp/oDPxE4pTVEMQpudl64N/RRu7uh8tievt4/9xcwX+U6D
UFoBPLRT/OcT8Sn7u6OelmKHBvIbcB3vXqOAyoswQBben0v+yUtM3kUIxK2jb9kr7g6dI58XJ/aQ
vEYFQY4OSRJ9hRu2amzTX1SJcwbq0/PPaphBPIz/aDIfEeGqBkk3khIDEEw3hKiIUXeXL9DnUM8C
y7JB/JiVeUCzgMeo4G032W+W6Pv9Oa5uB/8jG+tcqz5VWDQOHSGxOXkQqaubAzZGy+eUjYrfuZ/5
GJEuj1PXGKt52LyeHGnvhNbHmQPrr1Pgt8yozUgnM1UtJztS3PQeOfPhB85G41hxqnz7IfSrFBc7
NviMyoLg6QJI/7zRc75M8LfqbZuE54zlJGrvFLsQ8jDyc/a1rFt5SB6wVYLbFLi2EdBTXhFAkc7G
vuh3lPP+cMTHHz5rK8f61Z1+GsgkoxDR4JabMJg/a66GVLJ8WMUnwRom18+bnEN6noCCdrdVtsDt
calon4OY1umrIh9TXeFSvKFvY8eFDBOWoPtvVXaWWO+zqBs30iCm4vXpu83bQQ3LKJ6TCt++gloZ
B1UOiRcvqbznizXVzC6DqsL+F6P7E0iJkyBvVd0FsxomcUJBl1HgktIV82j70iMdqfKYS4dkHv5N
PgtRRycfCE0czezs0LvFzXYHlCOHJQSESh42z3KPhUMCe0aBp30cROUZxiy2/TZ8GF3ja40jmOvo
8M2xGbi3pDkNZjP0lLuZt5hhwa0yTK0pXdDdqcAPv8jL+XFtTZ324HS5d/xxI/ZYudiV8hS9Va/h
A8fGwGLFbH6VTFfFuH48wDij9myHOtILMflV5NLilkTY1Tbyv/G7EffOHlAsx4HKq/RpIGUoh3fi
sPokPXHlFl2NNw0St0fpX3vAaXX9ItIiTUOv6Zl6DrVZ5IRJdFhObvN3EgMmEEmgN1Z7yPW0S3hP
52lvWLyP/annQIobNTAw2JgMeaDiacpP4LPRuNVHUTeYkmGoRO5b8CQLbeXW0QouKiFwUysmlOIZ
pI1ERgzoNZKTQPHTYhFGU4O82lQ/DIGqvGzope7brGdD6H0wZS9hwTE6+iYfEUIpuJlm8iIFS07G
hIQfgks8jtRcN0rydBqF39DtJbY/PdJX5cFYLnoOlhpPhGb/838WpJQfv34/uGlvjmXzS2Swzj/O
Qb6xs51nJzzGe/eMyuQ3pbn54b5CD31a+FIqkSUhd4axXmMDQHi6zBGXCyk9ADNA3PaqQSlK5566
FgOg5Lk5KHrPuozpiOSYraPyCRbelH1AHIAlEJiK1JQ+bm5+lA13T96fNf+z/2K/77i3FntuqCuO
IAk9TF4K95RqzvltE3T2mWkNf1HbzljQboKGReawtcaljnkuNMVmSu0VFrqX10uusK1Cvaryjdwx
CT4r8/J+WQqXr4x1N54zW/skeKZGfl2nFtgfQKSjAjtwXHRqL+BirFQJ6lOi9AjhmiR+lLc2SEQ8
/SvXpSXsWtzfP4XhRnejOgtgWTYxKIpP3HfS3h07uQiQIWV+OHauxECPfRgRmNgSYDLR6KGhgcUh
LHlJt7GhPe0W0J8sgjkubbCcffXxV1QEIX7nNItd93FGRITRd7pHOYk7hl+guMPHaAf1vsOwVkuV
TExhvfwLTyrcm9/hyP0LaEDCHThTTHBukH+SpuAnObumzthSUIEQ1zFf0IBfxxeP74V7H6Se/Tt7
SFB5eozEKnd8WmiRAo0iWCTkBRlDNW3KHOk3nYFwWE0udTDs/5TJxhllyhkISa5jEmC6Tq+qgPTQ
2kwIeoIO+/fviJnPCJ+aIpkoJQMVdAnsJtbL2CAHP+iNxLTMFqmT/jmZjX9OczEdf5zwyFsxaeYQ
e5aFQ9G22OJQ1J0qWGSl5Bi8kF8HHl4uQ4e7JL0lwpb4keoNi6UBlnuaZFzxTD/lckxZB45QERqi
HzLvmE9AJiZCi8JRw/LT0giYSOWbLVJ8bVxsqaUFxqqML7kTSCmlI2bQdBXc54I7Tv0oerY9SlVc
D9sYjhtLfXh+Tc/28pWt1CLgG0jko2tu20GEM/LK4/Da7tpDYr9sgSMk9V/8YHhb4H0f6UEbBz+D
rYU1rhSJaoC7BN9Aq2rpdxpruZtFllzlGv083cR57/DbCuTFHL/nflXC1VvCj/C/ZpEF/S5+dhbS
qvSRTWpzepD6y/IkW55F6zb2KXobZm5peuotuTwrLMlfGR/v+OnKUe/h5QnDHPm7xUTUJ55XtHCa
Im4FJ5eDoDrmtDNSzLcyWsj234XXNEtqkrrkQ5CuhUzTQP4cfbf43MUlrMVefWZursWeAKNt11cP
J8aKpWpq7x7yBbMMHEplSpbOFZvvQOvsNgUxAO7P/9sDsBkQFOquJosxbsSHw96GaLFqWDI2oM8S
n5/gxSK1KIw5uDC+H6KFF6fsRUK/y4hBRjNc+aDfLZCkYFo7rcANPrGo27nX9Dd5ey/R0VXOHxzw
G8XpDW/lzqkfnIBr64/U+10iF12apiRCnMcltAClqt1F2tVoiOlqPKjAbleeBjnXj04T8NeP80ou
xB2aF16UDRtpF+qvvG6D67OFpjg66UdMa5Z7Ktf8SaWU0+5kil97FWcSWIDIO+51hRJ5tlFUakui
+hD3xNMMTQQ/0quRGercknnXapLvVBaI/ijPxbJsWyg23PZYWioAQr9cTsjLTaqU8EgOwEK9zwoj
eTDHn798VbXapbYz9LANR6VaNTs/fF+7UoXSpCufiheEz9dZNRt9aXITzNFANk3aMoIDRZoowH/h
ZdJtyYPEKPZU7tNDNzaZ9G+9owCfuda7VWAMQ2CpImzd87dqsH0S3PIBa74Fae2cRyoGZA8KmPQI
ObF4YkAOkJr75Pxyo/qD6OIlWLzUYXi8n3AAQMACu7gMRsV/+88GrXCs5Hlom8XZ7FqxboC3sgf3
ycCU7XyZus5M0luwd2SktlM93+/C5a5tGVkyZFeit5Zudmmle+KGG5TPi4kOpm334/Vkakmx4pSC
sc/8iwzJwuyoEPu22uCwWlpEV7XhG1SlHl5ApOKT+Ez9l+D4p4S4VI+EPSfwU0VDbHUJtGPnwba1
+Hiv1BauHX2c1O9XPJW0PYFkkUZ61wH+nyfsOAdCJ0juhtRVxjgHVNFkQuRwP/NUBoXKbIieLQay
6EDVJpdWeABJT2p14Vprn80kdo+eavSAFIfKU1YFqGhjvEA/XYQjTPD2jkTVgIPzeLhH0KrLNGZ/
6KZeXHcDarY78E9/jxFobBZThybUU7/ddAh4Qba6xOeZB6IWS4cpvHFEQCsVjy6r9Q46FqLr5Pad
AlJN6wfUoyEfy/wDCGlaY8j4Y0ns63894tKgziVj5faR1zErvtznpkPPbMf3WmMJJF1OYQQFiR5I
pvDNiX1b68V5obnNwJzNDlZukRn/Wtats/snTiluTqP42Wqv2A0b39gSrkbg68HbxnTSV3nBcua7
O9wwVIOjEGXpShX1Lx1rTklDxIY3XmSyi8X+O4zUutuoojivT1Qwti9HE3b3UojZDDnN4QTA3lY7
9PfKsyFF6MSnaLvwS621C8e5Rnj9bWSGXfQtk+BPUu70XyYMnYiq1b4z47CiTnnqM71Z4CabyWqc
mgyAj45r5/zxjmhrYvBEUxJoCmHIN/2Bga2O2xVSX2l8KI/hOa74AIo6BAo+BaAKnBj8Ykr3LvdH
f5S94xTHpAKoU9gTf/AYAPq1x8mrGihBsmc7v0mMFJqjcvd5Sy2OiZv2BADNsCr5KcZ7WLk0FeyQ
tR0hpNRa6reK9iCcM/B2e6hZ1BjdZ9JQklxQO8EPHbgKoyvd1nhSh4xWHJFMv651QyPjIK2tsjRX
DhZSKyG27/vtMNb0vG5usm7d7LebHi5X/T3/zSO+wIS+ZIQmkUdnXC0/tu42KUcddHuNi/pK8rjJ
x0JGruUuPfOiDs14ZvVifzdPnTq/WqVYnlpnwr1d2H3O8E+LEy2IJRKNV1mLr3PRCtmx7UnmTq+a
VI07UvY/Soa1kI5zWBqI6LRveMR2nIvZh5ecuBxoAJSIhR+i/OP7I9/FPFG4D6IhjmDZa7oFqw5X
R5vnMs+MvnRudnKCymJbThzNeQzGu98RJ3llBBb8zZyDbVd3nnXMKzPgWlVrWd6KrICbcYV93xWR
pKx6Nq8Pecp80iqOba/K+bRmYZnwq+owMmkbdrITb+z6A3CAKEwsL12uvC5i1jdOlf+lRMX8u5/6
dkCVe3Eousg2JiP4Y82YC5eB1jJKxtJEtxVdi6Z9FbAnrixQjKpmzMrvPdeBmXjmxc1WsOfbZPlt
Iff+QPTosIK0E3R3HYdN7RDHLlqiy4df9z9gCSVxA40uCTRPzUvW7rqMUzTJfzYyVOCq99VCh13S
xNMLj10FUcr5p8K//ZLmqz65T25AqP5fl8LFneRq9bC1/ugE2XTAqnoCP+zJ3i02BP2hKz0+N52g
8Y4aJoZLk9sUgdmreNSq4hHsjQxmZxenaNb8wmAU07IqszvXDXn7gpcFQo6JtmarNKrtu3ZU9hev
cYMjwqrwQ5w/xJA5GOp1gouVtdc7SN5EcqbIMElaCJuFhtcoFnCH6VIBSmLJoS/eYW1SAyQonnsh
tyjQIEAhSAVZzR6rvcHRacQQxNpR9soMApW6nL95mM1mdMzOjP+TTc7mhvv65mcFmFfBoMOwNVJL
4/cHS/BOGv1WydMHFdEXG+XW3dBghZTm8yFFG1JKkeJJD/p4T6eOxf16W07y1rCavAxDlnRPSyyH
weOYTNq45VgqqZ2DCCXyDRKkC2416unL1WOu8sa+Ad+p7GDXBbeFGsf+pin11O0YUbH4AoJClROr
X6YUZAfsLe/zmrr4pcWv5K6hKxC9Gyywg3TDdb9Hso45+Do6z3mSJpejpdq7EiQfpR46mEVqUS7K
AI2+BXwS49mTMzz/fIEeqgW698rek0Vhum0Ct5+ov6fBmCPvmdC94AQJIRArc9Xd36pHzHcyxx0h
wRHl2Fx3rGA1A4/hSj5t5p8+sJcqcdhC7Z324l8eft5mi/Er9dY5Gwgw/ge8tCo3KBym9BztsxAi
LvSp1Ahv1sBkMxi5Zr1jcaO+GTCDN5wFxQbdC1ywI87nhU827z6twhy/GSbSPxiMYZxtC7FDcBBb
FYBuQ8ydp7BrW5q3weueneoLjO/j1ty+lAuuXKU1mc3Pvm+S1Q7w31C7rUOwh3//+14/M6zoLzeX
Jd9VR+aEVn/g+SAg1TvwR2YAJLqOiBaV/ncM4cC4zdhRa29ub2tMnDTCO3Fm7+FNCVd1Y7GQUIvS
rw/oqDrqBrWIIxkCsHx1vMDlKE7Auq0azz2ivevXYnpjS7Yr9njgmIepsGbL/uKke4sGkjE2vBCJ
cpzb6x2XDd7+p7WeYfRHLVjnY3nG2zkBA7fyqr2+98MB18+9slcaK2DAFtHRaLrjyY7d35tcH+l5
sFjjlTwvrKP7qF978qwJRTxVK5JQMGKcoloflWFGa3LF/wKwCxRnNJJQWes13W+ycNYf4z93SsQk
4/hoX7wx0N5ES/4bvukc7d3uZyXhw1hlPIDcqolCwT2avP7hMoLFPLbccEfBwiHWsbDEOHZZJcZt
U5OmijMaiHL6aILBEvxHrJt8PFrSHwXM9c9cLdludk5+MlagO7qGzTu5BDZlFvDiOu8bj5Sv3Rph
g1ZzL0g3bsMk7cZmlSaMz4Eyb71zJkwHhSjariIyNmV7kClkEzw6VRu1R99CZNy9dq9hs4CuArm/
drZqc6S4sdaQ1yJGArkreaHbeI7BYt1HdQ9er7sbZa9/7GF/lMphWr88lQvU0Ec10W9NI0c0UjIB
2Pw9p+gBuL+kBrljUYMEmWezJQ3nwlHKzSGnOsHGE4lVunDTXQQySEZpPqZ1R6nBs5omOz1xhQid
1li9Yq5vPzwhv23O8bjWYz6e8tWr2jBCQqa3T9IlUoc2K5I5J3h6KXBXK2uCP2YXFJ/T0LurPRU8
QcmkKxAcfwiOB/iSV6Fa17ywb3+7UktjEAANclMcQj1fWe3D6ZDfvBrrGLmxTWK13VbQ6pCLZ+Rd
hj2N076Mc92zDO3Yvi22dbrOVZ/Shh1R+RQZBDqDKX+6vp87JtrmVvQdnI2lkRl2gEWC5VrYTb8+
UFC0UErGXp/SzUq3fSh/vYgKaQ4Bt/vsm1jDv+FV+K/Irj+sDF8ot/jXVwBw7RkSaK4omE3Lss9M
0MPJ1t6+mqHXXknBRZ1Rfe70BA9sxbA2yT6ivaNgTw2xa4FMVk+ChZNIoA5ZASgZ4UcBhW0ZLAw+
acUoM/Dz1cYCWa0TNnFPaJdBeXnsu089SXr/UC0YDeUrusIzS6gj8CrSf9TDuQhvkePm1NQSMC01
O3h9Nx+DrzJK8QC6zT07IRxgxcRAcFuPEkMJKjngf6rRkalFC1pJUgdFK27Spvm3DPAgR+cd8v3k
MPJe9BqSKQlOxU2m2HeAzqhyzXCBFlphLi2wZIVGQUcsUdIyMgcUrfsZ2BmBx4AOA13ky/G6NMRi
n8T/MapGYt/nPk81dAU1cqTqUR/q6O+NOtmSR5XwoU1XWkhWXROPKWnbWho+7UHXSvLZBiJMmIxl
/BMlPs0qP12SteG+914PkiUaBNon1r3jmbq/I5pGogpx12IlvLMfW8VJqP6TWODMfs6d81sWW5+c
DPgKfBzw2frWFAPex7i9vHT8U2MDZ21rESCgYnN+Lm51AURRbudX1qA2ZNriumlpVe5wNTmgS7+y
AFU5E6RdppYK532a0HgXzsG8hfhn/2aUyyuwtQkBI1ONttCitZFzLwUM+yiXEKz7hfWA1S8FYYhS
dzHFE191Gwj+0XFzpyFTdoJm5UhWfarQ43BE9wb5aekdMzyPtY473eWR9YTgt09gRIHcVroreBp4
3VzAECM3GQ14E0+2pi0Ok9tzj5gXwRoUb7e0frnjKrZzQ6sO5IAtx4ZJEauRdyGKXIiWfC3pjc3C
x2TfIgEyljvY2ZxcxkpKhj62w1M9AUQTqfYIkoqILbX/+UhFhn+HIjBYltwUbKA0u7aW2XSHQ9rK
usT44mS2tUkmXpkuY0/4uZTXEKYQzHk0XcW+9z/A/WBHXBc+BETBRbAMgAFhOyG61W7qKmDrbnmv
R3FQb5clp15UuqokOCEDlAw81Obb39ylVD1DlDga2N5UUEg6Uak/Ryhi9HGUU30q4/hpgWPeCeQY
pr20ulpZU5vfqq+CNbggist0vPkH4wjL5Rop/o2QNibLMGEjJJ4w2S0+bTwGTsCG7mcKXe7+AMte
F3tKKHd0X+von2VbmIN/Zlkp28lENkh22vMTx2q0xKjfnUTFOPSXgY02Vs0oXXNcNYTCupsjnCE6
5XMaiyk8kCiJGbLKv4MYc7Hv4ClZGH2onkOSI6fFxSKRYyZcJdg8aKbotvobBTjATEomDNPMmFk/
bPpoQDprPnxVPvxEdzGuXNLypb9U/ECbdBmoVpFsTcTjeBGdSyxI7Mzveul+0m2llL+dtIbQQmtz
TbBxR+aZlKM7bupGLE7lChfMFoudu909Uw73bVLaXE0sHLHNC+7+il6kDhz4T0er4U6NlJ41Y8yc
dsEzNYJAtAibQgDXtcKGPrc7EGOLNXiaMY4FUFTLduFsKexf71lOyyF3X0Ger6NA0F35ingU101Z
ZW8sONu/iVZtUcAhrHHQsWrF/GvjjtL3LuZFkWjTVO4QsPn37mecp+tRzUOs4iKMIfdf1qOzwRic
lJWtexx59Jb5g4fGQRbiMS5KXZCzea/qZhvqWiLJfgTQ2A/WCort0qB97HVKsa7cp9waT3IoxvEd
DV9VbsAwNax3/7Dp2x4gXwFTBxuno9hXShusSLmaWL0fVgQZS9Bvv3s2TcVd887tEUE3uHazzJMr
MQfk5qh9Y97WXdD5i9gbqzlvdfRKD2p/4aJGpYvvb9M2ZtsdUUkIvoJY55BViwZvfPNrw+0JFila
Lhitvg4DuHDSGD4ZREtE1sYKIGF+BX59E382OKZDrtZliE/p063dfULbXsjsX9DTL4Geq9bXmBTG
7Ocju7ubxpJMHbvCS72y1m4H4M9/4MkDMMPGbDap63lZ60fLzzefF6bgQEDSntNVbqerZVouYP/G
7uSfUcbr+luYq2q0H7qzb5PNJ+McFAd9JMfFQ08I05oNoBPHyNg4vRs6CONYjGJPqa3Sm5YxNhO2
syhFYSeYnxjvqCVuk8MqxJGOIU2jVvnVUO2NtMqmWkyzSUJ/cAx9jLS12XHmwrz2Cv1HvT6tpNDJ
5eYAPJp6+m876htm1xEwi28FgUh6yPvCBIiH1/6InqFiCvpx6upibbq7zGldPFfZv3qhdpxOyMlM
1Z38BS16cDZCX1NOS+5z1ve4nRdNRW0DNFGIgriuc5AgBELwrrkQYpz6SMoKQJaajxQSarIU+ySc
FqO8f7xaTBVl3EJAf0sRophsA/NKggaMBazatqwVCOMSu8AujYKefDHh9aDgjve6hqGAgttMuJpc
nEhgh6JZUV85pfGLHESneWCUzeY5sKnO4cZJKMJCJgx0YomX1RuLtZU4M50qqenuxuMzphxz2N1N
IlYsMJSn3aXurmoKhD9boJD4cP0f9C7bRlJqHa9QVKIaB1+1XE6Ao7fTiPTSEOw0rV9UyxoTtNXv
o38QeHdEA0BFKT/nFSdkJN4eQSDmp5eZmX/crpx2a3kgttbHubzhoLWrUCdncn5985aIKGRn0q19
yJ65Y0dc1E59D9MgoDg2McKzooQ21hQSp9F02wTDoBqQawLWky487/6PIIws3FdUg8iaITe/x1YU
/97G/3xwvle7tCzyoiDR/hzQndnXniNQ3SeKuOLEDQkAnOWnnZ+pY6YMbyF6LSN8CH5qAzG4K6eT
Zn963n1G6/Lh919bhH6lOqztoObI2dqKfY+pd1kh+xLSo3ndDVQLFpAT8Jt0/zDEkOvZ4yCmCrUa
O7R6T+rHUSFwENrgh7DWTwH2T+pso34UVM2xaZWe9dHs6SFdC8p+Lq+dny6MtE6b4Q5mVYIxVt0S
t1uT/tatVDQRpzyGgwvBygpyeu1V6XDQfQyt0/MiacHk+34Np6hQVCCsL+chK1UeRkCd/6VqPixM
gAxaNQ3BXQO4S6RKUu2w6fKT5DIzq6BfQ8iXwgeYrh2hnbs9GJZY+L8YpilF29bbPTvPbI/xPCWF
hrX2Rsld8GrJ6fWhiA4xfRz2p3PyHe81a74hWMqN4Liyyt35vE2MmcvDplh7H6lrfjQs1r7gKSIW
QtBn1yNudrA6Vxgyrf0by2/8l7S5chq6zdyfdh0O4iNpUN+x7uj/d0TSDIuY+7bBlbWYQQuW0COD
sw+ZlzXcW383/MrEDekD2fHc3ws58w6ETZEounU24LsC6aCTQD/2RKc0uEr3Q4NkepGCfwyZEzZK
7IqLieuv4c/w4BKb/NR+BIXLsVsP+q86Rv2i6TeBAEz054slMT9uOXWjf6/OMS50OKal/0Q9b6FX
Re8zcEpg9RrHswoSqMf65V4E36nv7OF7/36b8OM8F3RdBI0xnaX3KEgIwGUqnLhNinKaBWJh8nqc
vFUe2fbOQh043gbcaWMEiQULh8yPttNgpwqixBq85tjRMG15qWZEsnsnMiryEeUp0omocxGR8Qy+
JeOWT0Zf5nX07zgDs2MSsrRt2TtQyjoSpqBa1t9OqXgb3aSTYa5fNTezzdbpB/PkcJQlAE1YV0fc
YR6pLeMXInNa6+yxJ/IIQ5B+lZ4A0uJM0bxLpMDEVZ0JPF4BGaWvGhcWEEMD8KfymB9kAfsiqh0I
VocPsQ/INPRTvbw0o6c173Jra2mHJF7T99MFnD7hQic727/QsjasHKJHQRWuNsg9jzZmObiQhovu
PRnpG0I+DsYSdgOnzvwLy6jJU/Jd5TqYt5szWgzaKlBzZd7QguncjMIKQfmPAUqaV5ElAecRrl8K
f75faLLrIGNVVUnHWYG5MQsZgT4UzW/UuhuRR62+IS/xLcW8IIfa2Ew4KjzyeHksihPNbU+QPcnf
3dQXaDhb/wPUX2OS7NwbaTQ35GivGLl1LnSUDGy9eBAmSIMWzMcAGLGQ2DdvrpJb+QMRnrS2oSWl
y5+CTpX3KNapGfENQ2tXhUk8MX/xPrB7xBtkWtI7w6i1GqtFpIjYsGTGUqQNderaGNmEZh73eL1m
p47Fr5UUXafmAxAIMvzT+c1zTjrTbnFR2s5kEPtVXmwS3s93jJSV3hmCPAfglvRbz+TMd7ZIN8Ri
oamXAQFOVanqwXM/zVo2O93Dgdn78ICdsow1cRFf/e9Tbl6qCl/kbugnzGzLgNMHeO2zUp13cPmR
AuEEWIn1+h1vFhfrCBz3vVlOOXs++u4PxDG0frIGyz5FAbFKV9LlOys5XMpj6R1S49D9HrNpm8ol
nmz8SUXhfmWuon86Ezsy6e3Xah7475eEsYLIOlSBP0+htb7QtztCkDVfe/fq0PuEoRfxh7gmlUr9
kyNi+Xen7HIMDT0zkPAq/D8D77ub6t1IIdE74c15htIrqNypWMOlDJ2tZKpRGJP2ghWCiIw2q1n4
eHGgwQhCeTe9I2s8yPYl2eawc2heyzbQ5xnyqu3baLlIK48jOOg09xJIBHIQh43lswtibDsuFKyS
AR59RDsHRWYSlt28wnjuJN+M7KbjnzjecAw+Bw1Cwz8YNirjQArPzMS2uluiQJb1AQw9utfhFvB1
j8j/jeI0iaFJLAG+OSbpdgtjLOiKqwX6Z6+Ai/rQyvaXLJeBe1cESvVU05hSPsDpPVLpspSQ8xdD
MZGGkGork7yutjSvZzSGNBlzJMcccstFPlto0kAlgVHlLPEmX5SCn5y1MjESSLYgDMkk6xVXju2I
YR572XJUXYsjcw8aAY8jwFlIb9YTMb0/O8kGu6wSKsqMMPTScCJ9SZptMozspBn9It8wdeI57y84
sOAE/F/XpMy72rISXpntM+J/NqS78jIGJbLwa8W6o+jgZigaAtkaUxgeQcQbbt8DkhKNPvvYo636
5MJpH4ugSs0YVq4bPnigGs5o3zkaqjbGCVZzNB8QQjZyWMFEqGEZ+I/SdxNKSwi4IOmb1gk99LI+
tli7fP6ab2soPZtcBkMiyhaaIbhHpzRMg7Nyer3Wd35vjB4vjob4KaU0ajKZAMToftLe3N7awuWa
ATJAoqULfW3aVRSICzsSI+GKVX4InYBWrEhO/G1+fV+5UlwCkSXY/CmFzaFxyun2v/xM3u4PWdg/
27bFVny3MEal/pMBi6kLeJ99odJCyycWsb4DugnXK4Om6C/VyRzkjc/D5OKNU1j5jL8G+cGqKCta
aVmmJZrWxO00a1ulAOckOv12BlIX8QuXIZf0ikHdCbXbrr28ZBDiLettyHhGJE029ud2qzqW/B6K
lacWPloV06ESX8JlCv8XTMbVtzXRbWGUp75XetdkFN5uvD6p7DUyojZ8w6lOlzO/wR6gT0WX/QBw
Hv9uE8Nd1OZDzyvLAMlz5/A2JPEi8DF0JBF+7KTgR5N10fhoOVApzSOgb7HPDWg+wnDB9Gf990qj
PvgM5JVI7N6b2xi0CnCBoefHesJ7ix+e+YzNW9Wk2DPOnkiHErqPRpQQLGg2lxFlaxAUr1BACfNi
y4CfnLDEJ371DWatnM8vzO/hbONPn6iCEL9wFii0O8o/Plg9EQ/D5SIiujBf1J4DXbYtjftuNZoU
kfdHa8eHBLoyZniuea+rBxueXHVx3rM/f/ELKqAOkL0h5xQb2upDxu17iOS5nvFPSqJx+JBhRiGX
xcQyMNmw+9hE4OB8zpN2fRMK3uOJh2xAdUY83UVYPiAfYCDJ2pYi/778RW+98W7v3U9go8Y3uu8h
RjnncmH4s2C7rYHmyr/8tHB63tF+f/yH1j1p2TjZzr0KNCaFd+1vMhn/57ofWSw5feSE5ci42ARa
AQ6y9xsBOzx31FQcKfLKB8rbd+Cd2NN6VG5os4sqMohL1xiWiQUViaBUTdEe2bTADl5bK9C7qa7J
uhvAx2d6+IkSJRah8Hg0Q0QYc8uJG85APbHw/XIHGhJETyi6LAA8K7J/YcxgDp68Q5hWlgLf1Iho
drJ+qLFp+SNxXzYFBbWXHOvHUoKPCivHXOk6V5Gbv4vV+BFeJDESjvF1WplN2JsuDdjsYQA1bhmY
HyXO+5LxvcHU51u4xk3xvTp0daV9SX3bS/VtqYv1mFVzHugrRDQe7vUEm7XJJDoS+W5kIfoUmj1+
NBtukqvm/wrlazBw9msRWKh0KsT+8NyZW5CKkHR59xhSxtWAdSQp9+jN5wB3wR+VTbxnDPcm9NdF
R7JO323RxCzdkHHk1d/zBCqOCRWBMqtUBfWYkXIzAAOENN5bG1/71RhoVIK7SAyLDmNkhCkIBeh6
Wa36Yr8Q9EVHEcN1imPhX9jNfjcn+fr0d4LKfavYumhWWzmMVsCO1M9nCRIch3G4/aKqJUELeQVj
sE/RZWoVih9tNOOcy13VnZN6QqpIwbN0kYHP+NlKqsqF/qj+ms6wHVsjifU560gIzeyhEt5Ja5Nl
OH2zp0tFQ45ynW/Dtl0Cw112ADFvnYu4TgJNntugXPg2zix4g7T0pc50WSFPXMm4tdu3NVrcnA1J
gcj1bddi/CFvityo4Ce2GkY51K0WYojv5GyO1VH3Ep22Z5i9EQIaYGAg1EEq1TGuyEiUN0wfFwGZ
AxtuKrUbKDMBMRArpwmNPH+YUYshLWkfikY7hUC9EasFPG8uIz4J+Uozvifiy9aXXdKs2vgjEPm+
C1+dMa3XfgXkqobAGRn9uFTLJu7SOIcS1peTYDQQtH8cOW8kGNz0pN8YVIQ2piXr//7VOytbvRg7
0FGlQiBXERYs2cVGZDzwy+4RP/01jtucf8vG16PYHPzSmJGDtfNRc6LjfHgdHgICqq9ZpYYrjysx
MFK+7GCLelLCZsvIYS9MioGcyK0OcxKA4wPE8fUePUNS8RyY4vPmvly0oPbjtuyhn9DFPl4WghqH
fC9Y9R/ftREHCtfwN2sXb0PurjW6U2MADiyl5mgwU+hS3SpZlLPETjCDNynXuC41o6SfIXHlQtd1
nIYCGtWrOWr4VG8Ufl8rmzuusBzhPi/g1ewVy5BsbfM4z/KCi8ADsuan4K9coTkhWGDwt0OdNlkQ
mR0U4yGrREygShPGHdQY9WyI8yeZCoxSDCY05pLrSDHKKKpLkmOKyIDWmE+Nm/untUrIzjSNpdrR
JZ/HJ7186nego7FPlHdTRs90dv5l6T8Z5LBsQmP4gscMnVrbWrY1/If5PkS1a7+5hRa9fMq/djjf
Rc1beWl1YNARAWEJbB9HVJIDlwqf6TE51WI0euxINfy4qmo7ICPRO/b6sG5tTwssP+V1jWcbADk0
OAyT5GKN5jd4qN3Hel9vM6nKTeWw7Pu40ClzKma3xu0koiGClqZosUoO8Gw0tTkukEeGc/XyMuoE
bIozxRRw7mTkUZoIuEWdGTnP0vjTlKCO8antjfPh8sLrNBQss/bsamk3XUji6XxWAWNT0Nw1Vv98
zY6Vg930YY3IbRFtZmtx2KkuktL+zHwZFiH7oNQlDiAbwt1JjVxUVH366I0x/Spu+i1sVPaKBKm7
IJIM1AEMJz8w7E+8yQ7Qb8byPEPG3AZL8jkVuMPSV0NsrIwEkxQDqjQtkA3Cxaf80rFvJTEw+xot
h9KMty/uUcThIMn1reVUGT+rKe4PpjWi2t5Y0ji+ob676EWUiHcdC6wJGNIMB4lmUIe57Zl6GDtY
T6LQqYRWlos76Sj2Z/FyEa3sg5sAHyQ5lEn2oTUINYeNb/zVHGEIS4FP+LiZ8QPFAyr6x3xOq/XM
KA2k8bSHJdOQrhNZuDqj6xHzL5ZaZt6dkyiI6+uXqCrPPeV12N2/0Wr0cux4ff76PpnHVvS1XTZx
wqkod4LB90UXpYealmhfeeJTVU+585Hppt0EAlD6OS4fkTd8CFjtbwhZn5qAlcJzf7FUjRX8rpP0
2xS6yfsM3aLrPrg2T6R9CysgsgXhaZaEMro43MBh0xHbspsgAcHOYWWGdxLFFNmXHA2XmL3RrZt5
zmo5xkH88q6sY18PUk9SQEpYBNLl9OmfRwGILJsNUQNokb2uR3Bl1E5pvp/njzV1vyq0Yl6cK9G2
yPV/ju5b0C+eOmZqX2gFfTLH4eK8qsX8ZGEExTz/vUUS0fkp+gzqsXy7uTJlzQaJ7H7ZQWGQNTha
G6vjbQVnLDWcLjl4ccU+mOR9Dy4dajXOcHYHKXpiKblQt5VJ4DV47cjDycQlvsIJQEdK8kelNL5+
5Js86GpHe/0crIDsdDMWrNG1KyLICQjVwVuDRO3fC1hLpfWJzfiQhe7rRmDIGTJXIRPL18NFHgRM
Ex7bF0xztdagaLOfK/WAYBBvZcAD/4RkuYEFCBDGfIyWQhT+ZLmJqKloWMmIsFvYjuqBX5Li3FVh
m4c+UN1iqWU3AklAS44jZzZDeb+H3iEKiliKRI8rWhSwU41PzlFnHDB863CpnEkBGbOBZTVggxMs
a04gtHEOPEXPdtFWx8uLPkxJRfLeo4zKVieBoUCkn4hj1AWNoUc3wm1tXepjhZX4EJewB7rFR7nw
T+4DdQF6bJ8aznG6QadjyoQFerJqHNVheG4Q0+7sBWS8RM0r9VaSRSoUeZAk8P8l7hZ3BZ6jjiKJ
WwEYrmui40PKZWt/FEhpBcILoxeMM5YFhQKPv1QvrnJIk9BoZcYXOFohhxuDrWLJOTu6T4IOKXPJ
agQpa9zSwQncFanV6Y/Atdb8+c0VtBNcsLFwUpNDroN3sb/XeRMY41iRoisOxusNm+lxFS6pyH9G
d9/SdU6fJLGXTSveqL5I22Ynt8TtuRFUtp8UjWbNA+HPmC1UdQ0o+z7wjmMnb5mIFLA1ZP7Sp8pU
ZLnxuQGXhLwaH3rKfMPF6B48VZepgdFdQ8YNlh4l+BdOfYkQn2qlnaVTCK1/LBmld9XNFOSqJ4ZF
T3VlYc5VQw9wni2f8LigA/jLclE1NPJiJ1c6whkscuomkK/8gDgiNbLPED6Gyj2DZK9/srcyM8gM
EFXS70XYTBZlKRUvAspEeyf+GOi4bIuo1BdMwBUpA7j5AI1ZQVcUJS81LUw38vnsf7DcAqWkpLWl
Q222QalFhKKmq0/HLh6a9YBEs1yvudIyLBK4b2nau8PeIS8bsvrJoOLffcAIaFYxvmR+vjlEpQRY
64VyGeYHxtTAtwhb+Zi84HcyiYdks/mGC/m4jE4xXWgKGOpGrbSfCxNH19H1QDZPx9y/xOpJev1d
8ncYMLs83gMBPkdfGAyng+4/7U3LsJHf3JffQxyVRKVmCXXco3hthWRp8uFHcRcCy/v4o953csfX
ygClhgAOGsWpjx01d/m+LKs0vrSTV/S7/4mqSvcErz4eGW+G5ghOLm76v7kGOtS14ulP5qJNvY4G
vGR8iZP0iJLPRGXYMeGPAf4y4WIDHT+6kSYcYb84qfgaCUef7I2JO9THHhG+8o5TszbR6C6tNY4M
STYGO4YaF9pwOys/JRiZBxKRI+eHFvgLTf2A8/Nc7wSBbPhDbkwWc/UtD0nghTlauvbl3RYytZVy
khrRRcpTd2WyqSkdKOEBZDgvtRQ5807/NDyBjhry3IF02vkymytwOpjcu+MQIHsDJVh4D+L2zkSo
2DFpPRUfnH6ql9VnDIQq8Ejcxf5H2osdXFHcpdhjuKceP8KjjL7LcHQCJgp1juvtnrc58wpWZZOx
URtcf4NvKmd0w7mUYtbFnKWJi9eTWDRW+6ppY3xsm4/IXThJjX6t2L1MQHtozsCzSdcUzTFgf3We
f7TVzlbLaGq0FwJG+e0bB/3fY8vCQvZvrLH241BOBmX5x8JmkXvjEwqF8mH2eH/V7oT0CAikO06P
NvS90iijsbQ8Cx+MaKx5pP3qzH8sF9LkduKjIJxt5HSske4jcWdKxTTUfJeM/HAXps4hMX9al2zB
ELRbWoN5y3d4eLA40Fu/dNOyyKpjU0y3g0j/4Scngwk/fgI49Zq899S0ZPd2IQ6VZ17aLat/C4TJ
mj8b4jqfUX6mNzva47wwC4XPB7eOFhmrIwLDk4w04p7IbJegn6zlwLxkKl9ypp6ta6I6bgUdTsB5
yXXQ3CjRc+lnFpoV1xxWe9674SH3AGzbSxF8PG/HzocvDg7FcJ2zB7m3qrtV/Q5ebWXCG9JWNKYW
2nOHmvfrkT4GvaQsLI0ZYIJLFvV6nwUr0hvvq57lR9TX5I42v5ne8hNJj7TolN2D274aFUpyiocz
tDBLQ+0CEmlCcmSXVd5bI6E7scolmw2S9iCvTi4FZvlQzdf+ceGOp6VGmT7BYtgGRIy9Ok2FjKu/
hxgqJ0VjWlDorAnrOy6rPWAtORah23LH+ZoPcRCpfMD89EgGdBwWwHuCdChk3jG30ESF5oizVPXf
vEgYodkrcKmOjvrMZlEKOJSaJCJg7BCv3CqdZvsjQOOtlgj5E+7yq6ZtGVO95jPiZsUtZ3aynB99
C11wnPvN617fzgkhCoablakhphv7RwORBPaP3F9MvD6S5q1yCH90BwTMmoNhM2xLEdxIlSBh2IiJ
tXipKJQoKLWUqgipjnZGqbH/8bH9cTUbGZa+GtADqCmAVIuP8YyHBAh2VndCj0gCWdxVmzIynWUi
6473QHoA3bW74hDeiTYHg0I8Q4ZEig78o0nHeyYukj4Lc/tcYT+lLLHJn/E5eVX35kvNqtDCoznt
jcx066teM7lFUC33sEr5iwg3nL0+HhB0X6pOe32PpFIGhGh+UT9trmRFhxVY65b3Os1gu9/5CQd3
KwuZA2QgL6B+12gRiuWkugZRQQXBRBPP8qJzLktenXtsoJ90eWk3N4hvme63l/lHwWKg5NQg19pm
f4GRpfkEYBMXBcfvCKY5l+K9340ONZ3I8qth4wrJEv0kKrWEDvI2VACiSiOTRTfZl9kN30i8rsZH
cMA5YQegzwp2QcY0CbaBry5o1c2phoujOLTAodD2r0fVvBlOfzAqTQ0PYWJvGuVRGsbdgWr4Nyb5
tbgK9o9NTNv32SaPWgHqnYqhvDCij/9BWOkB4PvO9oF3C0hEc6XPzVhiuZWdyfiq+vmITjDa0dVq
iw0cKssj4SKokCYKTSGn77U7QvivhLXeT7d8bvd6shrCyY8lsqX2PVthG6ohVsIruJpyXnwCgMh/
C/ruWho3RiWjGRiwXlVwDUlnXVJMlQGxR58e46yXv2zzE85cUG9s9p1ixLF0v8RS6Ptgm+3tY5T6
Fufynd0a79rY7PnN6W4lOeLdsr+yi1nKamUn5IHFvanUhAHxCC2NdUebamt72Kr/2G8vnFoiswkr
1xDtjfoG+0l0GG2XSDxStxZKVw+g9oJBIWZWEnt8dqqQ6aQOb2wQVWG9wWXZpAQS8LwUm+gh+TPe
LDKeCPBQITIXTOF+hqh22WVL8LSgUrFt6TPPzXgszZHU9HIvXdYHqJBIz+fpzSD6FB1OQmwiu9/d
GwMRTBUfWizjYYmr1LIk+gH9Kha42aAtT7rW9ROAmxkM6AEbZTpjo4k1jRosp2xWbYTjfnX+dl/m
ZT6GmtdCivlUuz2qyk3Vwz1MT3uTzvBQb/61hWbBFssAg7sKtg/E+a6NTE7p5Ko0BLkpUfMGKni/
j+A4pF494yq9ASNodbh+FGizC5o9R2gz1FBjn0z1GAb3+Yp3Km/rLSaN3q62p/fcnq0Nv/fpmEie
URI+rHYih6yOMAr0fu/jza5b6uqvAd8Cbx/50bPSg6CBz1klRLCdD6U3DxBBnCYvEIva8TPo1RMH
fcuHF3ytMXyCCjmFaAxSpjCzkDDW9C8Tlna9Jt/V5r4WC3BcIJfsLNXCaMDuBHh+sRjbWLpYVX79
RP3sFWrhPcRlXjj+jVmcdOkOYP7CsmtBv7d7jCqU0MgZbsZTL/b9IJR67ekNsOEW0qBQWrjoKDCY
02zqichM+QmQ46kzI25ywnkmOtA7H6uoH4HWfg6D2z1JG0VzkS23DI5nFxVnlj5jqXDwXAeSUfJH
L7HHiM4sRIS15b5rHwBQZn7q56+WAHphEr8kRv9Aj8ifatjlT2J+qSbRdoMmh3vyBs6iLuy6ZIn6
cIvypNx76cb8e7PRgK17nb6e7qvt5OffFJQ+QHr8zXO9z4unqDUlG7+L7hDk1Fa19JKEUJhlZb33
A2/1TX8Afj/vhzWVowlwImmCSUnehBaRYMTGsnfqpEBdj0iImCii781ID73blmVHqS0WLd4STsjL
Uc2X+n1C62iu8JSG5tBWpDUdXYyF2KkzmPKuwaxsps+BfEDaktpRNpz9rXwIHjMwi7N13qUyH/J0
3eJKPZNamYaQSxEcVDHlaI9yMXx2XWvDQmAfweltwQZoYN1mAALOuyr2bd4SoGWS8v+nATlLERCC
yWbW3cS1Cwb2XfcbVttCUGuCHB619CLWlMNL1CsT+FYEq1dutRdGOd8rght+WzlFsD0UUPfRAAsg
2QJZiUKt7Ufc31S55mHexLABXBF/5dU9/ovicFrmfAat2IeChuNuwfSf6l8AEqSNyxYXsC0Nlawp
EYL7WDGYtJ20bJphjYC/zKOfY12MOlybPH4r2tYKwYqxpNFFAnC/4obdFA53pDTLbtMOPbzpkvNJ
TNOhAMXXGrrivQ7Cs3cuMlPZNC0wPrhwM9tZUKYSEYYKj1rk4dBKtv+LkifSpyyEQ93UmriPcg3v
/N4+GV+udy0hWiuASheres2Wvy/tyin3O7FYtkN5Z2GmMPsPb/BmRMNxFpH83kfAHW+udkLt2FFX
VOWk8dkjcp8b0bEOzpFo6Dpwp8Oc+0gz75qNTB9o32tiELxgk/NPa+8pXMR2ziQttGy+HT2nYbX3
gm+XT1mYYfuPzk4X0dlq+0m13ODRzb1BVhetI76HQrYfWAdf5cWoaJe0N6tT5TFtIqFhJMGqBOMx
mOUwTth2rz7KKgxrRIE4yxEtlTbylAFGbOQbb80cf9N8jAmd9qm31qlCYFwyxjLN3eRfe47IKaxo
qEE4/9FKCSn7bwQ3I4IMZsvk2WWrhpY3+rlxiJpqDYFB6cS+6Qlm5QNu3LJKm7UjJ42bY6hzft1i
w9crSQeTTtraZ2EFjuP+L5UjcsYVTEhit52NXOc/ev1EYwk1MRLA2whreq9PD3xV39oPOqyAmdnf
om9ir5N5ArCKL40eA2EpPLiWpDblxNTCgwZO94cFcsXfYfyzGSjCsRBFJfkhmLYslHL7DFc232FE
NRXA2uI1sWV8fRheHipTUYbhICpCdNhN1bd+NNLsJvsCYEGP2ygTZz5MbK0v2RKxrXmYEk0PI7dE
oVJgw05XMfGav53mUr2XEGu9chFBI7LiJeuY/omnf8h3Xkv2e5oVUSkX0tMSwRo1BNvrF/Tkmi6o
ogmHv5ldSO/ggrmHT6YTVx0+gXQv1IY/0U1dUQI0wuvLYJKfueH84bG4snFGtV61oJe4vm7by0Wa
16Wp/teFwBPfJVtVrfkQFKEVrPmSoSuhAKFiBfHqvuLxbYL5yoJjdvzX/PBU3zE9q4FLuCYkDk6S
U+KfoAru465yNki6AEzn9jPt7Yh/QYW88p/ahAcxX+FRm6Qm5MagzGTdm37Z+7VQ4o925LgLv4B3
pS7huPDDZqEdatO6gSweZKSmOazVPBE+J0jNB2EfFfGQhEs03/tIQKnSx/Q+6UFeqNGgey9bUrdK
scua/DEIf+jU7sciSQKeCSU21ma8uBHaWlW6J8vy99O8RuQRB2GNUBPIkPHzLrBTSFuiJPPDyOGW
fl9/iBnQf6EpPXiFb7Xn9DLXJEdl9jrKfoWyqpPB8e+3MdIFF2q2eiQhGuODWgYbWXHeyPucoz54
DBrzaDAYezQrvt+QnMiqmdqrz3+zOWdx6wpMzMzM07MBujinpeEtSTZsLM93nbM1fJXwhGjYSBLq
uivr3Jrz5bzjIEZXhQwnnafmQQ16nzsqBoOhSuoYGI51mTxGrHG9CC4VitCMpbv2fiMY6tsJrazK
1yWDPV/1aeB31WHxuVDNcVY4Hvy+fYz2zADUtryct+fhuTgPAVhxuf68JzNP/QSAubSCxIeLcSLM
GCeWsIlOr8QBIapa00d6HtOFG/B9wrXuy28psWVBK6wubuLuwbCEiv4XVNhEBq1t+d6SfYJtkfe9
RFuxDKWNdN/uS/P30QKeM87FAxbU4D4FRk+WYSNTkKO9nxCY9D5r8S7nY/efc0bcQBhLp3Lxb4az
XOYbvQcEWEwdHznk09vTOplKiTMUwuNDMjtgICE0uD+9csa4yeMh8Sc+t6tpXm2PzPWW52CRboxS
lAOyiLXERnOTDTVQu323AKEOaU2IO0WWNIH0cWWjvBv0gvoGuE6ITA+UCJ66IVAYQrEjdPq8RIZP
DWvsacJXywnRgeV84pHWQTTzTl/+63KwWVZBkjme4L8NlkS5EVqAxmI5m2Rb4d7Vw8rrvR7GApyg
wGqcu21qWN1tdKqkyMdE0bYOUn5JQa4SihKvnIplP+b0JMy2RBYmIyIL9ojAWy7TMR6ASn1xWk+j
r19kHr3pF6hb9VMns4Z2GzhMpkkcmiY2XG3VKFvyM+z6K6NObWNCfj0WtrvsP4Ui/GvKzGr3jdao
VqhQy9wOkGKBlR/Y2b5ra4r7314H9mpanshVyp375v1FhRgqR7Ynb5m5Z6t5ACDl4kNEcjpGznMO
ESjbYfJKfmwb1HLr86zKc+s38393HEebRIdBc8Chqeq88nnr3zvutO+opMGnelhwGdIxIaJrN+0U
18NdyDd0QMR0wbIquQNuHngd5OlB23qqiPLAVxG50iBd/DhyFMbU9AGHPkI1R+iABw40fkEUCMk0
IoTIC19Gs60DXgmaV9G7e9lJrL0CewhMKf0BX6CYT9TtQj+fpNGf+XdXWYn/9nBm/BlAJ4jbdE8p
CckFjY3d/i9h93RGGOAsAoLh24BYw8mlOWxlOytI5Gdh6YzXc5na2T/CZ7BUHjXSC0vv9xs6UUVn
xapPTJt7PxNq2zqFQdrgTA/+U+E2KzW6/4MiEmSRgdJQQRGmrxW82S3Ki+o1ixjRQx/l/X9JrF0U
dQJ8fBrufFciyfbf/Thvp+8HmajzlbOY+osGr4hRfA27qMwcUBT5wYfmx5lQkp0w/778ZRlFWwnM
klGPZ7wmvB168I2ANinwMMl1mnIYssrcfAwK2MI3Ve1oc1Zp/Lr4Un05UD5oix+Q8OPgaJ9vdFhX
yWA92jZC6y8IG6OgqHeutjydE+ojagFIglHlfYPy1sYGly2UYITKn4QBhPURyDA+yjw2cfW8VjkT
y1g1aWKJW4a+gsntBQusOrSsgRUWjQwF2C74O+A68kfP9nnaqICANExqbSvCfNM3LCovosjR4ctN
Br5Den5aak7/Peorv+3XXBeTD/cAFs+OmEHm+ER8gLWlGQWttwRlTMZQZ6ApBPzwbKVW5lgtswzg
govTyMYPLv35oG1Wgb1tiQwqeiSXVrEzvDstroSfmQjHeJ17/48rNnLC0zxVRvcka8XN5goioiCY
nqED65GdbPgR1AiK5FMk7zwP84pnQf6nJrRhZwnVctS9JaBGhbErLuQ9fvJe4nZX/jyBOuXWorbZ
foXUSOhh6Xf/kAiO0GbHZZPOnSc3efcyVhaA5mzRwHFzb8FGx1wkljNeeh+9E554ErI4bUaY06Gs
tBIYrUd7IAerJEvl35AuW+h1k0ZYtHZpdSQWd1/TDsJT9JhTlffZrnYJB32nwlbcLK6qp5T4D7O4
JJGIeTAQa4DG2L3YQRYfG7+xw1sMyil8WPaiYDG79WhlLEIl7VMxy0nDxoqQ7kro+vrZXGZ9G+qm
AcWphJOS5TtIgpqx68TNpdPz4cbJ01GKu37Fdb/IX5nkKIvwZ1DSoiXEVYEy/fCbRsxRTm+iUN3w
tHA14OH/lLZ9Vocw7PUOc6pdWxTPq445D8P/lYq9otL5mOCDdyZVK6lH5ndgNxarxOES5VZXI4Xy
hFo4qe4XxVfiK+0RgThvPdtTvnXOm7B0lCDsoOSIBPY4Y/Nb7RcriuBHcg0G2bO1f6yRcngWFW2x
EohmEn+bgY1ryC088FzSlH/BzoBMdvbojn/sIlZdwMRMKXMkDZmoIrNJn7X/0q9ApdMEfeReP6pu
TKmbkDSGQxtYbxLEJDQW5LacRmQaUFIiACwkayf5mpSLsl+akpi8nmc4zh457HnDynv2myxM3tku
MwvZq16odiyg61c8HgALKYAjEDbwOTE9vvoLBLC6PsJ0yk70UzZsJLwGAhVyHdJXonvyMTJ2mFjP
N5LM0BI/3m6BfOlOrXS0N2ovruGVuIyzJQzIa8sOELKibczKMZQoIl+PWZqJ/v8521VtdO70ZSHP
K45z6peYWZhV4Ox/AUZyo5G6Efcb/4nkBQjSJ+kWqW4821nQx3mlTc5yAI2JKo0Tm8xC5TF52plr
Rla24MOZHfNEKv++92xDxwH+p3g77aJqLn0lIuMrmnshl1Rfqo1LHv+YbZK5KzGsE2it9YgXiUfX
9tPTfUaIHlVCfVvtN9aHiKBZo9IlZpSU/K6/5l2SrDqW32KJh4CgRdeG/KST3VDH0GKfhSRyTG7x
9QaxjlxPq62DaFpF+bs8Dyjg8GO0008SfUT5XM8rxOb0v2rwK2umo/RP1hFQt0U5lSfZ32dR2faS
Uaw21p74NMoXUnE3T7DUj6q0Yg02syTK+RbwBltV18h+AbkbKA5D5oR2APll2vd0424zVDHif1Yh
u9t3qJhdcfEjnxG4B7UKH1fKnVCN34Z4Rn0xASA8jofiTo+yocbYeZmrpXIgLYy6nNaqHuqwKpGE
iowAvLArPfIyCmCgkgJt3cSYjNgTzdreZsZqRlj9U9UD62YKJ2ZebTusHFRduOonphEPIjoPcukO
TCaVWd7yaxr3RBae0l2Pib3TyoN+YeN0Oytgw6M2hKaodPENla2U08bDLvFXvHD9zIa5ZVvfvsbS
CRKxRE/5XOkSnLvhf93MSjL8DNc+NAnBJT8Tt92MF8FHnIYr8ArgsUOelHsO1Jd3bY7vLH/hmaLC
7+Z7V7egJmsxmWlJGWmG2oLifK8R+G6RxtuxeikImw2PgZGoDApW0E0jPlZvsffRyMr/FqEeD6D8
PHfm3ccv3p6dg44rwkVZj4NxfFoupvtC3g88ppB4dDBG2bwBacQQ0vTUCVJriWGNeyuH88XGLQZ1
kUmApeNsSpJlZQiFNs2cnDpcsddWcrV/2Pjyi0osnHUgR8WvU3toIwVeQvBVQyJ3JVE+fnvJ9125
3cAKnV5EuWVh3ecknCiO3eoClNb/eOkb5bW0znvEOu352lBqNZODmZFlWzyarOZJsGc5f9Skg9jS
0UINBnPEq/4Fj3GoNlevlf9CLjHu4oDXVoWzotyRNcwXHVgcJqvY93AFq3wnBTyu+Ivj0wDyojvr
xbg0jw/vAeuqJkfon+Z6+kYSMfUYiRUfyRQiFgM9MZma+7xY/iPErvbpUUOhpdWXLgHbPZTuqrmo
KFQ7r7sSwyGaxVGeucyaPpOoDY5qwQIvG/MwV9QjJDLZG4LXViYg0mnIg1VLHdigU62/UZs/BlV8
DHeLZutqva88Id8CynqfFhwcwIBgdT1z6bG/kOOF/MRbuq+Ax6qEDuRmkbW1CRD3e3SDRI5PXITF
uIjVWdl3+i16il5zAcY41RtMI9pXAFQI4lwkI/Huc1OpDZAc+8W3RUNjGt9gK74Dzn2QaTU6kZJt
Ppp2x7Vb++COaLk8qnuT4Avmuoe3a8Tac/DkFobQtK3Un4y+oojMLW5wQ7VFG6ByI0omWjYuqcPQ
KlEPRaxO2+tX9Kw82bmvL8w8EZZXnY3q/7SP5GeS3fWAVVuOeSCiwiF9uYgKNxbf1qaCkcc5kOG9
ntoL67dscgm1z79g3Z0gCgqn8lmoNJC1yJY+Ue+TvpD4N9GH3V2zzfKeUkZXyBiwqWt1rq0ESl/d
/E85l0Mtthdcd1/yu3UYFwenuV8Qv7w64JLLNh44uucnQWswuAGxLgWAoCVSvDibQQiW+d+ypJ94
js4/9A4+A9PTlwWT8XBZmTJpJEt8KGh9GFl+lWISxnw+/iFTvVBTFH1+6wh6oOttJEAIB1MehfrP
rQmoGjqE45DgziXJDM+gnDB2V/MTNuVLQ/d3uCj/s2nAjnhpxQs68hFxwKWZdph+LxXNz1PsyCcy
GAASESziEnUXRoiLJvmUxJ5RWQYvpNH/T2Q42Bc4Veto7hWrDUs3GqShiTk3sWv4Xg9IkpNQAe1p
UFBErEBE80+1J+A+IFkwi4D40yIanIMK6h9Y4mtUKKJsnwHr6QmFNMyQ85Lb54OaxzTmcYBRwAEv
JOee7ZrjkUf+aG5jB6e0eJKCn8MP3FUa23k+rg33w1Ewon5A7frQwVDPCO2UxPMJIduOtsvOe4vg
LbgKbyI9B+Z/iteJkM1jlAlfoDFK5/M3WpwvU8EMBURI3ZM/KrDx06h61InFaqR9tkjHGIPr3pO5
X3EBG9RavopQnsxogiJWUxFEsqRLD28jpACTbMzzSNZpkwsYDLHPuyth7QWx+bS5R7iuJ9HCxC1e
gFGeG9nzGGqdrLqYn4EvQ0oaJ/ZfOo1m3g5Sal9S7hJL66gWqfsIaU2f42FGoKxda3NAeYsBvzS0
9uDG1Ah/MV7ptGtfJo6vDdln80Tm6GmQSoe5MCFsIfNh2WU4T0M83wNwLAxa76csyi7RngHAf0cG
aX+B2aKV47L+RoFw56xzSxBOKRtFOKXdcIlNPt3T64zCZuvq5GBfqDyouXCeIvOEogSXMMaNg0fq
PSzGT1A8OhvHsupovGHIRSOeCVKe0Vy33gYF9dMf/sT1ol84UnRNNm93NSkKyLInMWJUMPixW7l5
RkDTrluDxNo478dUq/mLmtwOITr5XAGLmCLzcQQLNdRhphS1ivDz1j5X2LimmRKsdrgx9wGhFTSu
zRkTrT6GyxZzYe4SU3lEjAPYc1apL0DpI7p/srHwC0kfjfbMVhidSb98yiXSqb3xehycSipvujDX
wjzIpt4ZVzUFq9FDNcmmMWK4F7tpXqjnbv+N4Uwt7HqMN9p0Z3BIbI4RcPX7l5oW0+ArJ/uMpNek
Wex+whkIFAv4ZoR8eRL3KnZtz0UnPY/T96aZ1ferK1D6rrvM1fdTBYAKtBEpOIdhiwVr0p7iheUv
qbFmBLR5NQg5PqS0BjcVZJgx/M9XXCktWkFPNQtcqhZfGWnMw/qN6cIWUZ6KschoVi7cy/4XlgNL
19shvw2Do35NwzcOCEf8/q1yQSHqSf9SOffHmZ4ka53oRLKp8wLcvgnHNRZT4vlBYPIU8Mo7qqyO
rW0Bah+/T3RXDthyr0YA5dmwUJvQ+Io0GWJ1k7lDY260pb5Acoj0Hl1DtsZIll977Y4Hdm7sytxk
TWfpyaajUC7mYMqlKFrJbrUASqSAWSCoJfuRjgAL3x3waRzpJlDps3aI56RLIAeyPz4UxJUJYL8U
B/jnsiP5ac96SIsM50uIYLLrfj5cIUd5Bb5fLoEuuwqaCQms2I0f2ErGp4eUp+9z4lyfPOX1or5V
KVgdJdkL3GL3RTBZ7/oA2SSjNt9oXkchnGhXpWoCX6JypOI5+n6UX9EWgworQqeUMxUmMYoZZgGM
8RScJLM4aPtvRAlg9mgBQDLcIkxHDdMEWWK0spMubas8DLh9CI0F/WHZ74FRw/k/DwbxycxEXu0V
ctGf++5XfbRc55DzTfiECiVTnIAfnLDM7u8IrC4DkeVVqIZ41EpsZMosh0lOA3+pxAXbt/U7ctgT
hOg0jlIIOvfzeQXbk+Cba1pCKkmfs7SBDqgjEpEJO2LmECdB4WxRRTjEo37Ljc0313AqrMuobhK9
juKlk5EtxG2WIDURcBLlcjVrRmSSE85iHUYzHfxxA2sP+avw0HrFR9IEz53hu+6vmRlDZLyKF3TY
XM86tGrsPgMvzr6b25bat0oa+kzm7djKk5Q/bnrYx5D4tSeNZkT1HrTsYh5E5cJjjRHtm4fn7ARb
R89NXV19DrpKWRmzu1yAYoz8vQZalfRqoukakYhq6YAiesCwz2xihfLQevAUZMl06RVrZfGvTknj
lKw5UasK5yP/yP3s1Ss5Aa0910UGMSgaRpEeaZf5THtTT9KWNXfqUmPGDScH+tYTmyiLVN3M4ZZL
AmcK5Yg0JjxfRYZr2C2WfopCL1cDl6FLlSP8jQdrkKLCYFonOH2hof/Y+mxoU+FeKLBvlzxIDrZg
3K/ynGKXSFTppfQh9T6D8xy9e2sSl8WvqoaPvHnG4Vpg46VB1TF5YRr8N06HACrkAtaZfMAq6mkT
LIooYJb7GQmuwl8HXZ6ACGPiXk5AHl588yddVgEL/+ImrO5jwgIqFw/oTvOnQQhKyuWxsB8ZltUN
dviTOTcYOSx3omdPUck58LkMbf6Tzh5TAOrYESVPse76DUo+/cCUDztLTEKCAbmiJrJFSReJDezJ
36oEXcdbHwVTpP6Ztwq9EuFxIxRXTbuGYX6e2qI5fP7Vj2Vi9lcLI+cHIgeOXS8y8RGyPVTaqcaJ
QSERWXsQ3dB8rSuZI0kPMkZn9/LhVvf3US0SAjRLl+HnJTP+PuFAPuWKBmyx5rVDU4MAOxYObc7k
9eykb/qW1KtjdXbtinoRGVlUR+eABB33uNRugein4cFkjKSphI3hErapPtJWzAlM89IDMZgxbegK
CJ5FeeTjG/ULQaeiGJQnVlRk1bNO88bglA0pP+YozmsbbXmqanSQGtVs6coUNzFjjtZR/1ENlHF+
zT+kZ5eWbfHuIhA9bt2rVN20towWa1EE0RiQmSmqZcdV49uOpDcMwY53MCQtitAJRcU40OuuzF7L
K+8ud/0luFZ19gisP+RQNKvMqDGdYf62Uo04whfL7tERdmDYlTSO3WgoXmSoEIg52x1Hjf6d5gE7
mDCob1vrUkW/aEhXrWtjtAa2lX6v4TAT6iCUcOl4qgSOuXvYNCuUhCaitHLx6WU0G+ok+WSSgEWf
tmf6Bpnu3N+qX+8H+D0LMwdBhPa315X8t0GR/rD4kyFCUOPSfA5CNU+VCAkrXmEaK+XDCr0WFrit
oLhBVFfOM7CuTO0EYJUp0dSAtjecMvPEyOYXpJtmSyXCMiCU5TfVC1DoRTJKPBzSGVFT0za6A+RN
O/Qj8b5ASi6eMWMh1a1eK1bCMoWVWgvPkJ/y7NvxuOUcKcXaoVYJiXra6IUuJGaYSaMbkcJbYKK8
qwle0YwlbT6vJ/omruQY9DW4+8y4S/qSlMzyINxLHEzV7JpxvBBArokX39Q93C27Dzs9056n3GTv
uX/0BQRjxmcWBl6/LdgnxAZLoWRevA7Xwqd9895btC0eTB96sUrJJrErRWoW8c9w+5uuu+/gqgkV
wn4OebZnoHCGyfOVTiNIRF3IiwcGSMD9RG6OjnUWT3srVDtWNqQjj+8H4S3Sc3NYYWPJGy11ej1A
pKLs5TH+aG6FcgqqglcZft5/YhYGDlNvdLiQiwbNaQWCOR0eA+pgIpwwesTFO4IU8JviCBK3I3Gl
wwcdbf9wkCYRQnaSzRvPR6SXjSLRM0L4QTRfYSB/JBvzczs88/crON2ZbumYRhjPqHcdqqXkHb5l
uWrSOAxhhp7emHXsIcFtsSW+sCH7mZI7TNeYVuD3K9dfikxNqZ/nhwN3vVm6VLoQLXI/S87ujuVX
4Xpoic1uG+hK6EQLFicpZwaDEDkx3jCZ5lwduU+UrOs3EsIrN4mD/KyYcFe7IohG0aEhIEAd6Hyc
/5NmP/9DifAsiBax3s9j0tRTQN5uwfb4sI3Oo8+XrmdcDr55x40hmzwgOOnaCZBRfPrQp+lXAGmW
Jr+0GBG3BxzQ3YiEtnKwZKzjaBDJ+GNyyXwKlvwRg6erj2bKhQ3W2PavyoInS8Bz28yzdEu8SU13
GHwN79qQfyXFZptsZ0UsbBxQqiaD1MY446gEb97kR0ZLBf4XFkuy3o/8UsXKvYzZPpdFmOopTEea
No6ObHOqtdwbW5V4ZGsbz0Hs0DjJDtmHNliUNVyPfKNPJsuDQcFzBcBLg2efRkGod7C57sNqKXvR
T6UUN05oIz06GDKvTeV9jVTUniLeU7JvR/kCJQiD4hl6wEA1uFbIpmaL4nN0TOBqfk9c17TP/iEx
wR/6WllKYRsf9+E0CI7YKbFSmtK+FkhY4jPfVr3Ru+DOOBZv7g6/NyWa0bx2byLb/X1DvZiixNvT
Qps1UcRypS2ltSMDRjth6pD4rfONfzX4Wsq6smHzi/p732xqtE9bs4BsfEcZX1MKqZqtOIlc+WiF
n0ZVLRHs0TAXB/CA6ojtlFx1tomOV8xdSRntdpayMt40Wo2Fd3soacsiGOEJ9eBGpeA1HN3Sv9AP
b1O83WF2ZHIKPdVP8RLk+6qM9JKVvRfnQWO9qxjgxa/qcgQIdqt1uNHaU2kJ72cwsmXeMfQ3xeAC
YMmg+jv/ovkXUGTNChGhiJQXzB4/6EvSsFnCgQuIdq+kuXGUt/Ogk+Xma+j+O/F4eQakpcs6ODOQ
TAYCGhqo0qBHl9Lh/ld1X5Ztgi9U7LrKHbyJTfmGiQPmuoEzsAX9K9aOHUhpzEvYQlcu89xUK4qq
v0muDOY95DgK0UBtMaz0xeBveR29fzm3RUyz8tiK6qVuNyWMJxZHk/oRgFexEu/sv5n0XJKOfeH3
elyUi/+7MstOa9tCBSqunnOZ87WWiGuwhRzIvj1LJirXHoce/xQyIRYFyoYTs3Ud0/EDHpMJj92d
YsHqb90ynqZcav7Tb89az5qMI3W+xkOVLWteRf5GirnAPk5+io6LWUEuGGjSbZJ3lDBcBUldm6Pe
SGTdpKZd5n/E1VEFBPPsIMGoeaBTM+gvx22caZY32f+QArux5gweoLJaSA67EhtGvl0Dvws/SSVv
OSvQXrZ9sdC7yNWbRDHI/4qMs93hyBScpnSEREx2XUTp1hFBR84hKnWktOFXxK84zdw0CAwa4xbC
wbVso9I8/h0ewts4XXqhewvvzwR4sSjQgcNvXSHjjiqu0LokqZBtCcyt/K6ojaHjeKe/ZnHkTA2D
/CM/GyrX1ZLH83axkJVdIgq7hiSN4JvUIkdYgvuz2v9iaVzdI+NzKWcrW5DwYiiZqbLU/o0OaxDQ
bIWWRlTIEyLtZqJlEI02X/w8+zMg6g8f8skSRES/DEiDTNm/DQetBlCDQdqFrg98bhFoofFJ4Mej
8pcgHW0JO865djeGQ6UVs5dlU8bQcCEDM8Xq8RcQRNyHZ+CGMh0837OrF+O8n0s1PAkcv2gJ/7J1
MGmy1UboCIqCrjHUBTZi75GYFP2ggZpKXPAuNgW8Z1W4fz18F8p4WzJrwSP4LqO6fXw+1Gz615np
GacPrV9iPdM3WTrThCVuYi/flehEcB86WokrrF235cyTAn1CYj/qx78OGjISiNlEEifFjdB+HeMA
OmKbWP/KJE9xzhsEdQQ/aMMweGlMtp4CQ+dtxsRle7J4qg4+j8DtzTrgTxdjnHWm2Jay1B4NNlr4
I8w0vZIb+l5752yDIsYTh4bKXxdM5XdDRvX7ZIjzDJqZlH3rggnUXfloQZRypwmMmzFsddS8mqas
+j1C6rfBy7pMcHTR8zNzvAZM8Jitazr15V5hsqXY/cueJ6Fgqi84eiZ7sBBsz6sP7rq654KcnbNZ
94yTkDXAPBIhmrW7MAh0zoFPSWtZdGfgdgWNqw3qR48NeJ3RXGiPZYcxASddWRx+ZWlpO3nE/GWW
oeFT0pgEVJz6ilDUf+5kBjc0pWJw8+ZEKYn5rAySNo1Dv6loHJucAeePNjy669L0ojjqMoNk0axH
QuEExC3xA6ks7PCjvgHJ8E3PbpRCNLT7UoYd3ya41Hyh59OC4i72pbRqpi3cK1T+0XTyUW48Sarw
UoH7X0rIUfXZatyI/x2BVEtJ9sXoB9hFXuLlTELj3nYou+bP6h0D9qQyav6qa730WSGba6qQcsuc
5INfrO9ZYt5P6I0FQpZd0YFKQgwR8kF1Y3q2Z0+ksB3jhjP8mkv+kvn1rm4UPY26Q3Ot9NW8UJ6M
kYjcxx6bZNnIk+XojP84lM3xARDDr/pK4EJshnB2SFq7Gr5vO3isZkHblJMFGHf1Clzc6YAfJfwz
Z/xxpavKcPeEhxKp2E+Z7fErGT0tTX6ixok41gV6IvcbCghm9zwhnp5oRtT2c4wSIO48FC/ygkmG
Kp6WqqxXAu8/FYgvZxkEkY1hmtuXfzBKfVo/n2QuAC19z1GauKLga6yNt9GqqiVOL3rLEY38y8qV
2XLP2PWJvEKTz4gMe99w3sjBYJqXBoOPHJm8CWw567zDG1EipyCntSOWlmqf1Xe13aNVxMcrCGG2
rrJYsmmqWBqqAPwKtpr4VbyEObFxd9CDU7Q8aKdZXM5v811X40JieoVWZuMJPPPATLH/q1DcHxsQ
BkXhQOw+y96v8vPu7dPWx4WmxRfx0j9PIynQrS0c93U3SOCj5Ly5cv8PDwYQnWrw4dAvSlVn38NV
yRMs3WH23zkU7Rw8Vt3N+yGelPUGmhNnSrBI7ZyvZp5YJXzWfIQmy88uXNapbbOprHjoYZN7bIiC
fw9uUYmTZQozVgdhlnQkPNaVojl9Rc1lqSw+k/SH1ndeKttHYEcZhGXS3N+4Km240L5oknSIUKql
b/sgyK4ch0TDjrEb5VPTrekrbBMzN7F3V5Ip4RnuzwFQI+TuDQWeFjOGIuTSBLSJa1qIQCAJqxml
t+rgQ5DS/EAipHtvXnpv9adgakVFVdwYC8tTo5/ARYBY5YHU9wAyMNAnG7EZXSdLzCauTQwhY85f
8X6AyQW0W+H0hOWI1j+B6+aDxCS1Ti8Mxljt/c537uGoBJzkmtSpcZSEmMVJR5n4VGv+fzJJ44nz
wrRGaMxAz5oIR4YSLmltCA8mTJjfTFMkAC91gbbvmdYIUwzcV/QhpYUNlUSjoqUFayw2KV8As4ut
OGVvtMtbjPWf7dmsFxNJMetiALzg/C7acHRxo2NnDOGAIyoGMQqsHAuPOZyDnF11A9HBC4NDNkFc
A0xuHAJk3J2YqGy+2bOHoEdzTQVNiaSLKxUP3RbcT18XwWqf9KqV5ZNMgFpFRA3tcR0htGq4hGoM
4xL8OCMaD7JKLRIIyH5QdR3dILtTl5WyRZKachMnnPwv2geSmbhSqeBixQ9DzzFy4B635ta6RF/t
yy0Sizvk/JEht2dZPKLRqKHR4oy/gQwvtkMR83E76isMZYgLBCXt0qg8U2VmeMXsN6ptZ+eKGdxL
ROpxzFE0Jbs9QyQlnRJDdpikv0CFJANvl2e3mfBgfel2oxCgXSh5FV0pDqQDINn5Qx2xRWR3dtpd
GfuPTX0iLEGTQwGYF6kvgAtTXrJxW0TOGWEQ2UUPkc95kgsiao4N9CtD9mfxjW0DMgyfzudoD3xB
ufq7G0Rhm/CoUn09PjBkDevhRxFdhxPQGQ7hh+FjJgTuEOYXFHmFrmFya90WugqiVUmb+EjXu8Qg
MOtODctktgkOz5DIpAjh05TWEXG+NUED6tVg946NFWVRGRfNXrwx8dvDixnUhQaQjO0oqQFmPLJS
Gv7OuQA5Naze8vSTKZNZoyTDz9U1CgqZI9AD3tYhaEDJtAYGrdY2VwY/1fBAmvjvaQ9NFfAoXw4r
Z8KRdIJaMaFQy2hYUkjj9T1r1DAN7tDEh2SXhtcAF00bCCKk55mE5we5aiPyw22VFcp+MXMAvZfJ
dB8CMfSFfuB3gv1Z1+h8lW24sdpkjgses00IM/YTo204fdqA4molcgRQY+4Ap88pEdWHXVQ+Kzev
YnR11PacZbGsFlDDOV36IIzJf/CafCcqa0pdc0Vq0qRwNAl0QK6FrGqU5d1f4qqF+RpalcpVtRU9
gTqoJ97FYx9chlHlZLB1y/IhjyJ7qCUFnsTTR6BeUL8y8MIuZ8xKuJCBhes4WWHpnOO8eIpxn0dG
3UsGIxHgcHDn7hhuZYlqT9KF48zz0MQ8DJP3ijYXX4Ts8L8mvyqJiWqtmhVPoQ2et3tSMNZXmbYH
klleb3pE+VMlStlPw6EfhTvZyRRx7MyBkSbjMEmnfpge9rWL6aPKR3hCNdjRC5u0IhfiuVOJ5kn2
pIqFa4oH02L95ALy5ZEZbyzvs+q0inPzJ2UQTk3uuo7k2uLwovi0IIZ1cEugVljVHB93sjgGZBE1
cgJ9AWyQOOeUCzpS47/LdWEtvZQgmD+blJHNfknSaAqb2Ced7a1SdqvzABAZ7UZlFHAGVVlGNB7E
IYhDiwdOiYpYe9yJ0BAOMyLnJAXjlvdGk/wTpOTfZTcyvbbFQyfk2R9iJR4I4j7BUp3fG6X0FRAS
DsHXrK19unE/BA2NVszv83Ol/6UxsXDGjFmSt6SxV4dKkUZmBaAVUdoJNkaxw6NnU+w2bk51k1GT
QkZw0VvD694TgjfG6n1rRrLJxFVPbF0P/M05/rfyMhWWda/bB28otqnWuO4BvrYYMGlIBqPrJsdz
8+bn24YWv/QVH09vtXYm/vMJf+FRSjjTDobGyqd106jA8XJNE77ttE/6X4R8+vXJTNGpEOhuO3am
lM5R3uVLsnSslss8nJa0zw/g/RfLHBiJH/PoFTOnOP/DjCooU70ca8OOKw0k2JwFAPViKkJK0rSf
5HTkzG0XHTCf1Vzckz8zCIKFdbEk+Z2nOqsD1X/0co+tUZIvBprKdojaFjrW1X6Szs+zQdJF65FW
UnY7lQqOQPqd8INOdDIG6Q/r9NkorZ3Z6ycMRFnXEHgK0svYtjpwE6V14c2/yC5xGBnw2FAHssC0
KwWq+3WuYMd6/9xHu8TEJq6A9npD/Msv8ApCi8d+KNiZwnO+kdBxDFtJzFTIzqLZONiVdoZtalU4
aS2IPQzS+yyg0Oyn/1fXx45TUaVvBcKa9FJOitD8G/9DLHO9dX1888Bsx8G3ZRMyVT1RJrGOJ6GL
tuYMZYAGCU71QYR/2psVdp4FxdIET5hvE8/kLt0Sj2Hk1F0M8xKSv5OXBsmU31aeh1z7EiOU4cfF
yhXWd4RRD8AzK5x8JO9j/uTw9QirXGcA5+vZUDAWilSMbL4btv/rq8Urhd0jUNMfNIer4S30Rghs
GQe/ra3IB7dK8GB+MY/NYpzMS77VJR3iIgbCTD3RNfwbGCCrwZzF64WDto9q6ZQtmyAkeKX3dKmd
qPJOJJgT9rdfch3IFXKFxZfE3DnigA9iUMgphu17VxzoTW3aqXXeoEIEMLePNcd/BtlNXH6oirdf
7/NscolKTKGr2aXLZzE3SI3k5g6I5e54Y800z8s9ungYBRtAzp7H7E2kteW3lQlSjbkTuSLFpNIa
k4j6iCdliH3GlEPphR2KgB/t7eTexsD89d04B92NgvrlsESPVA2j2gbXL9h8ubkHWaaeYA3De/3Q
PBq4kI0I6pEzbPEW8t0NIvmqBc44XYiMs5rlTWXwPkvJqX5QN/wiu/CihgaOCVPx41NXSYp8N9Rg
TM3YaBoesNXkQGv0ZCfaqHNqtRgVeG7oJdR+VjEIYIi6WBGgmZo0KUjPI6vMoagEia64cfrumKkm
E9xKrOTGa9wOEsONPHX0CDQuGktTwazzRg1VWyYxCPzOqBuRffhncfH4RcHBXu5T3B1NgY4Q/Zwm
gMIpicLw0uJ7r0Mru1yoE9IvkTY6Qn2hSdV3doIpRzuOAu7xQGQY6qTMmc192Uu/UeZtLowqZtrk
5/zT0QwpdbLFG8vTV+j0CQDNpTIdHDc4C7/XmOFZUrgU1hAmMws2MDMxq4PlZfJiXseLGW6bfdqP
iNQkM+ZuPTyokmJchaZXF+3ZMUi/S4YX7IfNf6eEHbylquMVmRe4dJvMaBRmqBjlxMzAxZGnXIbh
dbkPoBiZX8F4lt/gs3R4+drco9Z9Rkorzu+gURkz16Fbr31b2XagzyjZHzL8Y9eDr2gcjKIroleJ
rbn41IL7skoannrbjOmiIDBrilxM+lzcvjM+D+KNDxvHMvYIyfEbYV6Rk7Rh1Vav/x7lN2houqRg
W3490dIqzJ1H+gLTSeyYUOVFjzaat8vGmf+n6WjcteFVnZw6ZGrdbjHYmXtmOjg3+LNwoKWDKu7h
CFeiDVaksvPaUcTA/fcwVqbVfn6W0biE1/I5uKcFIJYUSlp+73+WjjsfjOmYA7sgcCezT9r6CM0s
GuzdH2pX95f6TenRntznvaB4aWSRA/sa1XWKVwIiUj88U7NTZhbd/MGeWFrLbIWWAB4FOGL601Xi
Ri4SRE5+9fhTv0ErsE74auI0wkMbCrbbbx/TSZqCeG0n+tiK1ogDipmaiwlZoJF3BPoSBEgQIdSd
0kh++VvuGmd+dkEhNoGA+XZrzuBdIQUKpdMt/pEqiI3Beqx9TiB3PVu+lEqr6uikJ6Iht5TZ0UNQ
71X8CsSlxuJJ4pL1+LIGtf603o7XlDhXZeAHKX6rcQ/mc3RgSJ9t1uSaDvQ6UgyYE+kQziAhWoBj
R0YiH6/E/Y9og3LvO+500BWcQDuBLPIQ+ev5ySR7hpAa04U7XLq7jaaO5BRrqrconI0Q3ee2OzXU
OlstG09gNxJAWrghizLNfqbiezg543P7XzoY3HEBWU6x8YypZyZm4SFv+31g4DLhYpgJb1G/uHUd
BzOrJ14qfIA19O4M1dBCssPayeAk+oiTbjFdmxvqS77PbHOmRc4Eug435OgJ3Y9Ih6qsozbidhCu
ktS480eecuckPDCG5cXRzccE0LMAKKnQbsASqiR8KWF7xV8i63+tnnYSahyawt9NGL7EvGM7JXe6
3OVPM2ZOXDWBFdJdfy6cKu6SIqcbS/aKMpc43zDu0bUStrVa/6EukKsCpa8Vls7tWjIiIDkZK98T
4CN4SRK1FMgChPoKkL/gjo43bM6UwOvQAGAGCOmdeXrb3ylRgPKNsEZA1eO+qcOMvsuJyOm0T+cu
RhUKscPEkHCAamJ+pyZJAFCvELqNFOREdsELSu0ZNtz0EinS58VA8RoZwAjpNDFNgUdHF+VGyTLp
jEIdECO+28Ej02/V8mOC6nIhd1h0LD85YU3hGUujHX+M6FwLKgcwWcg+1FIoIWYGfEM15839R59g
Gn2Q2gIypM4gLNv98NN5Y4vQtQpU/3BNsDPif7E0j5Yk73HBBtl7+aawEgv2tLuLw0ifR6mrkUlG
GRxo+zYx8a9dS7eCG0+t+doWQ5ECm5U/tjtUzext1o5FPT4wSFaVwOfoPvX0Mi5V5GZy7LupmE8O
z1ScWtkJ0H3QxfPXNA05s0wupZxExrv+NjU9wc9jxkTUAU0kamkZo/PWWWGCbmhwuoQAfGRnaYDv
x5iXQQ5SDVQZtexij2kAfvFU/HP99wBlJZMYXUqSKJ/8QjgoqwGa25aOzfY68wlfqjGL+XgJ0JuF
40zs9l1buUnvDoZwr1zZ/QdBinRlod15gG6JkrowaFPM2sE8S6zPrZXoarR4YFhsr5lT4luyqGmu
QAeXw74GXzRPdSfg9Vr0EleYazdr30F/jb3lwuyw68rERzLJKLRkSGKbM5UHNYhxw8weOepUUPgB
46kuKkRBMr+8dxiByfrZMWmH4HLoO/PqFzrE33JG1XAf+dMxMSWn7Gb2R4J8+kAbjSVmt0Zq3F0f
qy+VzPTvZWAkHx7nD6KSuvtAvq6SJMn3rS0I4shZ0WQvshy0BWupcGqFb6qieiGwGEUhTW3YzpJg
gUYMlu5gewb3kSmvh2jWAD0O88ErniLVsWU9DTDJpsn0stNQ2lo6dr/2EPo2kWCVpjANgEmGZBUA
78fmp8QMYLayHv3YkoaOoKceTxySgvqxzE1Su1CqUXuvMW0UQ9ojadtPNwsZvjAdpJkRdKwAGJGp
uydFfkzYutfW8ZzE0y2/bnQKvK4A+Ew1byFvl5xVgx3RdbiRyuoBLQbSgmehhdVSaYPf/TAdWiP2
uozg8fDUHHmeQ/S9MmCGRAE/AKlQxHJcmD6IAgQLGOBC/ZfB5rhL2K7VOJA6aejsGWs3mOpXl1Sg
LjcLABl2RG9T8a7L1enDidGIGXy+ogKLzxNMw4yv1L/MRSDOqjzplC4NTdbEm5b9kDF3wOU1dMIG
qepufuxFzPankRP9Jj+HizP3MveeD2uTr6orz88Kcsx7cowYoRcp/P0DMzhC00e1qWqXd/IQh4XX
XcdBdCBhccxOT+hjHKl8XX6rf+wiXyyFdKrevr5P4UNETgtKOhUikkcbkga+tpvtBRermTVm4qM6
KXs5uGoC0zSPyGMniP7/1W7SFnb7gA0BerEWVbiWJtrEIMGZSLjcOeiuFVOThxY8Cb4zPer4DVNT
ISnei4I0IulO04EPji0KOPZ8W0oev9hiD4cyJwzPgkDALvCK8u8SGlJb1QA42K6ok58k3KXStT8Z
sIGDElz8ABILia2922bL2HgNNtZh5uGKz1EsueFM8TsxGMAu5RNJRlm/pFh/pwYPIakE9z7UU1ZJ
VkBlvvdlAAzJbvetWuelXhWiOHSszSgEPVj1D/KKvchocFgJjnCENqMn/zSHlHWivT/chDG9K5U+
pudhdPQtM7MS/SJBhQ9JSrGQWUbtt17pCcFH3LiGIdQr4G46th4BSobYjJhP1N7V+O66Ge1ngocV
88FPyGn6ZqFWmQ4EQQcMvmKdMlpY8PVYwWzQz1Mn8Sj6nZvqlMnzRBUNf6fUH7kiRyMDar5VdhFV
iqvV7N5t95eZ5jKZ2bGJmYx6rU2LTyNklCz9N12P08CXUNOZFfrhkuBnC+1bQOb7bjOVWhUuQF77
BFFmvdkQ+2HEjrZ0CZ2Pjfp/hcwThVol1Br4wUbOVP7wy6TK5bZPeRAnAOP72cNofbhqC895KvAT
O4DpkBjE5YYq5cvv5ufd+guCTD3uU4pwLMqC5kFFUe+jWHWi0ha4RxC4hPmqjzsweslhmQvG4fhw
tIHr5fizOUPQSfTdXlPj7+N+k5pJ8WD/D5GH+7UGPJ9JVvjGOfsAiXmqB16Wgx3A6v5rzKyl9DEc
Zs/M8OR1WoJwSlu098ir5TcO5b4OZ4cXz4cFFCFcX4UPgctzGbNl4209m8TXUhboMv8Dm1QfByMG
OCsg1jI++vzfdjnoGYVDD5ZRVMP9P64ujhNq961dDyuJAkx5iIOC+qBt6RfdyRwK3CPdGd9eqJ/U
UQ/trjfkyVAq4ACeLPkgxNN4wuZtm1H25ld980bbbslEjodbAdjHzsWj4rga7GVEQDeF4Gzkdo+J
DI05A6uAjuydg+/qKp+nnTKMriWd8XqkG2RZwux2Yy/W14bgnwK7Wr7nyN9nyCD7xqhMrx9HDynz
UXG2RAFf+RjALJd+RFVAU5gwLiFqvmUnb6nrYN+JvhYTqotYnqbSAxyfArHjHlAGQqMmgPvwIpBr
LqZO6nHnlmQDKAm72m9PLxNMXM12F/5Te7gGPWRthtcgH5TLsGFJjQtY0bwC6SjI2cA5Hk4EFEia
pImb8K9Ir2XIauYhDb45+Vc889l5MR81IltvGTZokc7BX+jLi4mqltupUnECeZKByPlnWA0Py2IB
S+NqDux58lcYm28zynk5266ZzHZwVruFafdN0DUFa/B/6pZPZAncu8NlAVEnH6HyblevQtjIL2gR
+GpHkqiCuny35sac4NVqWOttlpgWLPAwxRrPcZ+dad7lGY3a0YjeZaPhvVKFm0zCXe7TzGDOYmaL
V16PBiODx0+kVFw3+GyAr7eT26NB/DKe2oAlmSOSi379W4TkdSrsXdSoPgYE8SUHxD/4PKFUYzVX
VxgI1z+kOl7KuLoq0jdVhNmRrgdbtZW4ZIg245899+8GWbld1DHYC2DY4qQnmuFbqsj0JzT5hKDm
AKShgItumMzdnoj4qTOowQVJEIyHGbMqdsp6Tsp+0+NvkXnELYgH/ZAV+jDvUih97aAos92bHw7Y
yyqbWfDUlwSp6vtQ7E0rlPzxsMNxY8G3gcvclXUZIbtlMhEmxDagf3L+/JTPjjduK/RxhrfFkvsP
bjyLzUfPs88IiGeeOOr62ByWQp+lGe605Am0OCaBk0GExVuHg9E7ieBBSytbTrpOD+95MdXpliHX
GQak3mOvPWtwVxmo1ITMT6hYMvBfRXWSkJvvU+Kcp0TmDnKF7/g+qDqSNZp5rAeSJ3Bfsyv8CC35
fSO+9wDHF+mL6cQNwUNK2Dy8iO1AM7dElxNzOm+CqY9Dm8p8xskjUfXaXH2JCRToVH+eZR/lzY5u
DRpW7Gp9/ZqermAJooM+V/PtR+6HEHZc/FELmu2cJNq0xoKUJTq2M7s4v5V/8sGjd7Y8QqTypBAD
omLoLrELdgMB4cRq/i76w1AUgMGK2fZS3DLK3oTgwbBaBoNqvplsiW+0Ow0CHuhpJcpt77vTQY9J
UjGe9uhXirO0u08ZXYQmnSPfyPssY9ARK9FkPFsNGRSeXJ/AmjKHEC/qXgWCP5Qvlim4gtMA0O98
wg0W7qY5O/GGKW9dxA89b8s/3dxfdnCMV5N+aTfyO6BpH3dR9ZZIYbele0wlAuXlWFAFskUi8ouW
CALxKsgzRkdPZlMwG+9Ni0bSdqNO3fD1f7oewUpeVGcLTa2N8VFamzkD410Vwm0vyaOkQnmbfY81
VwblO7GeetObQncBLTWZww8xk/YHFaSgPjboYYyZZUPbBoIhpRGKcvSmNN6DWu463+ZSdV5CF/2o
PpetMsSlsqSgD/UZwkjuEck+CALgT6cciIJ8diZt3u8MDvOC7gOpFD7Z+mMDMlzQkRqBy2QmzNdA
Lnne5YjSc/gDJv8W32IFDZLyyVwdy0nne68WhYAxtb6L82wQj8v0Kficf7Eq4zRvSlfXb0LSAxd8
eKdavA6WSm9xEat9QoowPLp/lLTDYUzo7zhu7dtWjitHDUmWWm3G48OAK70+H0k3KTLgrhJahptg
unQ+oReEKqI0gr2XlsIQPDT83rzfNFJFczP0FBZO4Ar384beZgL/hkEowD9X9jiUMOPLzMFtL/Mb
JU+09w7hOaS+Zo7ujiF/kWLWlPzp0uLqVpbePS9oksPDeZEvZSpCyXVULlvaDzhNR4I4kkMj24Ni
fTRD3hUp81Pqe0Jj9cmTDTirDKW65LSKsJ51m2okE2TBA7lsBNnzPBBGL3sPIeSAPEt96scAYYHX
+S51Fz+cTANZfhIeNx43Y9bwUEDTCtmvW++C1FNm0R5yW01vWliUcK/Z2JmEoUz3xKbTPzMIaP28
Gl7ZD2bFvnVs3dGFwuTRNtbpqD+U+/xxndalq/2aOeJumU25yNI5HLyoCWOvFSEwza5d/eig4wIp
2VFWfRNeNKV6M+apOQ6XxpLiz6Rnd9Gs69wCTT6+nwoTWwkDtKV3GY5Cpd8WnIM8FuvXthwAKow7
QJ8lNrxUy5uHLGlUpLx02UXfg7TPb0JipEUPO3V6GVMuF1LfLp5EOBt9NrbFckaynY1IrIBGjWca
FqClfhHsGWXt2e78shToI/f2atxOGk+4KsfHfjYu5M/U/g8bGvWdACuNqH9GfTn0p3TuerdGM1J+
laIRY5sCES2wFa0anfjQ4UN9CAfV6rGHS2SvPvoUK3pl1LLo0VvurgPeVjFYZ18Ey6SS8pbY951C
Nq2zIDOiihGJr1krSYkd8U6GdL6IWgAFvVV0rsOjxILiQ3N/nl9a8QWxbXfbeJ3rHbLK2WVk6quI
ZMdkZ/D+Ta9/nbmZRrVsO1djP/ICRI3mR9WLxWG4aMdIBF9gw+SGZSlzEkb/ZmLMWAsfhcteUJUq
D9ZpVvrXKgflDjTTznjGdTUhjHgUMi251KkcnWS++q8RsGUOb7s+ul8jWOdr6/MzpAocphKhUELF
1eEZD6aR0WXFdAScBBAGJxNWrfV7JtMxyRUwIDpnAJ/Qt0/RML4e/KyOkTpnj86cYID6+mxC+FAi
CPOL/pIrUE5BmbLjtItjjneteaXaCa7ckGCmyhsiiiyXWetEigfTgWXIoeFoGV+Kef2UGjK0ZuF7
Jo0FL5WnH+OmbgtWKfcyhiC+XLwH3lJT372d7U2tcfDNJgIPLVqlIYPQ3SQAf69tnbfX5mXP1faR
31u1j+2QVWq2/2jh55UWGSuANX2h+c6701ljeO3xriEu3PeDKMgc8sw61EB5FF1K1Ih0pCBa2cJR
7BbFM/xvv7ZftQp2oN4I+GE++A8xddk39UvgUDui5yiauOlHvPYmrIfsRtgia3PP1/U8cugJ6NR4
6a5jgSykHiAjXWtHhelxXK5Qj3+SDJX4mFLoHdWZ8KD9ExsNcCr0/IbGXE2H7kQmOKuqvdMT4GdB
MBVjXY6LUMONszWo5BGEg96oJ5NLN0J/UDmC4JTZKSv8Mj9XfhZYVWQhFY+BcfQYHKoMNVeyJ7Zr
VEWzIsHaKa8MkiVEkTzxh6BlmeWGubrvnbLqMjSS8U4Q8TdW5zNo8CaLnBqUNU+FesDgMeQm76Ig
z1/uoV2O2Z1hp3FjuFvNli1013/TJ0QcIAvGyZpQNAdbrd4U0JGksBBK4wl1ZYd0dyuoIc4HfmQ5
MH/JNGaQtbz5qb8nL9lU/sIjiI1msJK201SPX7WQHSTsa8kU3kEO+Pj4WJqHxlVGz6D4uqaZOz4j
sEEQc4jOJhkGRzT6l6Zb3w341nHDouFTQHk6CAfNoL88uIO4JEzOXIl+rjqyjL9SjCFsGkkMqYwK
SPjxERDT/unejUkknasOWsarMeKbzq2g4Wcs8jW6c+Vwlkk7qGwVYfVSdYLNTFFQCqZJj+rkGqtN
w9pVZGvBPa72LmHIqGLr0qIVzWk//UndAp3V5OMG/kwo3u2jjtKHKHcEUtZXgMLX2fuoMVmSsEWt
FROXH7bOqfCndhGweOYJeXciF0DfcYVRU4uzfTkeuLN4dzYh5Hyp/0aHVom+xZ2GeWJKyNbWRAwa
uZu+upj+B41V2+/0/GOpyax4FjwGoxFxS0AFbLYbjPkxRTEya4PSGowebsr5FK5q8XLx/aUF1aeS
qMdBJfp6Ig8QA/SisBZpBT2ctGV4eJYjMe0oPUNfDr2u0Yb+NT12zc4ynUs7xVU8SlhpB1p0CJ7d
sRX3RN9XQoyYJCt+YnojvkLl3qsQE+aBFjUyiAvb9Ztklr9yzZJlps1SPiQHp6SCP+xKIhHidxGv
UfF3fC93oBZXxBrvbvvjkAvc1wnW0eRusNYJeFJhOTljvsQ8eSDEK1LVhUdJH7ffae0TFc8x5Wkr
5zKeH+irfs+aSznKTUDCCfRudR481jsiSvDqIJE+UZBVrEjHEaiFC8YN70wuV+wRO+ynhmNR91b7
a30SqxvNj37seA5ofaCI+eYTrZb7kZVIH93v9jVBx65bwgWOz2bAr/jCAJ5Ct1t3pvl6+JUyrtiS
YmRRrTk9p1jiJpfVDgPpQJwnuac5aQVjpsLPZi31F/ugpLy2dQPqrZa/ea+xKZ2iwqEhDDjuiLNU
msvM1l4NLI93ZP7rD506wLNSUhDF1/JzwlV/Crq3Hf0ah0nwA8yB3Nf7L7idolMyiDh3ywsw9us1
PrThkJH+IRUIE3HBHJVjjLUIrRaT7+lmqj2VBiM/7QgLcr6jpn5G85sMewZJ+Gf+hriEKCqq8AF8
u7EbqiImDRvaY5YWi7M8liCYh6wUiH+PW3A840pZdgojOyCV41EPWnBUD9OMyAL1Jqx9eV8rBpaw
xNuMeFd1Wz0qBogeYSsztS/H++6tjxkjTerhDp7mdsonvPSV5fQTSt92yKEQIN1OGWnZqKfxs/A8
qZDKbowTtKbV5l0AzpjRFK5es9nAD+bdIEgjPfU7qnnE0AgjvnpSES6gwXztXW7HNuiu57jtZijJ
ANnrawrI7tjtGXyR+SiPH8mJAbcwcVFdWh4MG9nxavyjfdIz+SQ540mQ+TYpPpq/thCZHMB+35ov
dQjUO18vAMtdMeda3fVj5F+uJvA+cSNpm+fuo2RqlfORDwPboUvmoIlBnycdxS46L6AU+rW3ZPK8
IuE6KUKunfQgpni/Mt2jl7JD5oOTxwl2B6LFn5S34bx03aXRXqVv4xTyxTfozkNvP5Wh5zJpVzD4
/lSzJllvpWe1Sh366XBOJxW6xWWnZubSfpbbRFzIiDuGmt1vmD5BLJFundNRU7Bej+I+GFGgHWrz
KamsZ9sg31r4XHI2YsvHURFy8sC5PilQf8DGCxzBGDftUGRr00jMQfrBsAiZteVyKVfwc7mweca3
w2QaHzaObYqxKpu1od2tGxWbpG9FR7S/TZkNxK6zzkH5cTqF4qQZPsoGdDMS6meAutuSL4bx6/Lj
/Pzep1PQaFvJMY66BGBRuyaDsmA8VAcAdVrYEwkiUV7F3R6g+X0xcE2/Zje69+TgrXgO1bR1BevN
ir19rnawUEPIrJJBzsxR70XIJVvKNwhPk/gnIP4U/UxOWVEKiKrdJTmaHE7aA9PQjkgqqzFr0EsN
0dPqatiQr41AU8M6stSRB6/mFLFw2qXg418cwuzIPnJqJIQSFDyvdrpTFc1WsncjT2ZHFAOz+d+8
rJlYh5f21wJUOhq2FubAfQIIWORNIwgO48cZXiWrvXGmTroXXDxucQppbOgQlSWUycSBkgQMS2SH
9kwOs4xrsrIhwIb9TQR0AeFTNAswrEgGugtSm6Mwf2EpjgsIKcm6R3tmTvjb19LZRWM9q7UZ3Vtd
g0UUfPZKAikHfGIDp95cu9KLV/cIPbAyVccYMx4PMepYqmXWJRIZp9rXkM643Z4iqo/MOiOBqA0i
RXtDLqFrA4UBpXfqFoo2gjaGr3FH5SsxSVo62oYo+0PVkCyiTPBOEyqGSIEwbeft/f1mPvjVz/rk
Z2xkJTFT8PnaJMdKE5e4UscAtsq67KgYrtoSlsoDDH7ucMM1f0abwELfNGrELwhXheugzGr7M76q
/NKIVTwSeY30Bs6PbEQQJsNcGWakkmmFXuGNmjxsZI5tw15Ufasf54SbxOUZGBSbDcYW7a/1TWQc
ZBMcG5muJZKEjyifDsen/jeAgWZ69aBmiCWrQdqqijJNj+nmsSkBYur/xUklRDWq8chLJ4NdUFxs
XrNzIhASWbyuqk9mcxDmbE18wmtSdAYeErjcMMm5dsKKk5twRoW0/7+QjSwNZc+rhrZwryBFS2Ap
WR7CsCSm1TSY26br8yz2Ne52S0C6+dy0qdy1Y8ivmnW1ZmjtaqUskqM2l8+Xr2K7PcyZzTzUh18l
EiSyC6sfKyzYeiTdmdyOCLjM4vcoWyvfBDsgt9CSwWu+48ZJh4Mk2FdMDAnribHUPuWKhW72L+ub
S1WAqO75J+7sgZyfl4zFPHF84B+twy3OGoFNN5VtnqFoaw6FRG/JMkdexRY6CMEkh+BTb1fn4Rou
xSTdARW2BnOSAnnjlsxCv410xl9vx05SZROjp6+l8PRGrErb3tdujX+gBM0zKrBn6flXBlhAbWZt
U+rA2WKDIYAnDB5GgPbnkEj+lS8bhN3uFLIE4YqnmVqvP6nbaAw26aCDT8NiAek+7OpJgMpIORz4
KFu2HcluWwMa/Odv4CQbO7qRf7fsIl71YP/KT9m5ladit4GOuH4GrQaEnMs9q8ahJ66lCZXySDNw
5Wtngu10V0p1aCGvQz98iwmlaqOMl9O/kZ0Q3LfU/w0iHnG+bZWfufWe0p0XtUYaunx+dZzvU8zC
oGQOxj+4c+FD0ml507twxzl1HMzIWaAa1HzZFiXBXOCBIOXNso7+oXp5slA9IeHe7K1r67Lz9+wJ
7EyyED73WfpegR4OacELeonEQ6Nc9C35+SjmGzyqBfroFrRp8IPPwlaqxKgQNXFUj647bavn9+tA
YRO7qId3NBTrHCfsqS+U/snoq+fz46+sTaBhDiifHlp5kY/FqKoi/zq+HZizLxbF9x7FwrBl5v+x
nHYxuhj1atLWUAMhI3tcqFXL8ip8TkXImLTV+X1qBdAbnFFZAy6SFtjRnNl8oGhuajXEd9uYs4sv
9AXNU5xfmnHjf9p2AhssBigy+0PK3l1EIL+yqF0HHmZm6Q/tiEP00L08NywVJiKHSoIv3urBITUB
1KwYHW61cvniLOykaSTOpd6DfzYLfu6dG3sAdw435y9G8NGFIsHlDvNfwWAL4rBq7S/LNGj/x/zu
h0ukXsWZz6WSwfSUZJyaFC6Iembgd4qsUIt183xqXOAcSdUO560l/7uXfFdUYMDCFQ8tVQLCJZgW
RoZwZ4Ni5/drdAOMV3IDZmaGh4qF7Z/qqBzh/Sn12hrR3jZuQw+RDmTQd2lch2w33HdI70ZnAyoD
GOsX9u8/3LfaT369eA6XAgMpea8tJq3yzWMYOWCUdOL8TAH3+cOs2m5OmJKr7V8BT9vbHap1X93c
n2cojqU9WxydEGOBElXgFscuSDRwta+IhAVD5pBnkdToawhjjq/zmASUcKevJEKaqjxuiR7yVI1D
GP2rdn2/axDairMVtxlUwhFIAYgFerw6v+DjdQShvgpaoyIVZnal/JbqlDi3eXey0gYnRpEBDzb5
OocQhlIP+tpTlcUzBV16QNFScvk0NYjZzxQ2SGyJyW3j7S7ssr42F3BxxviWkaIcOATfLX+zYzlK
gmKNvPnxRxqIuPYOPUZk67kgEZ31h5nBw2hleKlgejtHcIsua6JNC0dcak16OCAUgSjdvOeH7JrB
JDjbLMdFSq592iW3a8LRkO9bZWP8ykHRBqQvWfbMvz5P32Uy8Cvnc5nNZbE//pA5hZqoKTsKLdqO
MS5vCTybNFKka02HBotupmtH9grsnSEHPyK16jwCQL6xVB3EW/YQjBCg1OAX0A8fTqTKl1lCP3NU
oxdiXrFIhy4zJW64m48aegICayiezcqwXqwtKzT7XSmKQRXz7FCvN4sKYyfPXQl7NO6d055r/LLV
CGmJ/1haIMy/iG5xmbwn8i0o112nwGfqwrEJB0pC8ogWEs2Y4o7jYbzyGMA/a3BADENlVZwQVbnV
xHS6beK+H7hX+guTPcCagKbaYZyCnqMa5OXpdkmuMgRT/DMBxi2PuGd1mI8ow2js9DWNbYo/7gsN
TdEDwOhl83NbQe7sZ8ngnUzT29I6RIeMokwYOw7sMkr6gvzvcbmwjlzL/GCvKn5k5CbPlhORfSjZ
fxnEvR08IdWrWQ+FFKcy/BHXf2Xr0qq3ziA/ZF/vJF3AmPeOXeYPInJJwhoYX3ERwa7blVOZKePc
Gq+W6vIYeRGd4Lu3HygzR+Tlr9jGQ5MCsSwWizfz3yBzWeXxiTCReoRkhQiDWFwuPeRqzQdhybwQ
X/xMNSJveHWsL75fFmI8gMsjaPAEJG0HkF7VZQr0Mwsp0Uq18VTWNRSGZ/zqkvdirAu9Hxr2tf0f
Y24blwvAu5UHTy7DQFEXXlwolhc3HHlvBsBzGgetAMsAzDyWw+aTH2L64NaDBwor48Yuh4nASruH
2mxkNQTaQBQqEJ0SZ586gsAVxKBRUvCzLmeYeYRoz82IOAmGF+FPueaKu3CoqSCqW+scEWG4dEEM
NZ6b91lcRHiqKXEPXJCLxRZjtVG0KHP+KXNr9V6lGiZB0JMk/JuvpNF7a5qfXO/jK2Gwjw/C6+U+
4xrDFZX7F4PZSt01rM35Qx8CXzCEL+M2V0/rjYQ3ziHOhRjMgiPdEioCBhXhuaTEqUhAwV9TClfY
avy0IzOFLxVUip7LeNC8iL1ZR199ABDMJ+H+UyVUuTr4xlEmFABF/fSqrirXl0EggLd7Ep/2fMQw
pe4hJ9Kkci9xct5qY+mRKmYZQrFMAT/AJMya6GiYuLO46HT/j8jucLJebxyljqZ5WpX18kgEDRqC
YSouya51o83ZcpLjBlrxvUUxfI1XDf/o8BDC9AWQ9TAReAR6zbxK7BIyySpp2cDBCR+WQZgwo2RW
Yas89jXzdqTfOEUmxmxtSQVpMLmzHGRH5nvAojeSnlax/NQ9UwALhTbxeb9dxFnhILLOOBHKc+96
0AUts802g8OeyDvAYiQui/ZZfpwJbuE4QKW1y1LahXtyzFVQI/dkHtw0W8UjS9Xb5bgvIyfRy4Bc
1IntGsdh/VZUQ6IIgQkYHNvxXlmI2/48ytUz4GVnmtGweOC1RPEMHcPvyKKQmRVMb8o4O7XbBBVv
ZX9t6Sog7LXsbYcnGIwWBjT7B7unlN+1phjOHMI3tYmvyLJjWqdj8PqSxWntIaVItM8NJDRC7IFP
rbCGBvt/n5PPlVDYmnzqoD4N/bU3Ild2jJDyulgaoViCfhjed0Val0/OoAtb2RvdzhUTm137JLyO
VrQ5dtYd05rizQsckXGyzFC2194HpeYeVDdP380t+vJY3MWkMtR+kth8SyjkhaqgWO6jy9Q0Bh1L
8uSD0UCazJaPvN4DKnLgUKFEqLctBKY3MeqCt6dTW8q+mMzDxcBbyGdvLGc3A/3tNSKDcnaQeIXS
z0NkYTkO2DfQfqAP8+TrS1nl0ROTYx0ceqswRBorRqEzsik75ZFpgdsJDqfuXUX1BZZQqZqYPNGT
GQoceSjBhV2MCRhwiQWjbEz6rN6F4AO0QaGlyxMZLzGMsg/aKR0MP0aAb3ZgPzUVdAjyYiXK6/V0
WRkiSe4PY+PsRepjAvzPRyvLQZWvOdlkzDBjlbfhBDJ0/+Qzjf0TFVg7Z6jz5Ak4l+oWy5I0UQce
biBClpBjWTZfW11P9mj/X4v9UQscnU3T1U2UZl4dwZtDG1DebhcJwMYUOui6xYVpJqZl5qkg/Iq5
zmplBMsz5/AvEzgO1So4lLxJAedXzXJZeGtG/tYIaqdt2nAsOZD6lXrN0U01d/HCBxxXdul6Rly3
8Wz7G0aNUgx4x92lwyQSCqwvOm/0tu47tOATwj5co1nqNfLRkPWYck+dvWEXd09n8BZnU6D59JY0
Ox/Wn0g54EIfZte3+fO9DNyCT/XkVjPEgf807YGs9sMZogjqJlcjS20+rGHqIE56wVy3IOYnO1i9
3d4wfpk3N0DnpT4XReezTtd5KWvwODDHuZCOuvkxF6qwDswocEqgpkUobVZvMDS6vSbnvYuoqrEf
tinJFCvfJOaoGCV0vEwPWWDiQzJxWIElwXSvXI7ubCTkUaxBnIhotRrVYtxCT6ICeX4v9/5m5V1w
5xVgsoXwTpJxHqu9k8Awe+tTz4bvINzwKsN/KYrYS5EX91VLRJAf7jByE0now5VmCk/A2S4qOhxU
98Y+294AwJg92GfhzxA4zMHEeJ/kxhmnAhWbi4HfJRgQoC47F7FYWHsZyyeFHT5QVhcgB/0vjjIv
QVNojEevnaQZni5jAy8S/BXNVVBkpfoXrzxp9jJcWiYImMh+ztx2ndU+4Hjn81MFaUA9Of4o63cg
KNm48oqpeCFV/ZvGsF6FnLUhsHfngHQV4jxHTmUoLon97WRd9Tpx8Mmmv5eFidQhpP6FZkFRseI6
U0FdCw78BkH06n5U17MrtuyobzWCaZiCH/PRsArvOZNYwJEwb4Yeeq640DnDKIMPdJbcFkFf6wWl
PQTKdEeUr7GR9BKHjAZV9h6Ty98TSduEQprMRXQp9rJhddQ6iKSyOYH7BtNhJ2N1Jdsek7i4L01t
WK2fvuCvtNvU6PK38xtq74hHPSRqFMda6uE1Sbz0/rM7NnqIxW4BDxSBSaZtsoOHxXBXNVve+pAu
2I38HqkgGkeJE19L1cTAjviwKIJ2gxTzqk3vjesNu7P8/aNCVYxx9V+vZWKCRSXCSj028SX41KWg
/pGB61h0agEZjqqSdMdJ2p8paPxCvygXOcbgBI3isf2Ysa6AMdYnlu4P+lAlkMniolA3qGCzIEEo
6RBrQdFw7VW52GoTBHtaOHzJDpVBfmJJk4AGQLB6J8SutFduE5eAqKaxElziAK68c/Uc7l+SeZ3e
yTVBUDtlGM4DfelbtkiDQuNRB7O5u6XS+57Y4fVZvp5ykLrZqsJwrvx1Vd6GeTEla5q/L6EcAXwU
6bQ56hsFWdUT25EHUgPqzyWRAs4n6lAq8x87F6lmT8/wda1u/Rp7do2HAz7Wcn4kRY78nzG6g9yd
2cG+ThrOPTED1/QFk8GgbVfAOYJGZfg2XC7vsfCF4m729FozUcYo39Awx06/ZSncC7ibSoTR00IN
q+YtMd21ec4f1mu1qtr5LVZ4Kv5yoEZ4A/6c634TCQE2JcsAqr2FikZpxhguUl/M5/VmstqWarg9
P4oldz5qzuggy2tUXvyfhf7wsWYyhg31a/HEIwEnENake4SkI2Q7HLhmtzSo5Nxq+Dlf8DcK7w//
cetVmKhlxGy3o4r0ql72+O9uiw3BMXf1YlJ+Z46efoHIw2eNQcNRBuOEmydjJEMYvC2IwZrefe3D
pZY8WigcW5e+r2qJMWH9vLWLWIB9aSxnwWYZpQeiPWp5gt9RSFu75lwU4xwUy0dlJH+jN90fqOJ0
Jl6DG73reDabKrmEc/aZqqs/s+Kxvr1lzgyyj6H5kAS435AYtMz9xEFlP/VysQ3sNqPKgPvBdJD2
pW2/UdcQLlX4B+t6eHQ5GH+qj58vdP7cDZAgmGR+G1kwemKM6HTp3k9JO9gLeZsPvM31Iu7YNGT5
QlVJoApnYj0WjF4rY/2PhF9M8X0sRLTjK6ScJ8TRzS1Npfwagh9hZcJi+0ptt/lD79Wr0uzWncqw
muW6OIowACxFVZHxo+NQwYAOUnUhX50ga5r+oAeX3VZArjXjF5ZQnInubf/sXIDw8JNcSpR2mIxB
K106huzKGvGDh9xmHquACsHT3U7kZW8yZvAZ+O2xwYezvaHJwaHQV/R4HcU3kxPVIT8RjZ5K24Lu
grIwaCqpgtnqTfjF0HMTh6p2XTjnAOwZSesEEC5EaZxo0NlBDWlYZiM4Cj0P63vfY0hy5+4JVJ/6
5JGiCZAFOpeo2Q0537fcCHRXcpi3QMjaJNOfcDU2aVVBEmZ57zLM8u11Q+uUvPYdoyyZWnnv/5ss
M+IaJIzGJfIK787mhBo+ixwA6qsR1ysLvDN4MiGerlUpg4oknvH5N9YIfMAEWVtIq/acGZNJCyu1
yFPK0SafOdvmMUyetPUjVM2MhzFkvr1Q0sDsrrro1M4L8aD3rjsJl7L7EQHuJh/mGulKKyqhvdiK
pCckuqTVG7fvzdhmad/+bH9K+IKdBjYiSKfO4sFCfpSJTeY0dEK5nORqO99mcdYeIcnR94LLa1cE
Ujrrjiyfxa2V1tiru9JJP8WSjJ8UaAlyeve+RZsI+ehbA9U/BGRCBMJJDaQjyt1k3lcZjUG7RLi4
0GHRtZ4c+S3w3B4XcJJ1JnHfGKzYvA95THSurV5k1V7EbCqNVsWfvlmfN5TxOZG548vRxW6DPrHO
ySJlc18WltxCQx7pgvqxtoxmQUh+7bEAKBQVvbAoDOsduD/khsp24e9WAFrQ9cbyF7rsHCPCQ3BP
EXWy9N0e/WqbEvO97nYnx4C5nV1L7WTJ9MZOFFsyqMfJ1X0fJVDFz0ylDLoUWz9tjO6IoleN4Bc4
rkrf3ugiVPKXHZNmaYGgnQVBtvh9RYGFhCU54XmLnSUdVj4pPP656qHWBk3w+TjwQ26idPB2MZIM
JiAXEWLZO5F6N/5XiyI52lR77vMzCphFs2QoUwhK4C7JNMFVazaaO//8V4LiGjHK6HBdCqo2ztbC
XcPQW+aUa/944EasxFBoADyXoOEunqmi4bLy2ktolGwow803C3+n+sBeUr0F3D95y2ik66ENN/cK
b85LRGTD0AMufGtNi/n4m3+Dfrg/4Mpcj1SMOLC4Yvs8EIzi/otbBdgcEBV6/tgjLX1sSCQt8v3I
EJK2px3Mu4kg3/zGu/A696Qv6yO5TRHoLVQZpMoQiVEjbFinwn/KGtBPTK31OVdh7V9LeZRTtHm4
lrAVwWSXTMGAoLvC08j/wSD6+hb/Ou6Ni0bmuNoLKjyWiy1e+3PGlmmGE4ZcBYcOED0szI8aCjnN
AdAKL0Oyl9tgVI4w37jhcOXA4xlK94NAx1txCzSAm1gQ0gPjwBCM6307S35F8/6MiUYSzkfhZaex
oWqh16FAUj+cOvI2bIFM6VFDC7s77FdzRL1mCJFo1BDa7U2Mr2DiGJMCmHy/H6BCuYomdKk2yXoa
MuDwT3Lha35oc+2BNR2h0QL/8z3BrBKSl9ILKAZLa+VwK5GdxVtBl5oF4GhltiPE3gwC37PbmSFq
AilKChELufGe9BFOzNWjWpdCfovhOhucxJWDcda8hh0OmwdWsLs0HE9qTlsRmKIyzmTpiaS2QEpY
WBoNCViCPwUpJA21u8oMlGBWjqNzeuksGcttHC0kE4ltx9KNBhpw8AqA2ZuKvtH3FswwSj8BoDI/
so1Giz+y6KDrXRcyF4mMEHLwt1Vgcw8md3lYPcVLK8i307dWB7QkRyBumeVJeRQngUHhJejXFTxG
ofIhVwcUa/8r+Xtqa74nCs3A1EtJVa7yGR7PbVbRGCOwsaJu1G9wJ2f8sdcGWn4ZnsJYVulMVpWu
3mfj8ZZpYKTdgnUCVA13dfCr2GCsGoTV105dZA8Zyo8PC2pFncykA2stJft/t2+he0u0lax20BF/
kOJw6j9TZdDCGDgh2HhSJ2SSijX/eaHOGPIBy0PFlOaUINlRDeVumyy3zF2BeJ5aO6m/dcrvOVjL
hXZBXt3Dj5ZijPeACZ/lhu43HgbhZ0Dd4+IzhRKiVqs8dZhAFakt1zCiyMpJgjM63SP55nKqRjjf
4GqoB9+HcO0uTva3RZO5T6S3RPmiY6KMPG6LTm0C5bNAHtGcMIb5wXXshxPvsh2qgcCvn0e3QoAg
eL6Jz4d1Z5bMAV7ysdQg+B3h7pRCqWgjTFODkwlGroxvoCl4vhWKBT4eioS53FOw6i20+sibG/ca
sQAH8mUy8+jMl0t+zBmHUc+/sNqFEarTpgK0JWbBcnc6tfgUNrevoFqL80gZxZHRYddafPE8TUCu
wBXAOIMAvnf+qxWPscAsALtREUC+ac1PVBFcYVyo6lvcGMq/7DvBwqvDHTfwj9SfjbKyP1qGWjU7
WCAbf3UKr3QL1T8S4SThT1NUHsMN73lzTFqsxSQXp6zu+t2WuPJlHIwkvPr813XroEo1Dd0YGPdg
AhwCxMwSNUVZuh5oWiAqgTekpuje81lAjmXb3tu+A5JM7JjChO/U9i0I444QxoumbNCqW/6qruwx
4GPEQZVk6Jm/TY+A5eQdgxY6C89qai/P857KTOYpNd6AGjjVFMwZpaP7hSVy5PB37zXtWOp/foFl
GOXYPPAD9s2Oe2cdRMvepKXijq/3SfnBUrsGYl8vP4/mOlOPulwkrKRgl28rxgVgF57Rnm5BSxDw
qfJE5aFYEq6bEPjh5N8LFproMvIJxPUKL/wl1wkJdN37v5dH9/45pn6ixcNElP3ZFNWq4+MLdQfd
+6J5OdmKrcq/GLnguDsn0czzAjV71ej5fhxFw3VFUewT4z7846V4s0o65qDbFXbJCt+cuXoLMEOq
/NF9FEeYCKjbbxhN2UKbT6A6OoJl0UMCT+q0jQgEAQA84EpZ3YXazGQDOVbFyjtz2/lxIdrbeRZ6
9CzFQHQkJVyYdGJHtoGw52ZjFjSy8QGKeW8Lv/qy7gsQFyCnHUFOLnMUnKkyh+1BALI/OPKTBjPZ
WyqQU3YsU5tXCApnOkypIy1pLo8tH6rUIJ87QtAwB6PhlcdlvTJjxcIUz9DHrZpQfbUp2FEDYh38
zWFWfHe65GMFILKNmwqVIkXT0IOMjWsK0JmJMzXx5SOChGTcaYvS/LdWMB4DW09i7nQMvKAfAkpe
lRlER7ecUSReuRNepNYu3gSeFwvw+sdWLoY0BCFlCYNB3TjmwcHExt5+lxx31E0NCIL5hPcQ2OYA
6S49RSm7xFHfw/Lz7Og7L7F7kC/9f8W1Sle3YOjwAbaZJHvNfnsw9GwzC5YQd3/z0AHmGhStIb/0
8cTdMmL6+opg/52QpSMhEcNWvJKpSTIx7NfQ0KrefChexR7K9gnAKW4gylEvBVL5nuim7F51dNfe
H24rceCTWOZDlD3vCufQRFskONXa1Z7UoLM3B5ZFVW92xxUe81SiSJw7ids5TjyYy5wwFlKuwjI+
LZuXBsQEuEzMjqzM5P7nrsRZvFwhqotDEnAfFv8ViCfmRVagN6zO8z78Cj/+u7OauypHHiZG2qkh
UQB19wWFnjKc4/rDl+b86Xvhc/IZr5FLy2nZbZdbPEb5UwrObECBErQeIDjG9YrceNTm0RL5POH8
Wc4ad1drB6edsaJonvxa2NICrHR79Sz5OEKjLHSr9TtjHjvqY1VYoYnWjTc0MVgqzdCBHt9kVxIj
PhmoWe33LYVpbZFSL+1XxGFOst6qJcWnostlRWHkGt6gcV8g39URTww5uPnJ9S/scRlxIOGkaqQS
goTSdtHcFcTUPsrinaFbDZItTk8acwT6c427yyJB0wgKjB4oQiQsEAbEgx5HNRP7lvTaBfIxvUmY
dt5eXgloeZgqoyW6Jc0EMG/SV0T8FGBdyRN8gIWRvK5qMcNxWBTBB6OhO/IxSOmgB1gF/DLw3C9u
wbF1mX3xG2ZHD2gEtn4IWguQpA4AJ3KuDt+V/QuLthdyQ+4jl/ilbOtizqsL1yEQ9hG8egSjvMFT
ELQtDo1EnkKgD55k4zOKk4DA0SjeszLJ/ddjRqFY3DkWXGrwovhpSgrWOarja8X620iHV54aS96/
qs+ORgeNm1xI4LmXIm8b19uFsqiB2eYnsoFv9iR4Pe/BP3fFeDxHiITCK0AjppvXGwK3ycZi7QPl
J/LiJ6VJm5rcgAnxOe+a3iSQLauuo9WttfTK33NJAeX3D05cq3CFQn7ROQnCnsTh0AXDYGAIcgLs
lC7yPJ4Pyvux/L/nZ7le1GuL2cxZJQ0nWMT/WslwJsYSW8VX8Nu6WLvhuFwyS0YQIAW+6AR6HMIT
/QUD04a+/hPSN+NGHFWMJSFZutTutjVa4EeptyJYrbKsQEJrUELA/+YX6VjXnPnK1/CEX5kMWVwb
ePm+VC/Pq0Ps1P700Ppwr8W60n/Nt4SC9mvQvRAFW88UIfw/d7Nl1Mwr5STaL86ZnyW2VfzwcATc
5DdnRxzdG3zDQkmF9eMqBX412QQXfii+0GIXOxmgbXsYjAHNtwpcKhuCDKIlr1o4rEGXd1WeLeWT
NUJfP84LISH0p49HVCa6cNnkLu4Xw3iKx8mcOsiRaauQepHQmKaoYXu+W7B0QqnrIomBOZAFHZKA
BS6SdrnIny2fkdwWd+f3gHp83J8x9V+1LPYOGR5lEOa53QQvuWzNxTMk1L0vypgXy8anCvC2Dtxn
xKpwzWVOrh4LhuYxcQXLemTy8w2b70Dwl1hH2cojoM8j3jWYJfuD5XTlCsWTrii3KxEuCvYVzI6U
mvsjAMA+d67TMaBBGeqK3PJBNwrH+b4R7zlBQVox5yJs7v+O0j0CCrm6OqsBqImjFJm+gdFaVHIA
FeVaJ9fpwphiBo970K1MJBM91yQRpczxOpFgMLU7P+WHxS445SvV0SuxS+SzJ2N5LGcn4nKBv4x3
gHfyr/DEBw/X1XrbmlCu+7Ooxtnk/95qmAi4A78GMRXO9wLZrNmHBkpNXwlfikSe383hVTAcQenT
xax8zXbZ3OzrwwIqF5FvHKmM4hfPCw6eZJdMbowYFOfIqoBl/QofjINLVl3dwxwPm5Tn3SbGKZfp
ubX40QV+JWd3lUY169rKFyOd07SRDERI1Ha8qSCtNq4Xrcnhh7lYGDLdy6F3iWNziPTnne9r08IP
zS3JHxnFvJXH0k7xqa6Y9B4cSN5S/wuwL9kuhGQpMkWbUmwaY2sRqjlcxsOtTTfTdsyvVzkwI3jt
ZVfEvY2kDHGSpR+J8i8QzMHofK8ISGun4wwf/iG9N0Tla0oUNMpdPiOZfX/0eh+bUhkCttIM7Lb/
fJTQBYh+Icx8jueGDSpbIpGDcF9mojcrkzGRh5EvU0Wl6DBQHgde/HXsOm2zEMQqHlcgp8Rk+Ret
Ri97tlHydAny8oEQzF0uSUYlMQT+1G/uueZ2mvzYTo+WmYcv9d3LxrHqKkEaE3eWKG+Kx6g3ny8w
9uSLMOeuQ3KgG1addg0Q2B8DChCEU1uEL+eri49i3kUetKv7zpyft0KWTu9GEapMODSdMb1sZG1B
hXNv7a2xU+oi6xip99cCEcPCEEvDlwndaIVmKsGdzOwmO31POCrKz2N4tPtGMGL8H5V/GhdndniW
LMAByWjH+7N2y2fZWfJsvKwqouUpkVmu2II6ZqIXeL9/wmlq+2Op1N1H62Qv26KKzWntPMO4rQD8
nFT6m2FNGyYH4fwAJDTY/7NlclQGlHJ//5dNrSq1DKEOHmthmfQO4MoTL3yPEuJWXllLqp9hRpm4
+KwePlUEgkte4Gq0N3jourlNlgcmOfZrdtbjsYvOHnIgLtkXL4euBUpnDMNZvkl52+XNPVBqpIfI
h0/jTYBd8pwvqI5eipAcE4DfEYYbwCR+jZADNNsVBHAjgprHVf+Ct4KFOFtnRMw45T74PLN5koNW
815HNx4vjdQ8L4cLmDUMOXQPwmukB/JiNDtkIMMZHEj4KDgeX/pPN/E3kE0x9u0FECkanmEJ9I/T
SJySFxVfDANJhCTB7pAt/2gQoHUa8JppAY9W0scuf+odb95DQ6dIf0xgGudkSkonh2CZpE/oulCO
SarQlyQn4ZRVrjdntOONI4FPgVt0CXOpUyAiin1gooNKoRGGqpHopFSxVXzCm6b17C38jv9FnW4Z
gs01ITK8cXJTF4v8f/3Tcuvg8y4OUgsKqp2LgHYN3uZ4AHMjkhYMEd9H/fhsJwFcTxqaylsa61x1
sDR8cdwJNcJKfc3akIW/szjRTIvj/XxSNMNvCSXBnEbIATG6WTU+/debGcMfl9IN2KQI/roXL9nx
PMEvpTsPh7DZO2ieVH9tGF6Tj8WWHxPBlVnBlrnvptcZ2aC5vM253lRzE1ZP5rCmMKxap4aKK3RN
EAMSEEOMvYHIS866Fys6+NjEgbnGx36Z80c0mzkAM/H+blzWZp6koDj0JmdKLROj1D9JI7Obf0cZ
7g2QPwPDdh9FQ91Ydpf2Kyb0lVB2UANgY0PIQQeWDzG/+nYXTp3kj8mGWYfSbYEUBoO70lx8C1uk
aQZ6zoF357iaesS9ljPvz/5K32zk9Vk45d+r9faJdlJ8kTd8bqyNjBFkyqj76WvfOEOa6+2H6JEb
zNaahpmrIV+DU0quQN3sDo61i0s35EOCNcmiKzAsgYuNfzb/zWfnQwwG5TyN57NSc+VGQf5nsHsi
2EovirOghv+B3y4+imFXN4B9uI7FQ6T4PZ1C8jML3bAuQhBx8bVQSGK3sJgToqes/pQc8rUnBcJx
HHWPkLfAeiiDrkw4y+rW6j/0BKsjL81NKFTw/4wcvgPkLtCFD613VfwqRtxPBJD4HklcfAY1GvOm
5Gg0fMYcTzQ05Cxl9Mchbh7lhTgptRZvtQ0pk64Fg/ZbAZ6eoVqQRrLRhss0G1eytU9T9sQQyQdb
FE1qre//h6ZtMN/YR5p88QibwW8qGdylEX3rDGzfgAnNDqtiFyZNv1yZd3Nxq0uxsAQLn8a4u5e2
FwN3R9lxmJrhfuev4JhzWCQVe6XQYPGVmdjUxNYUEW/kYdIxetfcBYzrFC602zj8m0LHtylnuNzc
TVNzpdQTRqhV/eOffU2WKAG9iUKYU/uBg4SFjbskhF6PBCEDbdcLUdqcSEVayRRsS8DKBYhYQAKL
u/sxi0K+AoGN9MyqMHXLLnD6oRl0GA1O0cglFASytB41pIBr5UWP/a1jmiwfY3yBLTiXQz5R0+3r
GuP1UjGMtEblrmPuL7f0Z8x70f0nunXh2aDa5lhBaBwkSKv2NrRnwtDGxRCF56/vDNpSEdgWenn5
lZptGr5gNYQpK+0Q8voh0Ub7/Gfv05yGI2XkQzAz29wgzFvLuxdkHDGj2LINmnGLn6gYBGPeJuUC
D1TvPgsY+fRY5W/zwcodGkI2x3UdY6lguLRllBHlABxLyqHAuU1Q+D/QW+6vvKQBtV22//m/t+U/
JpXuogmzxbuyC6bCJ2OlUnTtBCK/yznLmhfgA3rZhbULLfoNTr652EK/5Mr8RxorwlTxd54q0lmK
kpEMbpZOY9p+xoH59cWiy0xUjA3F4E13lC1aPGhl68s+1nXXunDxIehug5zs/J/s/MIrauKdboHd
NBA0h0V+qboZFmbmpU79HboUjE1BBcRfb1U3ioszMz0Td3NoZnmGOzhwlsgk6vaXfZHatR4IN2En
1RbIXABzglBprPkkmE34s9YCAVIatr8gI0XIaavOCjw4t9ZNv+zkc4ThtNAhifVGaJPxQnoMvMwd
8MJIaemDu8/lBHbG52Af1Mq7uQsPbfJRcMK4TXiFIn2EhMTTOFVxOA5LkizOsGUiAjJdD/5hJ3UF
IZEI/GksJawOShOSFDsUmlOeveDXCvV4K6VLT6kC1Nj/+qRZf6HFhj4MXiJELvBXAGVsyqXrTDU4
KlYUgF66TFEAfdF4cc6ccGbCK9kOT1VjC4l4m3rWw2a5lxMLT6Y/sKhnMrKV1YiMmHr1ZiBb1rAm
QpHKY7BZBVpcHp3NtVaSAhfywx+jueWtsNbOnK78sEbjeO7gCYAJnncTwkB11Q1u5sOLfXhVMO4u
ExFLrGK7M4qfNCtReOGOtsWllgRjkbPzGOAe3mipwmYn7unF6vMurSZEqxPDRxkxxK/o+InadPA4
pmidjIHM9gKWRaEu6rLHIVB8aJV0quFR0kyRme+A2v7GkUW6D0F/5zV5rER68fsH5Ssc/5EBITDH
+4OL2mhD0AFYxTdTQ59f51MSsRGX0e2ko6+jo5A/h7yyzNkxEdQSsUVTyl7x4y1bskPpauf0ozNJ
nAL22TC/xvJ1gOHXFEUJwIPKfZEZN+lAzwVTULRvwIh3DeTxG+hOTZIY1PQlCFo5+iDgtKty7CEP
+vLL6SJbzS9rHRYL/5AsNRDZFF6V0pNHks9+sBQ10vzAX1bixLXau9YwMlTO8k2PvUDgJ2bvC9c3
ZRiJdqeGKWW0+MLbOp7+TuZNn9miA+B7bIIrrYG9HvHfUphnHNl5dvgl4To6HPkWT1639TjMr/oU
qWp6pp7lsuMsvkWiTTj5gFXeKAWxQ8ECf2awoBDkWF6XMijL7tiOIUuw2JBtIDaSsAC6AEGvrlkh
du8PKhXcGb6RePYgw0CwLSKNWEDBux/9QjcDHP5W7Qqhj/VMx+yY+5g07voLbEQagFfpAbX5jnyW
hruuWMJElBMsMLfqILAaAwxVfQJ+mcMytvVU4MhC1V/AlSVekpj71UqrLNUEz3zj1Oir9xQladv9
/b7wFPhp/7E2eWUHViayQ01JnnSk8ykz+T1Rij0bWZ/O3UNCHIz/4cwlES21uQUtSf3+4LyVpD9m
d/uv3mxxHDRcEAeRBWb8mCNvPgDW8O/kbUry9sX+BgoFZiskZXcVMO1ADEiiYWCGglnvLgXK65QK
oX8e2Ll61Jald8UyCUbqrPN5qtqegFcmkyAsqaQPgFKWkWSoLimOXrWoX800BJrF+Fh1yVFK3AeR
/nhyYjT9bIaodWrq9vjqGDLo+ZVaX+9Lr95ViuM47n/ZHeedPfBn/w/om4EYsmDQdtMRa/mKYhMJ
gwB8tgLEye3liVNSr/Ym1tE28MY3/jT46vAsUGnoFphj4jaXJiOxT/4TA+PUbU+8MDndpYDGbAEH
HIe+R0nn2xfZ3SZyUVNh9cyoD5aPIMwfeSBKvirJKqC0hgya+pNI8R3ScTDy/i7vwZosi9jgRrKV
QX476bOZtkP+Yq0fWXOWN2hJdyXEPGRv/PYlkMZwjX4alaKgc64/sZQJ9sXVZJosOKhq+vEMGdiv
UU49W2I9JOcfLV9QIawBque3hl8H8z+VDe5eEdbsLiPP0NM1jn/D3HVflw4ALCbtVZOZ59ih1bXw
sTW2HRw3eKRyfKi9aySgPIOjyJQsbUKqM2qjhqEsD440Kip1+fqsrLIrApveeLsZ1K+RHZXpEHZU
/TTayj5+341W+ZqFPqAippHM5RgoL284Anf6bmcmhVJpH8kDrsxP9kmC8qIhDtdX1gAuulcC/hcR
7eYSWf5mWKUiuilEFMtEcrXeesnVRXVL0SeMq8oODExvUvjl4Nhi5vTC8gkJ4LJt+gY/qJhIjOdg
VisXPWW/58Vf188Zz2m0uSDgCreTT8Tmo5w03KlhhGzsYG0OtcmPG7TMcIDRPNSe5NlYrvaWXVis
WmOsLCIN73WMDv9lCpFa8Zs/VX48H3cSBbvV+aZ7ZPkLrgLXLLTul7ZDz7xfgUVL/RNceCu9aD6W
ZLYESDs7Z/ZmIQ1Rcs0HZIwArkDrDmZNvI4nKHQkMTwuRbKA75A1BFiE2OqJ6jjOOLyaNwZk7mO4
lhoCgd9GlingfDaAJeYTXL5JNpVQbiUXWXzWH57dykl14bQA+obaiUPzf5NWuim438MC8gp+tuut
dW7Zo2/fAXbYD5LXUyhI9gAB1DUAq5spF5t71aTEHVE2wBI0X9PGJswrXh7H8AfilhS5H14fgGWH
KW1nzVlmt2jE8aACIdl3EMXoJ3JRI+YEhCtdR8rndZvPWGN28/hBRjb+Snvi7co9yZHjByzkTOAa
L6MKntIpBVWCStj98Z1Z/+H1nm3VF+YaN1NYmqeKuVruvWXu7gjPZwsiMyMt1TURLO/vZO61/0SI
sfzgp5y+VVLt09rSIwl/HBHTS+FtX10PRCnh86WzIyriPX360N8DTq4M5jT22HslQbBRK3j+uphU
9xdURMzdfmzzZkbpRdCny9TNr3hl8rAJE+mY5gS7kZE0SzWCsxIH5w8ECOm+27Pmqj0Feve30rtQ
Cq/us82I4L9+W5zZl8/hmCuoCMuAfU7orqwJ5rhwlpDevP1JCRKfYaR3nX0WBtcbn5vss++c1EEn
kuBDYa5N3h7WqMPImXbGlgkfkq6LKyWkFXks1155fg88nIi0ERUzb0q6o8s7wRKNLBgWdoCWYwgp
qEO3aTQCEfbAXbuglPTRpKD6dLI9meVn46xi6h24nPnbt5YnJY7JaWtIZyZMouG1cxDuWW37yrlR
qn0aRSNFHMTEnk3ON7t071hRC2U/DknJIG6erML6k2mnhsrYPBc5ok9yKrGeZwyoGBJaPKI84/UW
CyPrLgSKr0KJEj6EYGehqqqZ0Qi8ZekDs5taByOks50mXNJwlg4lceJd+GhFmjHnaPg2QGPjKTR7
xo6hhnn4sqdY0FAFXTyIT/sq5hcWtuA6x2lpTlEkaBj6loZADO61ZANcSIRAI6a0EPKCNNVKLn9I
AfFJDLkxpXfQhmioyVig+VWTUgV1AH6VWcxgLtED/xTkKFSRgXMKtf8EhF4RrWMwogJ6wpadMSBj
RcuBNhkPMZ0GL66gaIgXsjoqPHnEQ2lV4EGYQQa/uwFLH+1TXU5IJH9pceSuzkY7fMnNk7Ch7K8Z
RcMTKFMmTnH5P4iJKyL80IkJJIYAL3iwcaBvwTAsdIB8gtiYu1Qqi4+W5xHpgPKT6eigyf7KHhz2
zOB0b5Gs30LeQN2OATFbOFvXUTC2/AAl1Icqo/7pI5/86kdfG96cs0vaMeiy5Y4PUwFXPJFvt05w
sVMeC4ZmsPFW70bqZzFxlCmcedo4tjp6FgZPprV2hYbvjeMDuJGu4I+PCqsZhhBmWvLZprHvipAj
E88PvSywwjGU2W5Jc9FgRjRGK2kCSnlqk+NhT1LQMZ/kLE3s5IJKsufcJSHd0YNv2wfkIHa7OCNl
cBdjCMnM22+mo8jtNO+Hg5gCiIqfC3fiwzXx5cXgxW1UhKCph9UZ7Dresdn9pnaOxz0ZEgCzg9eV
ArsiX4GWU9ridN9n9sX54O9PT7ip6vstWvwaPeeVz7G4Qxjx2IKyPf1Jhb4e4xqdFMXywXji9jmv
rhktwRJpwT4uPXbtpFG++Qzqf2wz/60gzAYXlRr6J1YkUPlwjqdoTRej44SJjDnfoIEJNWlvKqdC
Owb71Ul50cIJfsdVp4OWwRn8ckFmDY30DJbSwWoc+TrqDKrF+ikcDnjjB99S+iky3bd9+CUF8irL
YMccby2PLc2Dnx0SDZycPpPbTj71F5qEBv0DfXD+cJVlOFXd4uvNi17Ng+jrru12zYxvtJlgeuFy
wt5QSmma1HdpWf3olhVkJio7eiI2lKeitE4ZosuisX6lvdrVa+0OZ3Zlv1cuVojMkVlFR8g0WJp7
X1rlMKao5URKJGpo3Do5BFw62CEPw9Xc6VFsTBaLgTk0hbUIhYZL8a7lBf0UhSNyK+xUTNW8VMSl
fUnGxg44hMKjkAIablHfdWjxOJYd6djtDJnTxVamAlxodOQ4RqMJlI+JEhY4c6w42FpMjw+9H0dj
L2a1FWyl7hIpaBdSe4AEc/RYRVgMR09S4CgKsWVi3ausW9EFLNnAHcr0gvEJUm8rnYOgAXxVEknY
xoi1lswkBaT67o7Rbhx5y125Hq9TzvYMmTo6+jdgKu3eF7qNrVtIiOYoRMdOgjd+D6ff8BKlegGN
axt/VwIpgMl/UCsE4090db/pvXDEjci33PVjvrqSDPvodUNaTrRk/eSPPRgHNB5utdnzopZskPpa
4DTukutHPb97zm3bmz4LZvEIHBGrido9Y3m/cijDHtJNVOAvU0JNsDoFk9hlRANp1ReoBQuqk9/l
kiQffSduz6s9u5lDipElOQN3CId75jUicjOPN2tGii8CSgAu5jJW772pNBXMROvJeyxsfG4y2vzt
25Ze6WJQQ3GBH4RtWFGjdbHVNoHbRLpHom6RtoGe1Fc8fdIRtyXzlv717vP0jRrb23XHXGDl5Lvl
tY6W/hGIQ1Bi+XwDKvQlwS2NZezUJXFUCIR2Mv/C1/isl7v7KsGyCHx1YHOAZJmE5WtAepbwQQ9V
8QD7vFzkrYrQGw3SrbcgQXrEbhbXxwv8VqjPcEALiMybDkz3p0ncxfhJiIzBHxcv5TsUsQ29egkw
PjJS7k7OSl8fSZujbi821Y/TRcUD7Locc+hLRXEJpMZ+Nw/hO1TxYG+COn4kRqaP33NNtrHrfF9T
EY9E7OHesyfSzV8us/l9izn2XkJ9LxJ/YeiljhBiJ2IQdRsDUPdq7bZcv4AgYRNyCp/hFQbeMnOd
X5hV0iNtQXQdRJr0OplZiwP/8hgtNV1/vGdeQioHBHta5MZKl3G7fNhC16p/vh/NBJ010XFvC2Xh
6wtnnAtIcYlpBO3jpJrDRmgYBXwTfQ6zcK/5w3X7jzwRU5OQFAyCc7bLrv/UXy5eBXZ0nH8DntNo
mXAwVesB6EtlhMS+Q7jcMiwDXwd/0cLt4mQiKWth7YKl7ypHuX7b596VdfD5yFKUPudvR3Vk7vvX
Tkw0pZd3GtIUWw6cU/rMTTFKcJyinOfZlfASxAUUeDDaTi+ak+OrDZ8F7psVrz/tCwYUyICoKClQ
4tYawZuXM/oI6nNoxDPaJ7wBt597eXa1e/zow/u9x1Bh8HyqzI7E39XTDTMtbWweg0wOtdAwQ0St
EKKkEo8s7Wl9xrsZ41iyBxACdSp6R1B+Bf6HUF1goi4EZtDW8j1lvGthvzzCqUhDbxBXHeYUvyXw
mLvWI2TynmwHgIYhJUtkY/0W4J7F5bWbAj07yTO+npIIqRHTlsbQ47C7PGdZZ6QJnnMYF8mqjdWs
4F3ulktfPiC4EVQCiAx64MtC3xbuc9qMtjSnkTLD1AI2iRX7NLZp28s6pNLDtZ58vWcFcqr7dyI2
eHL0uqlyIdYqeOstlxX42X/G0rVNJvLDIB93oqtleCve9t2Eu9cvY5oQonS+49eZMXPR/e1gCq7P
THg1qUVKJC/IG+fSsSGaQEUmBLMsmDlGqp9CW9t6aA8KbZz3WFEMpB1R4EnC+oEVq2lUPIP1dIQy
dQAXapSRnUGEzF7D6Yzp/PN3GMSrDERXlzYqw3+Ty38DxUKTWSKw1zci/FlziTsNzjx30hc79z4S
IS1qS6ywOIzOl1SGn7/KT1iLgXfgxHlI6IZGffI4Cw0m5/pZ14c6QcomXnx3IVg49dEVRlId7izU
fa31Eeg+NPo287SfdEmPnxiOAi6jp4YvwRU4GK398GFdHDr4lo6pueweve9wvhyiwYewvDY/tzrW
EmitG/Q8Ow5tCby0oL68qaAdORk1mt2zR5yylWXvxEUjNVjaYDrQqMEl5AHGbD/ceWIk44dvvRhi
hCwr65VqxOIolzsJMR6Zb9vmzoO3gFXwrzHcnz48jtAlyNrVHUU+4Ss8KnInZIZP11untohpqz0I
yLizOjj1cV1aIYa4wz3Ib4szEFRDexBR4R5S1umEasdt/iAP5iHyC1oHgOk4P52FLYYYki4NoCOq
G+cDkdIi4bNwcz41yfqH0nPTE7vzPihHZTO6joeG5Civ1P/8MfPhFp7U1qtkMYnvtmrCdGS7k/aL
O3cajBTdd9yCh1/genpT0N5Uzi0ooT8xCxQ1ZlSxWF55umlHNIcJnjHFlQocQzQ530u/xDQ9fUy5
TuzfH5g9YrafVkWwFbG3MRUResRrgAKqfJNRWTJuN56V+rRTzojUppZwLx6AUz63lzYEd5Z/1ncA
e6Lp/bDKrQZ6br+CTNdcSKub/7eNIl6Knpocjzz2Ui2/f1Cze6eKYruA3ep4LqNabqlysNIwJw1r
JUe/wRlfTN48maMRiHjj1BnDvAKWo+iPym7UDcM+ajSLSoLoitZzQIOnbW+di1ZkXI6wj4IAZkMY
vWfTwUTNVeuhV2GDYvHFyQHBrGoRH+mIbNrbRGbPAS0YujhKm+pWRHi48rLgLrQTS4Xe9x8+QbUS
YjhGE2B/BAxhEjhPCAyJUt3zgYSPXChzhcK6jdTegudrQpG5k0OGe42cxluypE2TiNsZFV8+FIZW
U1kpnRxGpDV8ETL2Xh7m0UxfcX3O6h3UDk+1lBdzBUAy5yvIKS5i8rKG4Vw4iv4QR9qPAyi4sEaE
l/dwSEXZ1/1EPQGq8eihzRiSjvOKefN3PlS2gvVZ2rxNZ7hn0hszNb9qfBejMD6dFYxdaoRd6hM4
RvDpJQGaFg4DK4jGFN4c9OsaMrU2y81tDkuv3/ialc0d4JSJ4ZtiQUxPh4NIVWWH5ImZZmRMOaGk
XC7WrMMBkLF/U+2d09n7Jnizl/hPH3YY+nFXJBGgwuTAWYKpNIP1Tbv8dxWX2+GXrm4XyHecVgyX
ifN8txOW9wcW5XcPjOSSEk97+wTomXPmBRmODllEq6g61Ja/0Qw2hevGN8bsbhD9nKtREE3ouIjr
vjuY5J9qKGA2UknL7C03gX6xPMw0jPtyGRxnxihnb2gJxEEmGm2vCkKirAAuotQ7X93H22NHlTjV
5ZnnRta4mq0VGXyxo5C8BfhjDkLGQhl9xNgGrQOY/vAQo44bmyixn77txfbeGj5bz1nNpMxrQnQf
VJSYcd1khiYP+c4y8qtADpAcQX8jbx0nsHMDh+VYug9MeTiJpcqEFmR/kePXr2sbxmy9XrvT7gls
mdmck4ViiQ0k6CZi9G1S3Bs6lCkp57oRnvlhSUoUr/gEU6TkURcjVuqroAyCwMmuzd67hxDAfBxv
wqXNOl1ZPfowPZ658YaYGIq/mYZExQv+BCVGAtix86790doLiKdLdf7nt1MaG8LMFiaW8JeT003Z
ce6iluZb5tIO/POMgqJvQ/PKJ61uRKjvcpwrd2vKW0BYou/kzsA0JP0lGjrxyeT/zuliv/65QJpM
sV3l2Ta8+aVUTFotYe2N24I8WHPs0nCi/sbuQo4P7SJJyEWt26LZFqgUTaKLgrCixTH4D0SeiKoU
DAYtEq5ymZPKXAkoz5+lsbX0faHsfUFYVFcD4r6SkY3dUCUUqxMDitDInbAXL91syUEwHdvpDGQ2
XviTEiSjLnqNCu2uFxEhO6y23hsiQadmg2GIt5hvk7tMfLv4q0CZJ7erGNkba3rsXBI7GIxlAf3s
FpXo6MiMIJDgfPT4ZxudXQnHVcnx30dhpAqLmIvm3mLHA6oLcsmHCRlu1YE9xrBsuomugGHR5Qlg
RJBFZNIF2UqiCbPSpIt6cCy1Gqyqic6iXuR3F8/1D8qotfVOrVnnCOSx6j2Xy7/TWHQetMWANYLP
MZyS6hZqlk1OEJF/9GhFnXNPvfLbBkb/+fDhQPcVx931euz1DdAGMLtZJ1braSa6UFs38tTtpXii
1XCrUhDNDvDR+dM9oaw/6+U2Ug9a1qlU5qfJXbEnc0gXHQF//SOKYGQvLZSNPnkwO2ffa+TOHk5+
F66nH+659B3sDHPF7bLGAM1OtCMiWXLjcY1PCWzGGJY9895atFFYhiY4W1N/PJeWxvakje9zONaq
BghlGwDxdGMTAiDVSJaIylvzLbLxNd+rhUOTlakNsd9NqhlqpYhBWBfichGTrkxNx3MSR841L7Be
38WnQxys5ZZ5wVEkhrRkX+YRBrgumnLzCNpNZBklOh+e8UUjDPC6k0IKJlGF24V1EJlwIBWcHVlt
gH7gfaZpTJD+qsn3ai65509mqLsMSqGn/nDtJDiy21xBw0bEeEdR4xsrm0sVPRKC/bFXeYVVY1qK
2JSsIRBM2Uomj79E/WM8SbvQHOSoae6/+LBwiqIpQXpTTufl+JFZHa3bf/i3UGuVx8N3Dw7+L5pa
OJ/RmvVvEImMOoSG81z3ikD/kwN/n0cNhDTeYlPMaQI2PR2xFXNb8+295rUcyTHrKJC5wFf/EZsk
PIjKA7dB4bqGQmNrT8iN2KNMo/xWOVFq3WM50vzEQ0vy88a9pldYpTu44Ia0TtIpD3nmtjvR20xa
jLh+3uboIwxUvGm2a62627/A9lh93ukT0o1Thed3avBS9sFHUVO0nap7t3dEs5xv1ijVFgrUxPgU
GxoUF3fPDlj+2/13TvHs0KvAsg5dbdswMOj4ObEGBK3sOiGP37iHQsWq0BnL8OeaDK9uFntQuima
G5vptbDm1oxHLFcbtRNInCokS3WUkX7jPvfCubDzma2puuJWcn6QglgSBayb+dvfdW/op77B5kjK
ChHLga5NAZ+IjJWRfnAD+3624288lhe29fwyM54joXSgtGxZ/64uaf0QdLfZ3BFdxKWL63zjUm3E
uS3E35Bdoq/rtxvmwMSxDW6MmAibPkD6ulXbXbDemK6kflOuoqznexeqM+TJAfjprtKKycx2/m6b
C/r6vcxCVahHg5UExeihgq8kxoaB+s3qwkVenpJbMv/ZELzVsdR9OnXGTZC4y+BT7iDcyD1b2oW7
OwMMqjhMN4qvC+Y3SUpwNenfR9x0o/SGOVyFGHO9OBzjkOOf+dZ5VtNYHpFhDomDtFxNUNQaOKxm
W2ERpknsWqVcgJpav5itgeaTIGPJNAbUKqB5OP+tdn6zhWdCEWrDabiz2DsMfy8n4dzCvHyiSo27
wfdVjtLhhVjAyfSryBVDzmS2Y86P4tqUp3CNXK0BArBUvcGTJ/qaHvAK6i9LhbUZF1REcgbxEnEA
aoxMCDdpm4gfN3Afctw1DKejoMsN/2LmAGKBaj9OK09KP2stTqM8rQlvExFNTnyfbhjiG5WC0cGC
iOU+nEHii4QOfuTBta4uKaqav3gwNHirrIKZRCCqeIgPGV9jwVvnZumWsxqKkwC0oJ9F9+fB5x96
86ho2MZj48v1ETTg/RtmDNGk/sQelKq41QG94F4GBgwVvcr+IfZmFUVFWSeNSatzkYFUeH5Xt8+R
rv+XIigz7yFpYPjlfz5lApuyxo5tbii8hGzj+CKAplKFy2VUbzM3WGAYbLNcwWpbi6oQWl8y19yD
/N0dCDv2phbFIYz9pzy3GQ0rdWefWwQlnzagFD7N0mZJYM9A6uOSzkBPAsAur+Y5nM8k3+asLSzq
6UVy/2Kf001/RSGISEXSw6Nsbr+bJE4u/jrbcB6I3b5hHyXZZMOVaPLSmrGGxZNOHYtvb9f7U8/b
+y2iBAuGqDiskvQhncVwQe8kSS/oGYOddScJCxsUJkKlVbJMq3jHlIhDZ7tGcD6W5UBzg4vgMHa9
6M0AJWpt5ssqHbASYFMwWiwRb+aW2SEqjCMU3Oht7B5//8jJZ+R55XwqD25wv0ZopIjOGFi4R/FR
MpGZEDoD2uuaPTiTTLZhLWfwS4JhimpPU64exIw4Eyw/pbQf67eTXd0Ne661SI9fabOaRSOH3ort
Cln72pChNhvvC48d23QycLRaobyHDogWQdLCmVmhRDsTekO1h37eSg0tonQMvjSAcVdaet2vUUfU
J/QW2hVm+cYblM++UdbtfPmP/TQs6+vzChao9n5mX6wzp12gzVIQxmX6EuzZRfOHm6qSRlcxfkHB
QaHpzJonnItX0Xa12pH1tHLkN/owEY1wpv6WdcXKPkXL59nyJe36QLIvJpEr6/aRvbDRmK4Rc3dr
iJqPOvzF3ZuVySHddqOKSNzm8IlV9fV9ekaRa+XvQJUvXIlZMFJ3d49HzdXcMXble638MFcyt5SB
ljcmipTZbe5UC8wfQcf0gmWkNWmZl1IsVTlvI2frM7LPl3uVaGE51OYRGK5nXw+NwSTrPvwYBCkn
kNkIBC/l7TGiatPjBq7aaB3powjuaWbiMA2pDK1c55t+Zf1JNqT3sSQMjT2DZWo4pPcSVwKCL79i
z08T4/YVsW43Iv58T9kx7+j6NUBDnbI6PJaL2xtKy1cDz8GUAZuT56CVw6ETHE+Tui6JZUqT7eYz
afGIBmQuwf0Z2SMLxwxDDMTSrQg4MoiTGSO3a0thRuflzXzA0LGmAFw3dO4VXHukVnqAsM2MFGz6
fMB2/WZu2gmY3MlFxbbwrmwYzEgOaJbHbM1jrzojVb7+jziGAhpPKEYPkTsgH+M6kJw7A8AYRPwv
m0QHMJ+BidYWbFF1kuMcfY+K0+JHdjnGVToj5rHudpe+yMR0pP3IQhV3aaCqMSVrZVPA15CJWSLt
rN7iSc1fivf+bwq0PB+h20is5K3rqZsUo10j6u29e55MduKq96zD10fOehBWSFUJT5M+6N+CfH+k
WqDK299wotdGpkp6stOJi50FtOnFlC2iQe5RgQccJywHah7dvO2MOkc1eQleGBvUBdYh4GZU+tV4
qPHzSuFbwn/MOeAziu8ynfOEXP/h5p2Key4mq0lbxxE9ngOd1CaRaQFAyfKq39o/NNxeOoqTIWMg
OZ6dHKUUVvR+mITbfAefV+SC6Zd3ecqxzUjDgtOAjUBAo1yUmrKfXMikJZzFsEo8AkuCA3ehGEds
2la0QCoJoTvBdU51+vKqiLnoIqo+77a8EgT6Uq0EFBpnhH9XGmOehgHLEVSJHUtRZdhAR1FZQMXh
KQrQmJPhUp3hmTA/Hj3kYJj6QF33PV/D2qap1CEThPYyrkkhNOfiOPns91yGyO11aKrwHb8f6H6f
Uz9TSNT5dt7XuBMLr2JrDq5hZrS/BFETHTUs0ekPZuGcyZ4m6HNb548TtEUqRJ8GAPWgJXz6Rdo9
nQR+8frPcVto3E9DoJSqKCq0zQ21Qroo1cNRqGfhI2WQ4LIBR4FP5AuAGOzHqAHmPpew/N+53Wyw
+NC75G3sJfX+0nYzoV2AvwHwwVhSbxMxgAcXrrynm7omKaBgpeuZBL+Af5uBxe+PqvhYJk2Myney
V8Xb/xwcaCBNM6tHnjomudLdhRh2YFMgtjrqm/+BY8SCkuvdGhdeUJ+uKFXqHk+mNuPLMB6stGwv
65SFjgPazRNu/Udf9LIx/NzatskSWglRDg/dHV/qDlJoBZP30cqbYPtVpFYYZvNAZLlU0avUlJFj
Rvn61j8HdZ1cv7chl+kP8SjT/ogCuAIVcSGhf6y/NDBH3LCtfwju+2ruUK8cC5cW2MdviKnGi93v
pSuJnh2Vd4gQ8MNiEulACvr4h0t9oLQgui3bkug3Dcgid+Fv+kYDq3R9XwMu1ChSzOAuU45DcI/k
IIIi3lmpUjDDzzsQFIyEAnch9UnRhQJ2Gc3hMy1wtzvA9e+UGrjbgb7XEhhs2FQwjxfjpbtdXHV+
qvbQ1rfXqiq8af9p+layrm/3zaU8ph5V3hQ9h6KU6pcNDdaNHONR4o5tCcPFLKm+nkpQQy3s7wD8
oDNpGwoaFmkVZtwbuuFVI8dTZ20sOlJJhrZyk5eDpZwIBy6uT0St7EF7aRWPRln3jyxi+VdVlHaS
tmj6oDHSnMK64k4NE+6Su+THqR46ud82O+QP8l0DFnUkLGSsxWkPUPTKP/1ziQotuDE2KY2X94nk
8HtkAPvbuc2YIbr/lFj+K5SMfDw8ZyePShAu6Trnx3VDewAjMMUNmZf1LfI7CZgQYTiciTr+Scw0
8cNDKkjtL/zUy1Ui5XjoCnQ7sPpnHgtbAseFPsuFN3h32fLK4rD4ZtZIHCAizwlhwuAREDj/8Nif
+J6JW/3u9No348N3yAnwX3czXBx/7Sq+0/8tc+0jryfWc0cLIa2SlS19Wq7bYcJ87xfEUunl2a4c
8xhgpmYebqror6eGFc1XHG3ftcmDLRbQSHjl41hMJ4e94ftvLh8/jsH1u6S0bK6sxpOS95qyAsjo
b8zVlvkbAKgtaN0s12iYz+2Hz6PL+taL5FYgC39Vpivb9mEhS7bkiYrgVXi0YNgwUiQ15ill4SLx
WTUbStrJi+AbE3fEZBwrbyYtiE8xpaFvlJ5DHl3mj0L86UBHBl1r1KvBWZ6/kTTtUlWS1aPH/2qw
DvJij5ZySQYmw1RZT9xvpz/u73C0TFM6p4gMNcdRAxyC2vyD11ePOh5CoHpF8bHSC0mZZ2oXJR/f
4eFHZmzfKjiq9okxwLu0U0OxIScKqt+aAM+9v9L8Wh2N7kDu8Qlb7HkWt3nD98TnDo+1F+86qIsg
HQ/8o+KIl6YZOYzc5EKdiCBR5AnyDUBsJJfHl1rdLrXrK/7tIkRR18TRLFQUC0FixyKZQspvmmgK
mdhAhoX32kPxMRzn/aJEmf/9C4uxPUZklaAduZR6fvv+X+aFY1gjrokRNDZw8FccQ4lqqMJw2T9Q
u+w/0FoODaXeScMy6v68sdYAFnbIe4hOGwxtWNcT6iJ2xoiHo8vb3/fuWfqE3MMpiysKLLB3QOaY
qTGVH+QoxOKjFsM92seXr0RYYaRDF3as41tfDJ7Uyk3r82oV8zXQY7udA7NSqb2G3+G2Nd0xJzzN
LyaQQGkhhuMUdKYDW5mLyOV8DZ5N4s3ZCRv5u6nQjKeDqQWwmhaxMRfBdbzZIObxxGn5Ts+iFubq
vFBZiE+8ytr18wYxNfIw8d/gqaYLn3fTdM7RHUcG47q4In5Bel7UlluU3mRN8fnuYDO7GgMmyBIW
h8AWfbid3/0LNWpgfSfdUMdqwH1xaxuVwNBsUUO157GoTx8Jd0HxyYowlS4TNJvdg9YLLIGVA0BD
iXmwyvl2q8eUhfh0xYU5A0jzPXZLVybqFRrELQZgZbaWVgWc5NhscYU3THcnV0XhP6BpWxcfXaKL
jnQ0OX1tT5cxb86AmNYfveASzYokjoiYOEc7qW0Gq9vg0/kCGy1l/A0cjgLVYG7O7NtCVaqkBL0x
YqxVmH70qUrN5q6G/0zBpb51yqsd3jdvhb1gYJutSQbE3TubzRoXvkJ52eK+OZETsKLngf27DRJ0
YDgz0zt1ad9XD8Z742Xsk6RzfL09I+6KpNh7sRf56l4Jp9ZOQBXV/oSs7L2YDKpzZcbRsXX7Im22
yd3uf6gSW3PDiDy205NWawCNhCsLaIbeGM2N4Z+JniB0N1u5VzWRzQ0udckuTG/2o/CsCpAq5Vcm
dRx8YboiWvkQn/0lbR9nautrPyHveFeMQHaxuH9OXsDtzQiXkKqxKtj7gVZz9RiptEEUCr2NZc6o
VH6xNee+mouKd2XBNfLaOWOHSLxJ/+JM00FVjbZNv2l6AVeh1KMRkOdQZW5IWRB/3pxY9Mk6eQqy
CevYdUOZlFm2SMi7jCpjts5T1zXzL7Lgqx50ypsAOmvhzvhDbEfIn2kzwHb1TIA/S2Df0j7yn2L1
X/uiOs/XGMVY+Mf3rDCs/UhV9JodRE303A0fEKNgqziurMy+02t9sGlwzOX8gt4HGkUoYh9dgitf
WVDa1XrUslm+4OK6t7GsZJWh8I0Kx9QV5pWasFT/7Wd40pNBVtJarmB7dG7q1bW0tubRe3xre6XC
3Z3dk3lv2+b1n/6eCvMNE64ktS3DR0ttYPv8r3r1UVqarrjwFh7o5/pP2U/Okgno7DrUYyyFnHZF
EEzu8ctd+rWrYSv3boY/KvAA5YecPpRDVvmqOkLAEM3W90cWzQXDuJ1z4vHNW5UyzI8bqxHqGuEo
MpyMclcbHctUxpkGCjRfhepUFGVxGsbq8T+r19UBTvxIsLMOrUTcWd1d9VB6FzDUXXocMODgE3gf
Jq9/EbiPKnLtJuOOXfjZ/yPKC4GmrHYVeOSMD+r8MyTLYbdTzZchsomUo83F0nDelRVeFLgrkDll
FjjXVxNDxROjagz9pZe+aC4E5U8wgUVs46fvRbO9o9mXUhjjTFsnR5+uHYjaKc2Sxwq4fwhObr4K
Wi0/vNiA1+UmAqCLCFnR5shvLiptVeTnUYhoDKA/fvm8U/U9vF/4YqbC8oca60ovo+E6k647wxs8
98loR5JAtmdeKmFhcWAY/Pz2JHZlsbN9S1qyZmd0IrPFoeOc4EDVzW1yziDNTRUUqdCYM4+jLBqS
evsNudTfcragaCVjCeBSqEvAHyLHF/tcrttG1RqzVuFCUgcU9WsEyBs63tCXOVU1jqytaXpc/Tzm
T1pu3EwGhIIQd7mf8mPx/yPt7/6PYQdFLRwsB+63qMtWgk9XAB5cAHC3iK8qFqLi9I6nJXEtFOo2
St4uGGLt7vGUgqwlE9qcdteGYt4KrmA+KKT9pq4N1J/VrrxpXgCUwTIVeUCI9DyZJJNbghYPoaVy
TN+Zw82oyZ0dD2/zbDj3GyL2UeSL1pL1g10SnP0Bm3hUHDl09f9FsCt7vBq/ec7Lc+4oLyOUH80z
SE3tciko6CWVElwj2ddJk68WJPmnJ15hqMBRDMSPh35PFtrs15oJZq6gLVCBw+dXPeI9af7vFLEm
Ifpe/nKXVhqEz5Mg0mqcw4qGj8gyqzSUOqyKxmLGKTJ0mV5gEA1bHNTvmPBS7okOl37CFeRW3rPP
+zS3qHppTyuNWVux/trE7L2y1hvVNfckksZwcNi5RaPYkT5dajKLK91E18Aj5LQmM3iSPEaqL3mh
YB19ADp6af7lg1NbT7HLD0JJhGopsomCJbUdrbENDqORftzTrU0yv8Kx8v6KyHueMd9gVK1quUSU
gEQQm2N6mGlwmgfNApZnQMo9jBPC1lVvTU5l/XqNG2bDSAn+mHEfS40jriprVmzfJ14ZGNGmCooy
WV16pTuFZndEsvTRlDbbxJ46asXoO5mpg+K0ztwlnkgt5DjKV5fmkz9AoxFV1+dtmnCKpiexHGH5
sMWfbhtU8/7P3mZxXGBYIQ6RPrGGVWNjbn/uzVGWhCs76kagAnXOFbCpXMU5KLZBqgwcPTuTZfiL
Q6j98cEeluaF1hOEhrQYnbmD5Os8sQnuWlTtnTWgNr5RGLD50mleAtTapjjqGf+WZE4ZMS9ttzx2
x2A2g5Tin9MSi6wk44siLawUTf/e6RLVGSU/uRt4aPZT3rwq04gGHQuvdgc/Jk7Bn7MB0PCgV26q
bwPiuQ72WVfM+oC7OjELT907pwDAyBVk57C3xuJXEaQewKf3XttDin55W5iUjVs9pOj99zDwf7mn
zXQNYemvF78WT64OdNpeJrNdg18BLHSwBjL6QwY0z8QTYtTiMXlBm7rqqwAVmv5glKI6fpmX5LLx
NhbI14vrgEv+KS9T/JWtJq2hEFW9xmfpOcVHYbE2eGBJFRs2bJZsEUklHTEvosedFNAPcoGG2F92
DSvJaEhbKYn00m4HTKW4yivevAUlIbaSYSdCa+rB6zIcO7EVW6c655eAtH/j8KNUfwi7PJwK0FdT
UizbPjr6U9MGm61N8+49Q+2Ww0/GkWjmwSHCUe2ytpqaHraNsMKDg2bBxdl7uJ6g0xIXJF5w0PvC
rs5ZvWj65UWsx9eyyeYDyHskM4xoCt2Wy6MK7EaHahwsqgDhagQv3be1j8aSmZEvXM5kZM7bPvD9
JFoySDXx7scmd89aPbCkYs5uy0Mwt981tPUXEXPH4AbFSJgcoKMtXAuvW1TnUIMP4dR/E8eU46Ir
U8Snyt5fJqyXUmNA6wEJPAml9ZZ4lsF3wnRjRlR7HmFpzWwAim9b+BO8bUs7vcpgwo+nvaRxmeVe
OgHniavKfnBR+p4lR2GnZ4Q3tZr+aOiAqGuEcrFu3r8UzOISHn4miCZgwPAD17sr6fm8wKyno+Sa
78WOKMoPC/ONJmPeK7VhSLwu7kksDa6DBUQQo+iyLyF0iNtLx+MI7n4qW3O1KgUyWbz8tpUwUZeI
HiQr60TTKju4ndOhP8q4+tm3OaYhXN0Ca3mgz6cUaL6bNimiQV9rv3WRS6IUBWh80G59MfIO4S9r
OwYc87hc8/SRvzNPQR+p3TkT6PVgg1eKmUhmXr9hwQQgK7iRAc/1Ll5v/4h7CyouZem5cyLdPo+m
bIKmJfVzJeAST7gS8pgYmo4VOQrguCZh29YsuncowTsPjE/XeMVTUf8bUkyc6R4MnI4tRfU+hqo1
bccYbOjQY2GTPTw3st9iaOTGEQKR39MKDZQQpnJf/YmzUtil3yKJVFUP5kE7ZpM3/KvGZFroo11E
zyTLp2FsSsmm1Oz29d7CgjwiJLvXFl3i7uImaft2JW92vBE1flI5xjgzKd1sEy63bq3juXahUEP/
LxH1TxSlWbh18aVtMG+5xvpGq3clzVVdNB0ePhO3+pppK7wd/+UFMbmoaxVwGALiZbiJE6Ra6BwA
FqyGvqPXa0mTJ4B+2NaZCnPin5fah57WmP3R1RmVJnGWHD3NCaJgnvVZrqjQOPSeG0ANY7nLGFpC
//bCha665YiZ4cv6wDz/tq9IfJ4o2E1nWwDobEqU+5Q6NWjUSo9ytz4ZWNZPHHanT42tGpm4LaKI
yTMh5CKruUfs1/F4h3mdv5dg+bjpZ8cHpqDcNFmwq0+CT+SeEffAB/F0SJIChP9gXMhg1I2AMqxJ
Z0yek+0PtBWDXKeMLaRxvlbIdfaxt/6LcDCtLZn3aoPdobQGd/dlBGqFqXXKSZcOl9SDGP1z44Vg
BPeJrkS3knH/LkLeFpU4FPFfz0v+5EKrjFRb14zYlyN9fhUShMZHT+RLqrPDlxjs+BIYRPhH6kA3
LDviptR4yOrIMplHiXCuyK3Jg98AyUzQL0uxc6TjsvDaQnSQYiJZI3Toj6Rau7cvd1zD8MLGwbl+
HAnfIBXCji4D5UxOmmlIepey1P5k+8LCQGfLIr3I29fLOAA7H21D2n+0K8l47ynH6DFnSUmAbr0o
bJDHXl4WFtBXHmM6umTxlcUOHHmgwOLUtToqPuvNZQiOB7uMlYvTe2ny8Txqf/SIvBX2mAp0F4b9
i1FIXeqqIeUaQKO+3mFETHKDiCeJDUSsizDXlw3A/FKJb7JTbgomfrQgLFP9LhngeI+Q+GnJ+zPO
4jEL57uuRUYkpFdhIOMtG4SXyG/yJzxF+723Ng5x6OAIamvyEUD1mQQlG/zGwHutOoFv30OByV1N
GF654RMwOCIjIJ4iW3jdxV5XfdMJiaTGluch4pRxc+99lahjzGuZy19RjhlOskowIBJ2QvaVeuko
qNCh7ogSB5qRGJRQzz0BRkopBcQqU7y7jNHZatXxUWOlL3WzJNxXHDgDsUf+bIlnPjztKm7pJ28R
xl22/ATkmfn36oMJRmPN9zyVct0dlLKuhjA9O0nK6gO2yF6eBqoNOxMzCeU/ssBkNADexYyJZG/y
MvMRh26G92DohXaDLi7Y9RKbt4jAFANI3JAcZ4vxRl5jy3lPZ70OJoNQSdQYDpW519JUgqPzf/KB
rDsazYLE2eSvs0JLajgzYs4W0vHg+h3fquyz6MEbwaRPYyTGWZk8OohW66OcIbz7qWM3UNeP35zY
msT5P4QTOvYBiYdvOe/7Lm9y7tBbU3nlUJLT4q8/jH6S8OYd7Bm/qoGYpg84PpQgcjMP/u8/zOQl
uPZPqWvq7P7EFKM2XrhbBbgM7feC7VReOlg2Qh8jhODSv/4Ul2L8oJAeRIQ23b3KJAzu+wa/9dNe
48hTH6CE0IHQJAnzPFYOrS6vBCEBJE5BB/ywFRbB5RWaKLFu4ZtPkCGJL8F3RsqI9Z7gaG2yHnvK
GKGvCQx0uuz8Kh3k/cpozpYMxayuKEz5OW7yGio2xHhVyRria1ATcpLOHu5fNTm6ELDPbtTf9EYI
SIbZfMj/KZCqnRZVcrMZSZcwWSyic64nqLuX72BfiAF4cojZLaOLeikWxq9CEh2OMz8qdYJzFObi
iL7pv3DxtPm9goFFQxs3g7JGZDeX9pqe59UZgRM6VpUDIv8bWO6y1XmWtoPDsL7xVKBUaBQWU7+D
ltv1jrZfe6zzEbAxUcwEqgMrpWRVYKSa6Jb8e771YWK2t1nxXWklEYk8hnlFexANOpswR/LJZZga
JSXZt78W9HZELO/mtRR8GWk+oXXlCEKgW0DqlKSdp29MOtiRuzmDiWhHTzwmhO12fCzqAvukG8Oa
niiLoJkyfecjkpeFcK5QHpB9X2zgsPHnzuVIR0EaHs0A9JoAgq5c5Mr207CBSW0RVLIbk01SXlqS
NAQUchZeOnO1k4SFK+XfQgzgsCd7PSRuU59PB9S0Nd1t/59hzH/aLInsV90otEK0c/pmIuSzOihF
gcLNQzmWzpJSappd74wSl/fjMSUDirsJBoaRa+zNDI0ZvqZ0/pRclrqALsX9QtQm8JA2Ppa/oeR6
UXrdySiPW1uQGNW3GtNdb3sQTiii7RZfvJQgJgAnWgRnKBQLHAUdXaard8tb/WCFXPkr7dkNeSAr
H0R+Kz1csVX0nLxZHmDY1DAIIyHQtH1YIF0EL7DgJqoqG/cE1zKwriwfHNm8HvWW0cpc9zLgrJFB
E8ovKH/LpQO0Qor900xf4F3mgIB++EfNGZ+yEt8a5LDMv32bvrdzz279yjSd6SylJT0Tt3GKfuhH
G09QRwWK7d9p4prvFEG3AetQdWSYcB2LQfdU2gi2r0YgGPZurm8dPBNPGxi8wbLifObkI8CNF+a9
1Q7FnQsXRwjbJzvhXbyZu2eUzHX7FOYNja+3dZCxISQDQ/ojhfdFAkF+tnc6/0ZHGxZNz65mAd1w
GP6TFol7oAGfQlmn6Gy5XOXGEyzv3hOTaPUC5CG54H/S6cT8+XsuZuoEDT+sKCzzWbFHXdmwRX+8
8XYgDqrMIXVdBSO7woaVIzjfiV5U10+Dgb0om3v+p+m37tJ/4WFJP/tYOZv2ysnipBXnuFYuLLPp
WonF4Mp4LKpj55wgtX+os9H42yyvoBFzrW8/RhifiwwvbYUu5G8bkfgUKLEAyxmCyWljyUrOeWtr
VH63npRmWV6N37v7lYDOaNh+akA6yW5aJJynfmrfo5GB5TbhJZ99MhRFD1skx2xY/9vJGvS+SdtX
orhW5Epv3xAIO+Mv5pkkEWXQVF/Ox2xJKyfIABWBoChAYettHQuv+UhMLgIlVOds4UWAtselTKnd
WNr2gy8YC1tOo1mRI1i23Y6J2RD9U1Lmj3n5elk2/hSqm+jxgZ5Rd/80GTk1rr3JUo+LWpzOpZd+
vBX7xHoMhul2hl40KlRTWD4A14DiLfKftjycgFgBYPLwraVNN9UVX3pGBp9H44t41qPfP1mTzBn3
+J7/0mY1UAtAukwNrKL4b/LDy7rXHLhHQHmHhzvxTYhNLF2E7TNdlhmeKiWNgw6PHNxlscfs+d6c
Bz2B/NLrdWYXPSpOmC5YTZk/Lx66dPZIKAY5O0TDtV/2lZ3EbXGmCugLSHaR76m91AW8zQVIJ2Iu
Zsg+9fswfgeDcmDkCFANiWG+6Um4SbrsJqMBHnjfAegCxUmsfAQSRI2JT87J4MKgpFMe/+orIzLI
XxUEc1nvau7uvDbce6Xzf71SLgkdvumAErLSfBTGZ7isQ1v1t0ldVEV+rrgtHrFNKlSMvfch+AuX
5o2F2CoQWUmutxRQUmrLE5Wof4LhwNihopuwAgJbUd8IaDu2u6+MgD+uWCcMIT5qkyYXCHPNSlFi
IMK0UAkxpY6KpqssFHFICnmWTFsShbnTO35MFkUFRPw7S6qWnhSABtitgCLS4Nbfy5OTUHW62e6g
yff3Azj5m69bG9dMvu+sbrTy09pyiZn3f+adxActb6dMPA8hdr5UNzPebgHpWcF/fTLfWbCd3SPO
jLYy3L1JNIDx1STxoFn52otDQHwpe8C9gha/Lr2K6QF0h7JBud8md3QcDtrhqLUOAdAZJ9NWDpOk
tQ/ZelkI/ECmwKTYDtlsDPXgNip85gGZGo0QEA47qhrjpfZ4FgZ4Yo7rUe7nMrQIui9/dUetsBAQ
POQiGSs6sNs4Ep+TMa4Jri6V9i4UAUhNTzPwNGxOceO2t12hNuOojhxLH7++BeVzf/jwVKF44XeD
1fBZxUpxF7yfctGmvvr8ZUBXq7/4anT6RbSpev9/aMrn6bdpLm9AOTw/fWXmqViCVXdUCov8S8Pz
e17XWm7/ls6oxX9qZoSkPiAwJEHLX8FTpJH63ixXJh3L8xNvd+uL2nFD2Qjfu9atMdzJRZgtQNlf
zQqVT+X2G7UWYdENkRa3QUQp82uDlqmtNV95I8LBwesstF8x4Q3YgDJwQPiMbd/VF3rH1IOzITZ+
c2nNrVt13rlKyzfTCVFBXHxmGHWV83UqCmZ/pYOfl4pA7Het37Jx42dea1LYrKX3EJhyN2BdvNKK
2rbMHUqYN/Nw/UmlGFsrYIBVJKr8i2uOzElydJRBl3EZfwEp6cPOvpedYGImQ/xhuVBO2DgUJwFR
YL97ptPAXXpcnY/w+2Iw2zjRHQTY6cz/gHa7zd3KXVjpGdm++egrXhhdgZdiacgmdauPMriL9kmr
c9zmgIsX/wHIxvvxAd4fxLlxvcjsR8cYo5wIArRCcOiihg5vTYhGF/pnq92yvrr+PcUY756vyGsk
Ne25CCE+APQr4xKBK5UQXfOf8p3o4XCqbZ40/tWP/3uENp3ivB40jW00TitmlTVKu33zVpHlxRf7
QUhRdkP3In3PnBdx0EEsUFEVm/ta1j4/M1Pyr8LeOYcr6LoorCbuWJEF27YPBqGLPiooQGKNUA9I
IvZ5FkM87tKLOdeDhtEN4zsZXZSTHa6lVSbbjGGGkUSSCa+PppLc79aWyNnTlP+tGtRNwaYnHFuM
SGr9Qcho5thMLwYsclXE+8v0TuPZZfZaWrFMVxGiyYD3i2m2TUMumsCHmHBHOe00MsB3wrD7I7io
rJnN6Dc619Vg59Dv0mQ/a5+dhByG1jWkr8btXuflD+diyfVpjI64sIDgfDNnxhAnt3Y2hvbABPpX
xnmFCHGkCXIEOawFbEQ/K5KAHX7pn2E4MBCV5FLtpQp97VPmcKRspcLfqw93lgJ/0ZkMnOQawlk+
JYZ4k3XanMBfD8yRTbPD33oLa0ToOg3BMF9K+N/aSA09+d2N1XlTz5tiFWVlDCKP4uODvlhEzsSs
UpWHZwyEXw2RnQldQ/oMHbaS/kC/vYmPCyWatdVkZCXvfNXh7/dibKloy6fGoOGoFtk2xGWJdwDJ
7MYJ3CJMY4vWJAdSEmctr6DZA8m0cePFEVldOADyZ2xXeX/XJ0UIoNRBhYgDYGF+DJg6nYoo6WNM
XMvLz12Uinn7jcrGn1pMTIhPgL004VZsTINmHQhvmXCmfHY84VQfANHmoGA1NcZpermRqI8EtXka
4v/eCyMygZNBmcOsHIncOxkzXFDpIJTfhowh6aLbGMI8qqzEGM11bvEmge4EVgjfy7hSB/wlw4RN
ZCl7BNsAIgEqSPdwq/b8nU4PJen1AUVpnvvKwtPT2NvxQolzaFvJuItKgNdJleqp1rxgkmc+05zM
MOczx1P/cCVbJ+r38sBIKzRG+frXeREc8zTzVX3EJECX/FnUVetBuw3XUxXjPpfBX9XiididbIC1
m4Ul5+txbHSSqcPveWomH4ATV5XIbUZB2yIaIL+di5XvcWaAGm+GTXt0jrUUlekAJLqoU1R7ywga
1kqFe1pKR5O7AOkDc5mh7JJGzOXOrv1j2JIXTL5b7bdLu34UKj3Sz5u+wOgB1iY8dJr3wAGu2T1q
nD+Q+DdftVSrnwX+ENio+VM3aIt9TAgV5/gMQY+3k8mVz6XnMzpQ9szUW5md2GjaoF1o83n8WxYP
PdVnMwfJhM/KAEZdXLdD0iYzk3kDZojOAhytu1VuIG5zihbrxFB6bZpuImGoGD86/cTHryeBPTIA
Re4gNjhZk68psBIVim9uSJCxNkDFeu9Xe5XGscLqmUWXKSiU6NQEyqFx8erIcQotl5HG3wf61leN
5hQK5hMcYLSw30Hhlt0BdDUCBzxRSKOLggUgBMGnfvddktEqbSBT8Tj67lnftGECfl3hURe+rhq7
0Pxo22DZjqVbNkyofdUibx5x8fnOXoSJSRYMDGIn9+ydaPcJgt6kyUDAklz99pseObIjD3giekYn
1KdCQJArxAx/UGaYUhCGUd8v5OHaa3etDMuPX/2xkmdh9fkVasa39d+x9Z4h1hS3DeXvAzm/Q+5A
6uDJV2qvbQaHJmRtrKN8bgLgvhsrluGHjTr3wz6Wx3pOzG7/PvCwGHBat0YLun6n5pMhTWPYOP/j
j1HOBZRteSqPrrhuFn2stTe1AfvIlnYXMilPhalnycffdTnNsy3PgZUo38ayK7ymtRoFP12bza8h
9c/57L9RFcBj5WzqZWak/IXoPiIlLp3g4VDR6DP7gQVzJLznw9+bqgot5gk8ixAU/pjcXd3xT+Sl
Dj+xjBJUSq+3i25AS/soz6IojxKPUHpLNe/8Cy/6wtTRXKX5nxt5y7/FWGKHvntrajP1wj+M3HQi
PaOnYCgRvBObM1S5HONGjmpkDsSQ7TDZAZwwIIeyBIKpkEVCKilw30je8FHaT/uAbxP/pZfHmHkP
BXsJtV11V6JVGdEIzY5EheoIADbGdkweGNkYsDShofkf9ssy/BJTuXD0/d0Vcm9ETgvW4slblFhQ
zA8rbouF1C5BIrryBNgvSI3r4mpWrqAezuQliQeXy0jc86/fmlaTa/W5Ir3b5W5vS6PR/jvFeCOR
wsXxjQATNVdowEgJUQDwAZQjxmcHEmeDgGqalr0tUMnF4GRdWnYv9RW+qIj3mz7G2bb21BzzQVmC
8RQ/5DY+19YAYELQlZ7ZZN6Eb/Jfp4PyJZ6dOoGFnEo9zDMrfRA15e5fvy5CvPwtG1/mWslIBwfH
5eQVMqfVEDTSBESCHKlM0uIuJ9kE86ulwV5pIEI6HZVznmIcHjxk7HiEgrqb3QniCxEgUBH9F23Q
4YtRKqSsJIQBSCCUxRSWNSMIpbPHMgmwe0oPn/DwSf/YV2+yOwoWF2yJusDalGu8aNMzpqgnsq+y
30ApQQp5JNsrfAHDuzKtj3IWiQKrTRq4sYmKTnoh7Gwn6q2EPdshsrnbpirmOu47nxeNC1VmiSBP
NCDcoxzDpcACjBCGm8aeaXPm/9U3Mwc90fNeh6Zw/cegWYVrWiTUe8ACKS8EP8kkkcd7hWq9NVOQ
vEA7rzjnbgq4gbKtEjp7J/NErdfNyAnN6/5i0S1PYKKgD19nAHAYWAJesnN9TleFBoLNmRQdD9zB
czpyQ7qhYPDAKUaSXiiVzdGezCNfv6FD9rYZkpxpPsTmJvOCMvRAfGHDYWFUf8qEMW4i3a3Ri9eC
BUqUTJykg0tq2dnfF/VJBEo0jSEaXjmBcvoKZjcmwT0DviBQzW/djPEAfYe+Uxn90iyKDv3KpiXW
dMmCShC9APt1I9GT8vRNPU1wGr/4UB2NODg//ZLKnFJ9ZS2jAANtkPRx7TiY9uvLCwkY1rPXAlH5
sZhXeZBJE9KOkdxzrB1Ahe1DRW4CQssbiJccCUfs0sxIqbbvm7qH1S9SRaoh4b/CUR02A0euKW2S
gmfDA2rgamuBFDGLvBF/lhHtqJHpsX2Dq3iiHhar1uyLeSs3itneTdiPC35KjOmN3HK0pLyzkywc
M+Vo1w2LUkOFCNM2dy1evGbLdf3nWgokhbFyFnEN0erUw2tHoIL5fGPvAKVeUBlreOm7rCQ4k7fF
RFmD1soL6iDUJnYHzwpTkbqXVKQcoCO2SVgnK+5PdYwooxGkWhkscm52t9VR+3RIyjUKZ5x7xY3P
fwv3F2t65pA3OWZmuPBYvTeetI6iitJ23WZ0fV0QSrneo6ZfCDHet4he9t748v/FERgDHAR0pImz
tJ31681gqascA/+WMxLC4mAUjfPicHAFu3NxJMJxJNtbsuJB5B2HO1N+nMLGuox7GxHU5G0MRDi0
y0KBa4YAKMXACWyfatifBSqYSRNNxB7kXjNt+TRCPOjgne3aRuA4AGLBDrVXAoTDDRmJdtrPzCcn
d1iHdVrHs7noPN3NmOs72OFuUTG3kA5NauucTibR0q+kiJPNtIyUKi/roFW9k6M4mYVzEq1R8Bgy
g7ldKS0rKecf92ANSysSmhZuW5AY4a1IMiP9qjx0pAPaSkYJ8AD5msWCxK8YoBKER5+l4tN2MQP+
3PX1OZaKl0BS+QKxh5nfWyPAweSmLS/Hfdh/GTtEW17V3v5qOo4iCshoOdX6IVTI45530ZvtKOFp
j6XmTexxqGaFc1Yg++S4GSIW966Rx+8qhVsg8AlteJgU6oFNfNMSHxOk3vY7Ohimzj17Xt6iLLGt
I4InJpl48wcilF6Ps/a/sWlEBFz/ZrlUBGysEPsdB8dltJggNOjpMlGyRJ1YnP1Q/kUMIGdPpn0C
gAF/x0kf6bpmHOeuelcMXXqhX7ML3U4UYxR6YEYzpHVSs2PrwohG1dQCWp7wKm+KYqmFfeVArp3K
sLzgPD0dpCElgQcRwxzUssXjHMEqrwQpNTAiKurzSQple+cSDT/B+W7c5ReUMTXBlLYLpW8Dqt1l
PJ4jUsCofLksU+qBU2lIaIiazYq9k5HlQpBXZvZWrOnl4St1xLc3cBP/t0PYjBdr+J8MkAY12dBd
+JB8LuWTXBrdtSM/BJAs/dqkEkst315+ojsVlOQHihvfiXsiJmc7/dwHf/2q7HDUpeq+yZnnvZ8S
y2pid8mEifT+wVzs5EXfvI4HGgsT8sy4twp0NkmcLJ48CO4/dFnL0juJRfCNeOrTTjHT+859oQr8
nGRZ7wye7CwVQ3U/6ai9NkYCjWqiekG9OnL8s8etoQVY4pvlENAxPaJi+eDbm29KU7nK7buRJ9HT
yTi4KBZxTK4sO0bOWKrCnPwjrgY+gXcs1QXnxqn7VMaOmWsxfDjvj/rFScJo/XrG0RZcNNUFwcTZ
S4aEZ7ktwCOtE/gfKKynp5AXQCCRlS8qXnXdiderCZM0dUEVItuUwOemKDQDjzqwPPSni5IE4fEw
jReESBRdeToFmwB6Q94WfP8eQk5H2TH3koJD12u2GKunh6jY6V811n+22Q3v/EMDl4OsBTIy3JN0
q88MkgP5a0o953axWjFvQxlpFA2GF0zApd3xQnNSKufBM/YnSFkmk0zpqEoUSriNpG1vGePEdw8w
XpJxo6yFAwfHIbX69VIrF7PdpuTPKtT/YSTNwg3tC8Aq4iyvhwKGFRsSqSt2zqkQNl9KDMT5ln+s
oT4CSCOdq3V0nICZp7VxwvkYyXDeMpEdeP61RXRjoTQAh0nBIA5Da6yk+/0co/HsGpssl28Rsr23
isQsaKmojKBP5Jm0Gla1hfGglzsklenWcuVHSmiyQtrw7LjNgKSDlWl6VfdBABGkj06r9GoVSKAA
8N7VuHJUxE840ambRM48/ayslNYrp+DEkv1a9CD8Mtx0BuJcf9rI5OMvd+2Em9rv+9bPWKDHZJIK
zmMSQgufLLSgcgjeEDMTgYjpoy2w4yJJeqEuyHFM4gFGP0Vo+9efuNimb85V6E9ccUAdZWNtiRpy
WPebqOUe3Nl4HQex0mxhX436e1+LSfJ+mJCIvZLHOD6D9PBZL1beSmZLHjVoEkVej0sNZha4QWJx
GFEZT+QqUCBlsf685G6PfeAJgRzMdiNrihlWvyD+Fp+aKN+isomdh5Msw3KzwENmZpQh00MZ9h+/
UFCwA/4knCwieg4wYjqehdGW7Qb6ouq2ur1KYzOX/JwIH1U4L2/LSUfiWNnu7xdyTAXwI/AAt/Mp
qmAfCBnyyrzVKYjj2arrVaJT6cu2mfrMH2r///95No15Ot4CZ7805g3rw8OTp/gzON10kAkwX3Aq
4LFeTinJsweu5S3YL/eVS2v8A2/RuRk2K0u9FCJ0GaqKSWa5naar6+Htm9dlVYi6dKs8ACbHx6Eg
teDjLWajHoKB2e8SNBi6msG2QBLDD9XhI+C4s8AwtymxjGgksxIYr4s6xSjc2SmrsK+/5WSY1ZiF
ocM75XLz7lHQxbIGzgN7IxOhbTv2kH4sN1TUQqgwqUsDqKqhJFZ2tZx2tB4/2LXjSFOHOMDGsOZW
ajG8pNg9xfZV3hcAPTt4/aMbGX7V6CMHbKW5pViw8kopzsLFKoDpy7tsXYoZN5pjo/al3tZR34Oe
jUmkrGdiWxTupWiI/emRLJFZCF3JRm+GBmqlsZIqyH8IDXBMzAc65PGd9Fe/mAtdWDvGJiE5w49p
2bMLHz+Xg14UivnzJQV0GBJTaNehckEHEj2lKP8+x3gjZG/k1aWU3YDAlhqBdEN32cdCFAbDmg/5
KgKDEwPk4BkhGBKjPDPo1fdEdGgPF5sJQZX2sb1Mq+9tJ3NvHnLUYGsYzMLUJp4Y2WXTpIkdDNWt
3U3dVDgqoGjZ12xdWng4f2kn9hae+CZSwIjAE5YkSoAYlDFlfX/nAiq2GwDjVp5hKm3CJhVxmGt/
28ym1bu0nuIZZj4izCWunuZMJK//JQTmerAnRaUINPxBOWm2maIbd9B48AepgyH/wwdF/izbAibo
CaW50Fvg5O2zaedEP4EB6DZYwFal0OYvtZRcsMBOxpVdLFUiBI/yNgn0HONq9QgZFKqoQG0vhYrU
/B/64S5fX7ecMKyPcwUAk2SiRRTY6MX4l8MQZdNy9cgmFq+5sdZ13tkFMfrd8ERDZBG0NiTVjDbt
h8IromMXHnW+xyjOoHQ08K5gjcoGzYxPQP130fk38ghsGKGsX4hrFPdO2xZH9hj5GbYQXa5M4OF0
KGxthHw2SIrMa/mnxp5pfYjwPSbOovWMhdzz4TAiSw3sp6qqEPo0B7WWwWmulZ0CiVjlXCl8XCS5
LmyI3uyUQSxmKo+KvNjP9Y3CzYnrKJbNJ/p2/rbUh1uZ6MiJxvNCI7mdls4bfmN6AVEsjxieKbRS
SK/HUFV7l6nUnbvIiy8Hszkhg3LvUoayqGx97c3/ZnbNpxKWxWD8o6DBR/R3FiI8QOFajvMvkjP9
o8amf8g56P6q/oV/Wx3vIvYF9tUBiQyPP6TcdW2vYNal8SYtksy6ZXU10GcCyEUroj607N2q01KT
jyLMf/JpYcebv+2UHrf1r5TwFqVLyJ6PGcXe2wkyCtYKTr4JUOiJQoolgF4hG5EcqhmaPQ+bwlzd
ArAiot/PrzEd2gpu5njBqxr9JgziIDFGsnngDo53KtWY7C6C8KYJXMZjzb5Mf0yAMtl/Tdc6RN1w
5KJX8lFrSxa+nf8LgWGDScTfoM20tG5Fs08/SpeLzL9ZYSPkbnhwpbBw+l7A2uznEj/c0SnHaChk
Ct/UjPpFiR4fHDelUt4OO9rlopYu3aR9FOAU+FRL2enbQhQxAvXp4TcT9LVnmeY72iGMnU9Jvijv
KopTCZBSOI29DbKuCU5KTa3s5r+VxngUGYN9FunwxCh/H6eb4uUEyjQrnY44TMyOhkXEjUMswL4p
siF+Fc4YsESYAkBKPj8wno7clNt5zRCFhAv9p4SFCRZSOudU8TujbezhgGqBTx1AbQF0ku9a4dvC
flLWSKkE7uaoiYsJMzp1s7hTDkue2PH10+78TIT87+9W+30J1LkMrX5KplXIRt2Ucyr34AdAOpGv
TKLpPeXA+JjpWALIWacbU8BdtCGLdIxaxFX+eSZuQlgDKo2J8xcG1IcXiosP95Ctgojz0yXPztoA
dc2w256fSavRMQOxhF0eTe7qvZlqKeM877vNWchBSIviaTEN9ik13Mp+22Gd2emkR1hxNLCCWkwS
bTkTy+EqKhCHRnN9yiIJfAs4u0pyK0AJT52aOvjuT4a6+tMQUZzkYqz3tIVRJJihTl6SBTdrsBwt
IVRd+RvZsDRPmjK1BmxffeAiAftkR+sYxitzqC5+GDIltkhjPO5gw9YVvDnT0xJVV3IqEWYya/kM
NRrKL5aG7MwcathVswRewjw4fpfIyXrp8UPDMYwhLd4ppGdM7VdQz293F9mCl9SezxltiK96irKD
1S71nQJdZeRas+5rW98bz3WwKDZPK/Ku3B3ypy2zvGhoCJcQgwfAoKcI+jssKp9kFZbg0Q8+O3+0
gzrIMY1Px35+n0IsD0jKAyaIMx0TlDW86vY9fG5tCU3iHbS93hBUePkyQtNap5OLqqTG/rKYhBv/
n813a5O3vflNYABVT3UZGtqkmA7PpsOsWK6a/+ph8Ly5cWAexwULY6zH7unD/kk83aPX7bd5D9S+
yGQzc9ygSg25qfqNpMJF/2cg9JIXbzWxPfCKAqz51pn4dwfJxNXaESIL6HIy9yfFHZwyJPENXJbE
X6ZvS6fGMtcxFHvSDMKQVxXSSHEUIGCxCbPRTYckyOebPGei6Iv3IhIdGKmEOLHoewAROLJ8+ce4
0Ae543O8JnOUH1TAPjSSvKhim7CnBOOgeTBkEi8ZuG8+8KIHMFT5oyvHQmnQby1oxO0IiHuNkK/m
LJo+S86nCl3a2rO2JRhzLdpSMjtQ8ZAG0Ed09sYkxKT/mvaaBg7SlgCmHVnlmnyIw73tuzP77L+5
KVuyJ3944Yqy9GH7s1Vh0wmi3niecSXuyD+ZKt3/4WufSco6oyOTwjZSdEk+BlcvVafsakA5uY22
HkIFNHmRuL2DlkBJR4jQFb2v8F4w6/HyuLoXo5dWHLIBb43Cbiw/KSlqI0+NKB/SpM4FWp1qUC2u
7pWNBSvz9ukpUSk7Zm4vww1fNyOqkx9Ju55pLSjoZidTEygqdZIbpplR3j6+ME6iTh//os4nUApr
G1YI2P6uRxM0t2U6HcsEIhZ+0SbWyYAnz6ePFWuAkY4YKcIr7JKIhmyoE8GJoRZZFNu4qL92ffm9
fxh2CgNOSt8+cbR0NhuvyS/CIS5xfx+2z5WuFB88FUl159Vdl/i6oH6/y4Jy6EH/YtrpOpmS6AqS
CGaZaXTXpoY27w6C3Ec4DU2CP8TrgBNd/Kgm9m5tgJs1o/PxcVYqgq0ZXZ7+IzP9yjaSJ6vdzG8C
vwkulwEkqxcWgZs+80t5o2VrCkaJLkc5TMv1Ac0gVIl33PaAEAU+meC82RZD/g43eJ8d4M7+t/6T
W/Nt8TcEQm+tZuoSUNwLvaxc5ddgQbWywYPqRpsXWb4diSlIjAJb0KKOS6eZ/w7RX9lDsqJdWjpE
ec4kXEd/ZZH5uP5jhsWPcMtgsSA14m+clNsJlYzhWKifV/X5SKT3HvTFG9XmFqrYhILcsfZfXMcn
X8cYvBjOaAK57hmD9XVgD/pmBgnozXbpBPOCGjnjrxoXhac7KmmXvTx153Jz6+YPOETBFhahuPel
ks+fB1opseZXJtLjjQCECMCXcHBVmkcBTa3l3qxbeo3Z3EBDoQR4YHjHmkv8LlqvOfS3P34O1IQb
m4xK1JGhE4BU6lQnWXHpnr/PaXg4+oRhw0LN2BfMNySotZoHkLvLeF1FA6a6MwQUCShvRnrxgZvu
XZjsHXEmjyBZ0b9NgIMd2u4odwdF+2L/tZpXZdhVx538zHmYgGsXWQv4bCrSqSAGeplTeq2PAoPn
ZPJj9x+QVLv5fXCo4QD1APUvHtOsnMkTyYfxbWoXtdnqziQMZiABxXIzUse6Y+eAGh6WpOQzezvM
W2VBAHPivKjj2cpNh5GRYD6Y4EiHMvkACZLx31Wp15vCuKVja90Kidz99UipcDN/gr4ixjTVCQQ+
N7+sE8ANmhdvVsa+qZle62m7Z0cfyTdtXBYxQ2x7ecGgNFdKM9RTFYA0uaqVAO+34i2cojPxTJPf
kXVoaPiCKnhU/sWwmBQaSXkl3bEOQFTar8C9/mD5sv3jnI/yVAld11zNX6M/vvnX8ihU5x7HW6Ot
YXeSOjAJEFs7rn9fjg3ZdqklVZrChwp1jiRthAROyjq+3Va7JDCqkJc74B4gJdm+8CUOsmveavKU
FURvYBsDPbq4my+Wy3Yywt+GLuIHD2I5TB/UJv4MaW41/eK3Bx6FOnAR4EnpT9LCpmQczHvGC1Tn
U5U/Ye7vXGAhlyDvVLlETVy5nWI+L3CLaWGM5PptvTF+gWbo2Q9R/fFHOlFAYSymIlu0+oATB3qE
ejRNhzsXY//qfCkrbalJaEChd14YpUPgd2l56vbvBX+3C6kOKEqr6BvRKurkXXBwxWDNcJf+8F0y
wKAfpoikLOsQPtZOz0snypz7gfOiPoOkWM7KSA0EwzDJsaQaVOupYttiiQL+ewkhJ4UTMrwmxsSj
9oVmajRxLWVK6EPxvm3r+hSDyDDJ6O5gupjXz0wR6+KTE8HdbJJ2jzmB/tSMcNOt4mGBij7PpunX
RkmkjjVY+hLZ5DzTDGHQn97XW/PNY+13SDgVS6r/37vedjWNoqv3Stli+Zvpx2wW9kW6z65vJbgP
RiaX6xqoYKk548B9MDOtKapLUyU3MhKnA1cw3k+sj0hQYCASWkqCznQUHRw9unzTQCdhFz4pjlaA
BRNhxtTLDtl03CS1FnAMy8NsAhe4gohGaghUKftK5lfWoBRm6AddSmLmJrvA77Caryh2fsQJ2GMp
lyxhRjKAm4/+WB6ZOgijBBpuvW9yMHVC21CKtxKUsNsoJvgK6yZKx6gmX9yxm0gVwtNFufv8aPWF
7OXZg9X49ru0TlvSfMdArVB5A/Km5DRl21OKgoTqGTTdcMAfSlazhgQU61nU0JxHXjQR58ED0fG5
BB08rLv4sWfNcLhF9sSjTDLkD/Dy8AB6K2Ky50iOJDanld8tJd2Sn9A8+KD9OU4pGEKEOjR55t49
ebqinl/xHg7ThLGtbelVcD7VeN1epCie9548Hz9+yu5l3jhoUu2Q2AXuRZxBLi0hArqucyVX0302
Ulx7+bg0++liQ7iYsXKm3hAT+99qXUPA2ur45HC8GsKAyajBFpOYsUaaXwjQ+a15HOx6y3u3ZjTp
dRVSwMIHOarEwWJVTVUD/RlXYuqCqKtrF6p2J1y2YwdFbbLUDXz0MApv3SG2afyGLb0LXhvIrpFG
X8xJ61U+iOTuRhkpQ0DFZqKX1NIkugd/IIeurMPOtwnzfZBz00c77BY2Lb8tfWkj8cLkNgO1tCke
mH9VEM2AQwfMtsLEpWbQrp5OaDgmthSTBeVBrNZG4wxaOfhf5s62mZX4galcYIGdEr3Kj8fH1BB7
iePijxGA0h/xHDbTuXwYxSbEptt1Jfk/EPysfPuGat4Pdg0NOBnGD96lD31BZ4FAokFn9uNSAB5W
kl1fbTHVvS0gxfKQWawSvpkVhGIJSTW75BGCFns/vOJoORpXLunudtH9OSVVoP1mDiFKTjA0+OHt
vstUwKwR0GDknfZBzDyD50qryi9Lr1YjkPvsKOcFD/7Lxdv+v5u+0SAjU8MrKPSJbVukJW0S57KQ
SxOkEBMiIxfqapZU/9zVzhWS/ITI8oXUjqGYNTWwwzNPPuMiLzRQ/U4bCUybDcJAxM4G5L8EQLLR
PLJkgbtxr4uuJNDdnF0PZwyt8BIxzTCqjpf/P6uKVawrXh6muCNCGJXUosv5DMH75axslD4N6B0K
TAykuALIsp3XM6UJg4HTgt1vGYj/sL0G5kxN+WkV0a1CsZuqgRDIZnr/+iZqgdyomW0bw0o9ihMA
c2mvxgMPTeIk7iFVJWVaQ9sw+gybJqP4BYI2f0TMzg8GHoc0lHyREAblDNg4P/kXH6JULn7YfNzo
m4JY/Pvdpu7PYPyRaMI3Yt1fAhh3Z+ag6fNbG4mpvE7rI3zkgh2sMy1bslqYwVyYlYi8BqVRGyCz
vqCeMxMYGzI3LflbnmbgA9FkHcHWAfokU56vT4aU8sC4+gj3KmqEqHKr0gd05/Acw4HqjHj6YEi6
YXXcZbZMaMLcXjCfMn2WHKGHrwq2wDtZRT02DAYk+L8IiIq8iGsPgnW/dNWai5rbdXNAvyEytjrC
uQZ3Z24j0iYtbRLD1RIYtBnGFE6GVrL4OJvTEyxc++z1cRhOBwJj2okD1yqLU43I00b4JWu1nDLf
d4RG53jtkz2aUXrG7lpUeI0P8Rw3cX7E08A1a1BIfbWD8JSc8bRIvkZ8AHVp1k4amHXTa4HmT384
PhzNY7RenkmbKp3wTsfS5TQj8Fec8tETZDRULHZmmgRYQAaVO8Y0FNXd67vEMONWQCvlW5m0lo7L
xSAC7iYKKfjo/A4/lzvo4ujH6EZxBL8f+axEdpj/GiZxOae4e9TXUVnFZpM1v6XP98qyKtAmi8/y
mUcYqI6HwoG8QNkQbj3SzrCODBCB6n418Ygw+tsvgE3LRLdAnQQkZ/tYcfsyfH6wW8Iv3f1fmOG/
M+WEbBkV7YHqSYMjUuPLxz3ak25spFt9lsvkOwv2STbSF3YME3eeB9RX0uyUFJya70RgNddlSf5K
XqCq3crMTk5HrcZSYcgn9oYI8iWf5nei40CN/rLZjSUPY5QsBQCst60Ri3ckQ+zmZ13V5Fiq5lhB
NJmze21DMUyJyb+fIH3WkXoL1wD9R4/gD46gdA6woIYQrFQCiJz0uTkRFifBaJmpqxfyywiiETVl
pn6pcQUI8czKhvCsNLe0cj2UDonzWpkwnCs5uf7H7ybCheuEn69uQktNU7CcB5uT0dG8F+U9/WOi
SRMDzO8QuH/aP3yLUWtygvhH3QtQR0QZTo7GCah7v763Cl/gwRwX+rUJ+45TLOGRs05UlkKYNYq9
mGCUGu7+aalE239t/W53JbpThqppdShnmFnbfqzi3dnJEzSMVKTgnxE0a/W/5r+9pykL6cpapmuD
ikEpDnpzj81p3tByIz1/+iaF/myp8zQIiBq2sOGi6wE+FBWebYzcEozRfs8DWfRyKddBygoHqzS4
IZZTXM3rh0BMVpkFam1MIk93r4FRWBTAdUqSJ++8DxkZuM86PQ4aziwZJnQsKU0uC0Bb+0Kiuyfc
dpblbDxObO0plupFj8cPw+QCf19YiB/32NT+WHs+ScedEoVV9luOsX3lfJLYxZBBt0xzdOPqFBje
fxJlX50nv2Ka4HIJimLa3DMWC2BKPMrBICmXiymx0hYDHC1q3+T/Yq/VhVPETbN9wJqlvWBnBg8S
0J3yQZl6LuBWCKmq/4sNIuvxwS70SloprGUTMb+a1tG73PTMPnu/WiiFY3bqPqfOUy97g5DDoxAF
QKcmIvKKw0jquXNqSg8VcIs/TVaYF1CoPcUADahRkWaviSWdx39PQfiIVKDoqA6Bj1P4OC15kzpb
c021GdIyYuC93E4tHVO2bMZj9qT+36UCOk4PNWfOkx+8uwU6tM5sNVxu250ndX6HIaAlgfTaVNFD
e9QhUzOzeokU+Zgnx2rjedqgkG6TVeUBauBNtVjrt6NNq2tAG52rZxM73Fm7v7YcyrwYfC4cFEno
fjW+tvlzujJsS3MQR/viB4oK5nUCuXxitw1kaT7FVhkqQvGy1YG6Muu9D89OvE7WOYQEOyMrWFCA
6jFIuez3iQ5GoLC7zpBgsA5gkAMdB5cuqjCNkhA041slaPy6IY6u+H6b5G4a3IZsm+yujBWd43WK
RDsAkc6L3wFN8xrkuGy+UlDqA42LZiqRLH05kndlMymS7IVCEBg2rax/V67/vmTD2KfCymCLiCFW
JaaoKuAQhcxXM6gy+GBuUUwgN+6U7UqHCF2I1m0M17ziNeWWmeplKDLNYerLw7wMxW10WRzQkMd3
EFLfYZAmENKzFe1P55LQsEwrYpHk1EQSqYmq821WR7o4jKuwo0XZEbd2PEF7FNIfXVtCmkAsevwi
sOpUu1Ou8aq+lNq/rKcBy4VOiRNMNHI773vq++OcoU/10MMQZaud1+c3Db0dlxBUTNGPf5OdKPEX
9IqsSRHB7LX7xM85DTdt2CYttzajche4cXnIgqCDJyMVon9jtBXnScGvVWOTdUzb4AVX02muCuTx
1ifBBSB56s/Yc+WUIXUDLAhlyk9tMjy50VTRbiE54WSErSP4i6iGROvQfLkjc863GYOffXiSGyre
BuWkF2bs0pd8gAdxYGrcpdWu9R7v8JEXSGGbWjBYm4agSxb7RZ+MqBqFH9UlCRE/0WclsRQuEH5o
M6NN5iIMxtWp0mvv/Rc53ZgM38DYDyWs0u8/fZigsfZnvfzv0yWiTsOM0zWjdBbk5uQR3psFSlG3
TUsaA2wg2L2CZr/bCJkudjUogD5MEAfUktHhbBnB7SEFNVWbf/J8fQE5l75/dfEYbFJ8Nm9vJH0X
dbD7D0a8MbjkoF1YPw4iTWBXQUI13UDrrXw61LmOUuAYjttiK4aM7CBfJ6o4UlYiRFBwZPdv8Hl6
F/4r5ABsq9JziOGHUhRQbAFJ8FCmy4hSEE88m0gFBfQByMZt/J4ErEvcm9BgtCgTog0s8c/8r86H
cb8esIpls7id1ScYdR5w75NBF0y5AjHLFIZol3RR9a6lzNWh10YIrKu/Ayu2mGVYuobv3XHV30nq
Aap0fwRFaT1cPZl94ud3EOQ66BGlMM7C3AWgXc0VgoVQUcXPAnooSj3bwLvGEVwTxPGzkqRQKkLI
4dLpZeH2LIBdwCVkOB2jUqdlasZwROHIBLT2BK2gKb6JBIR3ZSU0D1mwqkCRrlDX53nBEIBz2f7L
BXmJQ7Ve95Y16Wt6jowlkoPOUmTHAjvGGF5Hdky2GNtEXGZGl7tr9tBmyn7httjBPRuP0KwXxcUD
Y6o/wz/y2QuQ4qFIlBvkFDPdDVSEXne9u9GEEbzbSJYSsq+CcMHxljeNxEufR+NDQSNsPMrKcnYp
oa8LjvW/4DdEyvLDu56ehACd0lnm8sBT67QVrDYrnhlsaF5dyXiqh00V1+dCToFM+c3YvC30pUxV
ibrd13SLlfdTPkJ5T95Uz9ayoevKWbP2wYttKqeDl1olspZnmfHPlca2yGcfAPUk1sWqauGkKr+3
2f2/x9b0bRNrGt9qaeNcmi+8MOdFgwJLdcoWJCR8TsJgFtw1xDuh+NVAqWwE1IlzhgEZ2t43bqsC
NWsu8NjT/G8rtOKoFJmRvMang96s2Kxum5WFEM8z9AHcGZqlz9y8m/F/KYawRGTWfFg2gdXcv62T
T9k+gdTpTcIYjem+jQoQgUpysX5qkPP/2T2KcJ/Mf8/WN16LTQyxYADfwmaxXuyFFEGo6nXZKzhy
qEO6HoqOTI+K07mVoRZlhU2jBgqBENmQgZCFIj5998Zcu9eq+S2YmdDe2ulio0ucn8tP3FRDPfbk
6bCaJLzVPe6yg8yxj3L/d9Q9RGjHGFcfG1XjqNbRmyCM5Uawg0IXg9u8CqeXfTYZSkBhz3DSG4G5
EkFnOiQmnB5QZ5eDRvJlB26Gcj5jN+3XrLR/roylzaM7x/8wrw3HibGsSgHG0zVF6k1t8h0pqyOl
eymwRUKSn/Hou+YzlJYKJ2A6wrIZhE6eZ4WSUUEDL0OjdPSOrmCIn/uYoBviTNdMKWonw9PmSxEE
fMGVOgvICV9huek4gvjfTQjFmtrR3Ty443WctDA8p2+Mu7s0o1pLKyidKUJ0TrOgxIjjIVz3AWvp
lXsZ+aYECU5XHi20Fu0L7L5qFsS3LJI3pslnN4A8lCDveN0ubR5RdK8C97KJMwuCIBg73w6MK0Rj
UeTahSlz3lZsXmyaPpgxbGK4rr5c+Pc7Egg/SiZne1tYEJGV4XoEkWNeCEfctxj+rfQ+hR/u0Tlx
ONBdlBuDNDGESfMHvlhRREO0KiujppcYxuYdk7O3d7/ucXnK2dqOb3akQWq6xClxj3/rdxqd2ru/
v/n//Xke4/LEgMGL89wPYDwG41zlFJev0I+ft0oiBJe0W3dcQgt8d9pw16z5Q7ksIxsmGyQKjtVq
IGvtOb8ejWJNBwn1Voc3EEK+NQOWRvurUikmHweHyZuG4ZsHN+whnCRt83xYKNk9U1ZUNTamOV5P
Uh5RyrxBlFpC1ESRDnQONEYW4c/vvFz7cHqzDBL03AeEbOTsJv344Dzpo3sTuKd0PR/lEYTYPrQx
0y8ilUOzuDcR2acTkuq0fvmpt94wi0ZghumP0kYay+jGJmSx/YgFh6W7o9YduYBCgDrRSSSsOh/U
x3j1qPiGtng6fh9tpxYYYzEoVp2GVuLb2mWf6ZxULAyip4wSaUpkqzQBqkmOWIU6L5ttr+WmHfqG
RO/RyCb+Zenfcj4A2zsswfX8PU11mnHV/5PWaauzPO9yygKoCSKZORwrHvs5KhKa5bNFFV4NyIxR
QLEaj71kNqkLFiD6iQv4E5NPCzeW/SGlvUzoR3aGYpVY4p/q73wtQGTo/FGztjkeTaACXu76KWrs
/jJkDtD8Zc/6GtQ4XclOaghDKbNpN1kU2lM25cWvD7sMJVB5MJ1NZegAhi0oWYC/FC0Qhu9U4IvL
xlz57ot+EttQ1/Sz6O60wJw399sn+oQsTS5y+/AzLYZmNIf/WaPDyzHdgnscwzb87c/p2iSZ//Bp
OvYTgCDJwKLxSZDb2JdakbslZnFXssmSEi09N2Hu4tsOpJoHpuirUpC5PYOAKFztVyMSUnJA4RbS
Ebuyd5vBBDCNum6DyA/+EErB1uLFJ5AASxqT47+WJW5OziPuLyqMzR9do34Rusi1wljhXCL8YI5V
irPL+3EDQbYsj7Sw19IUpDPko1NscKWtJrypiYHtYUI3Oe+v6Mlr5jDrbhKdIXMbvs5mHCyZ7NSQ
n3CzJtKRfGZ6leJR8Z7C3jTpZaJ4sTg4ZpkRqn65SC5wHQioSsBBPeErcomJp2xP6TSOzEcBlO5P
qyGjW/aKdPh+TchH9U79r6rOFFcJb10SpE8k+WPgIgMXEyD3InrJly8RNlWnMJacXoshx1HAYqB5
H3Qpks2Whck7Wxkgm49Dx/ZQbrYzLEvcNlhdNS8ErluANXbnfztSZW0Y18rSt+EnpgytJvA6ruiS
fpD8L0RqfSpXDFG93dqJNnBv2Q3te4jBhhpgPdHN3++COIKBAbb3LkLwE9jQ+IizhWVPYsBmAOAA
II0MHBxqEYcXcLHybASeOpViUr1hR+FYV+k08cxhZhd3MpyqiXAgHHioG/B5VRPCCgiItO8xWiH7
VhViMxdsP+IoNBd/4TjnKqp9wxK40oq4jSivsYMfrOGijkXLXgdfjDIlxfN0z4TzsZnyaCbaHyU7
VvT7UOEpeazfJ79BjfcdbXDqQ21q1d83ESpsDXNDtGhQVRcvyrp9rcgtiOAPBIimgJewGZk6lEDu
d4CIg5M0KUq5gIbKss2wQYUpU9rLcxaCK6OM2pYQMM7AHwaBcs0qj6MKaES8rNbiuF3mWlcjV9XP
RW0XssfXx9dhyft2AXp2kl31wadVpM8jVVK+Q39rr3OXAwnLDA0yjnWaOtN6MsvnOmkWcyoRC/9s
2jNYNxeih2ILQ63reiCsWDNMOHxNEv7XGzx7oLRIfJ8haCR1xcSGeZQX64WZa5prMlml2weTbGJK
2LHuExv97tbP9xuRIruyOFg8gem31cZgaKY7cw/zXRIwbh98vHFOtV4+lhhI7jpXdbivdk6qUObn
1atvIUiqvgvYbQxvtNSLjuTHR6pJALhfFON3IuLR850vCuG8b9EioQDYBLkfkTfMz3t/8xzeH3OL
PXVDBBXNUqDzVwpCjawmpn8QopwWtLKf94c6hjo6xMAJck+QiwWan0hwegdxUgP4ZgHrifxPknuw
Xy5WdZDQkznErTvyTPZb18zZQBKhp0yCKf1dpsOhriO7dYm5+FhGHAG8VL3L/rI+rdc3aEjpxeo6
3bwUIya8jvlrKyfJPAxcdjpD6++pxEAtto8uz9aMaTHh22OSn9JHWRMBeoJk69ssxOTdHUYkLIzZ
vOmGZ1pTBHkKAtdKmQLO8IfNLXkYn5XBpBnQH4yEmud+Qj99AFtjzgbSy9RcPkFrkqnRhXeprSY4
mghwnk1VSYXMWxcgkI64B+2xt6ghpU7Xlvrkbi8WJCAcvzac8vIj7vLeeC36Qd0qimgWhnChm/1n
rupMlt3RZdH41I9Q4saT4zJM349JBnkklpWTuNu05bGwFUCBqPI6LiD9xVys3FLi9PgKbzjsrBql
IH4P4c/k8fmavh6ZwxuWPGlXwxpR43pzmp65C6v/r/GEfx4Y06Iy49x+aIPOYjMWp22j/KnpDhQO
ARLizsRVTL7C3ZWzxADD+kbt7t8WfZXSogbQC8BF4zpqRDxV+r70g+rWYHJsNO4K38NVthBp4kFO
taDQqn4R/bw75q0AbnDKKTStrKUsRXzk9tv1f3SoRFbkyQVcrM753GSEnDfPI4lwymJFeedUjJR0
IkjVVqJnm5oeSQ9L5yWFq8gS1fwmM57StPTlCT+3CldembdBGWYe1KVmHLRA2ge+jLhJpB6ijOjp
FGZcGWUF9YETiop4cc3bri3ruQ4VYE5/Y9Pc5bBdFW1LeXhvUksiJ87h2S7QPFBds/Bx327vYc2p
hesITgUjaDaN9VFPMNHJqGPVmOHAZ0ThAiHI+1JvqWt0EnbpbuWGRBwPHXoQCL8ER/ZWGsvMwGBB
vF6x4t2ejNChaxdmfV/6A9Iwocwnare9b+jp/FRWgP6JzGJR3ZmWVP5VxnxG1gmS9w6tWCeU8ACX
VSJeKrVn6h4AdVXSH3fRE2HASY3rZB+67LCSIlvSOGJRhvE0DFi/kSXv8i1Qs98F3c6jMr6wY+cU
pXChrOrD1EKd1K1/303kNnrkaiddrJar7vZsssuzvOBhTHtp61N7vd9QU1/4sHfREsvX3ayZA3lN
E7pI+0N8tWLMi20+10/d+/pzwTgNFzGmP7ouAKd5De1OltEmJYajgV28bt3bKzFudrZGmO24sIQS
JXSsmEr8CnRcmxX4BINR535xA6JCBfDMYnHrBIT3Xki7emM2xAMWTmGUA7hd7IxOqJJkndvVfAys
50Flp5wZ1RivU6CFntTRi05pOYODkEXouCnRE4EIhK0nelqXEEwSLsBOgWNXWiHetvl5de2DZQzt
KK+GaRsZC9GuSqQ5uzqMOTnIkgU+njVu+jA750DulrZm/6wFLAGOuwqSkQG07zFC+bNewrGR7oqM
p1NVDURSALnn6AhpojChvB7xEiFQmbVuP2GQKVDbkB+xWoXt6Dtl86MoHqXuRyYFJqEj+fRoJSNJ
ja4A4v7Xm+aDMgErPiNCArfo+m8esv+hpX1Kpfz5znt8NC3945DolG5Mr50YQmtwVWOED/0wecpD
fAD5gTYUh0ZWlpSgbOS3S30/sHODxmv4rsBmr/AllM4asHM9gmVVY6D6Y2x6C9JgFT/3nDnG4JcX
twlcz1nZ1aPSWfa8edltFnWtzhWPidmlFithCKnv6w8rmfPgve0xHt8VlzzMKgRrGmABT/kMSr3i
L7WwfgFRKuSBQnDN3da26GpKZc0+E6XNVg70GbPEr5YINvSo20j1QYJKBvBfo/JsFItM1YyR9Q/3
FGTbdxlrSzZL1v3TTLJKWvYFhtRPq+zPeFdaOGHJpyA7cOJkjTlHBBw3YOXBc+Wqk7ilKS6gwloq
EjHhPXqvtoiFVU5lzyhMm4vjyTiYeDVNeaxVYoCoF0YJs+jamt8/4PJX6+lRx6esqii33GuFu2BK
LU4y7BZEbbM9GSxznpjhP2tC9mVd5gLPklaZleYL4hVNK6sU9AUbtBFaVcz1S41pFdI8MPIns8no
yNrIvEneQSb1DxmflCfPHpO8CME7QGkWXf2yfK9sPn89d2+vyCnjE8V8ayA4G4x6PrNOIZ/EhJFb
jZRn38FhJ5l80gWd9bDUKTVWMQuxSA9Rps8X/hsU/eGxzrCtSEzCqeGF5KTFWl8HUUjzg0zfyanw
9Im3XsiGHgxmsVrLBxoBjmnKJe9dbWNTJuzemAD5w6twY4xzQH/JCcCnDDOjWBAIPrS3gWzLm0iF
Jc/9HP7nDeZ/54IW54GLb2ML3JQh+akDiIvgJacMSsl3QLNF+Zy2VL0QLo+GKPevyusUw7LuVOZ9
4GTAmS+YaxPubEgfydCnR/qVohwoWzpJ79XPd9FzVh8wMNAZ8Gf+E0gjL1mlsokWXSozn7yi8LJL
vI4IRRnuU+ZsrWtdnpG3KHHUj6ZamOqaf+ahK17U4jwQ8mrGC7ixEMACsYej3c9r1mHWX+oUc5pi
WGpS9HG62tj/GBlPtY7QnB0D6BZ+dQvtwuRx4E6NWOFl10nQbQHQyLOCdILklOIrYEHqbMNVfxo1
cTFrYHMrrd8UJJjiDzsLb+OF9MNGarj6vTPl+QitYrnbetpZ2E9ukk125EiBtRhVo9XDR10S6l/d
SCLGhXadoqWN1P08QnWhcTy727J4klYjaU32rfE3WDmqgVYMmWpfpJ6tOJDCsTCPf/iNoDEMpZj+
TcmerZ1mnDZonJz9gT0+5b3ZEHm7vNTutrLUbB4Gjq8aJZhJ2P56kEpCmvgWNqVCfVIuo0xCjYJH
TYGdIZadUW/W4ZKEgkYW2SIH7BoRJUEBi3RfiilbA5+AJ/5w86Esw2ZH8V8DTmtYEirRovT0/ApG
M5/E1jW5EiSnmsDlDn6CcDbzeRO26Ej7pY46AdFLGVaP2ZvXCwkWg5ahnDxdNDsYIwqoxL72Rq9z
mbv9Qqlmn8bIP7pLxtzgq5W0JvzknDFANjSE0MohipXdOjqxQBu+lmS5gDAKVj7ysvNbdKytkWpm
n7x3NAZsYQTSbYYEg+LHhz7oKmkf0YISfPe9Rfdg93f6e9m4f8X8wbM/cRnOJuDg2XexpNMSlkk4
GOvh7IPmS3LlNzbrf2GR9fi0fHmxE7hZYv/Cbg3+OuVK8So4RKJFcPGhCukRxevge6Zk0yy31KrJ
LjocJK7NQ1pNzyt63YCCQiQM+IYcGdU0mpP/HMg8UeimiO+3aNfXKSOWnmjA/3UIOvuVR74H6yfU
aA60vA7eO/xVYznS2G+GIBsoV1XGpFRwjSQPesr8BBabd6iIgVeUVBD7DoR16kLDKpICyxJ5oq3H
fFodT1WTFAuchfMzSWY8OOhliCz9vVHREJddY9wZbbGW+iTT/2x3Us/eCccOkJSof/HYjpT2tLDV
NvkMnmGar3zB32T0NJiNwyljjpjTho7c1GJlpWqh+51CljXGl2b4mSOPu4ccgEIsTeoIdLWOKRqf
0V/nEDvCb1EHmm5ghOmVTx+s8d7GfjENl/0DalpIOagAmN7Z+wmS44GB+mnoWB8RjJEA/nYPeFPO
XiVABErxoBPgq4GbvFU0oFEHAM/vf2W/hXRufic/mIkmIeq8YPb9Cy0kdWc/SwGdlV3ibc0Dstxk
4V6T78UvTUeUNJWi088dOgtEHE9tWqdBuITS7G3oCvBsvQD00pYC7KcEiYl3JJ8jKschrKD7hthr
5OiT4fu4ADwbRZZxrssT1t/oluVnZqf+Wr3XhlhyUw0QcE7BeoRT/SzYjyWhpphngHXf3MmZKMoJ
YwLdYeeZ+CeSPYP9rRt2qJwRX00aHxac3s5DLn2qPZ93KUbzA4j2bJ24xxKE0WppJj7gJ4V8fgzY
3q/9/+mPZgKqVrXtJzfMJRWsthRKv9O5O4QvM0VGw4eBMvpD6iXZrmsochcr4j366CqAyruEgNIX
R74vlV1sNubHJmWq9HsI3Pj2mxhxHW5uM7vT5Moa47RqaAQuwrttmS95KqSVY3cOFadVIfrgPfcO
HMz3MIKiayKxlNr1oLXYbDuGt7pg1njHGUDBTOYZ94rq7WeyLlEhyYlH4gpsoIKBoFXMWvQ352wC
vRwmbWHhCxjyLv+s+FWPbWszjmciFxAovWH88FFyqums0Por3BsfDHhyruHfNsSIc2B3U7tq0sdF
6NgauLxTylN4pjnciE1/ZqN3ns7AYHIsYJFVFuvVVQHNBoN9IMDL7bxlKrgW4fINsoDso4QLTobS
WzuvWX2kkIZXz8v6fGb7A+yVDr6xQiiUdnm7+rkzhPqjw2qnzsIOZA2VfOAt3e5tqsN/iT4b6zUT
f6LT7WFJjty4DY6yeqUlQeNtU/8JyBpYNPwUk+krW17EPlwKlZhZZmrUUP7k75O+LKLf/+SyUZ3a
cXYce+MApVgji/Fl2GGoLNddaXPaIbuQumEqWGDa6jttOqe3SdisuLZNlJeAcnrZ5kSlafD+1au+
6R0MWBCqgwwb0Io+FMvswin4I5vf3w8gEzdxXIxrx+J5Z+sYCptciQUf44IE7MDxAJghSjEr/Kel
8fvo+QvLm7+qgP78WDZtrqhlMhRF7oD+n7qvFmIeeYTh/X19YVaTY4qZTN5J2CiGHoesD2Kt5taa
o7vAVvP+Nj7cMr/ZZ63V5pvf+JjwZbU9w2+MSbCxM4196JINpMlK6CEYvOA7fImFvMTA93/piirC
H7DOg8v4LOvbmsJU3QHfHxxJmiz3Qo3VhNDdOCcegJmHL+Pev2WY6XqJqeO5SIB9Xu/wDwHkM0Wg
8Mn3MlisC++YHVnPRnTd8GEa9Z17ZFMLDOPpxbT6tGDds38kFXU8bhkHqiUXnDYitwBacaxZXHCg
U9XSn3BydHNdmsOIf/lVcseWmGWK0w/XHPYw+I743tJN3Dye0USP55VBQZWYfZQ3liwk9nDj1U8O
BvCe+8FYbvxWJ1wfuhaWjOlvur0AbqLVrElI4IL33M9BdpUC4WpQvSvAj7+dAUwKwa0VWQA2X3I3
/RcamctwddQr1i+Ep4dHLCvKBVepWYloAZ7cMyRPHL7TY6+dJZoGeWajL1rNjHsHP+nYGnkkurBv
RfIQuCZSVcoSOm47/K1EUPghM6mtirJP/oTdJ7p0FuW7k0c9HglqlQt9OykEaMgUj1pm/2nWn1Kr
+zdOgkqFB4T/MLV/r7tXNPs7/iFo/GXhWt1E/lqdNycqtcIviLJIyYOQGDfc5A3br6RwQrA91Y+K
NWWTYC3GhCDKcapumWxQTmKO0FKM11SJjr/EgUczuRECz7R7eJBp58ZwRVGfsX8TYAi1YzMtk4zn
Ks3chzmDwVD0Psf+XkpwIlSEoXVyti3JQ4K3FBuOmr7+l1L7sb7jjRTsReJGnYzwajbXQbh0LWqc
pblf0/R5fiomrrkRpB057Wzvunq/an17MSxR3CK5m/66Z/KXoYQ5utpuxkwy9jjJ1NvT/i3a/MOJ
cZstMRAQB5F50jnx5/jd+t7ddz+Iy76gS6cazM3IqMHa1AHUbVgoBU/+zgl3R8T1FUXHeo7dq/Qn
Nn+AlztLPy6mkb5LimExh/0agM7TnM3QB+DMyhdbEwtqE+J83mpUcx97jEhU5ZVh0Vv5UgWtZMAE
SFcpGgl8s+uQPPO2s8xwvtocNH08r52xqLNUywUzphvYpTTehtxF07F+96gD7nvvSwg+UujBCWFv
70JoXOEflEBqdabFDS4ua+DF2I31740RmD3Ow1lVqQbKGy3Rf9v7Ih5atCUTV5fVea2eo1ECmVLd
a04LNl7pwGtHNq6Ua4EqO5Gd23nfik7qJde8YW6zRrq8JY7SZVR/+k9Zbf4P+n5ML81mLUN8Rmwt
a3oNW1wqM22NOzZdSwYVDNMtURE6PHjTAiqw2VknQeXN4LZ72FN13TxrOgYEjmh8ioGNvd2nTl8q
Xle1lCedyR4xMjyoYgeVpTPfzDhr8jma2cHaLpViWO9wkG8rzW3OZ70j1mCJwFFhiBGs+1I8IQMr
weeCThvbKRaarFwwM/nMXYkhRrYXtsAddv0TplyWgjICMz6o84+Lr6wFrcyRBjGytNU4LKa5Uv4z
oiiLRYHPFP4RwtosTf6mzVtO78tSf4e7LnN47nauxMC6AHdj0n+SZ1ktmPovcls8Khyofp6S3um/
bSwFdw6nldXTeLCsqIG3IMcraOZqxVrdwqAm4LtBx8ZF8GM15Q5LYoWk2TYh8jHz+cdWeUAuUj5y
n7mLUoc0H38EKzexhKdbojjc+UvjfP3xovdBVv6nk/R4NZd+sletcpgDU2cUeZzyu2qTL3RirN6c
9DgvAwm4Da/+3ok9trLc58e8S+drs2A/qwkH9tY+Ls7ubD3/85LlsOEIxg7L2GO5IoW+eMyQqq7G
oguRUatE3VMNRmf6zQOwPm0pztKfcHTwhhCZLyVdOgBu9YJ25HynrxbrnGP2Bh93D+3P/TkGSX1F
RzvpmaTAZKUYtGF6eY+eNR0DvZLi83kTAuogDMP1oUPH/RNgAmEXg1rmTeIf+vBTVVWY7EYN4rf+
hqprZ6VRlPpZUkPaczrYzLBCMBw4ZkKq+IBd2qOvifksZCaWqduAs73vQNyaV3WYOrBUWmeCXXuQ
xXwlAggIRkzTDz2UWFko+vyrQ/IT1CKQ8x73qR2NaYqkx+Di2b5geQ6YX/bF3LIdSF/kb+4J5dPn
HItKsJTwNDnobjTqqg1PbRIaR6dRjUkLpKw6Myd6Dt58p2YVlUsEIJJ/reSyhnMO3CObONKmvkXA
q3mTP5dNcl3e3ifbvN9/vkGDcPQ4aWBqBcaBl33Fm2uvTYve2SnXZDcC769qgk4TPj2qx2kptqJl
1CZ77JzCOvRmAH1vu9eu9aWQOTGaIsSZnsiJReo7g5retjYO/9pAUTMqtMfmK+VPVhKcG6AcBofZ
ZpaagY1lvlFsbiBFNkJLsQP8RIvz2NX3k4vxcwuYaxRXedLmAC+MlMsK1hoSuOS7y5L+HJwFZ35/
oJtFg8xZS1Hz92EIcRKHBFgNNa1pDK7cVNveuTQCQNxzPDrVX+zzKy3GEE7kNZTcG9LshF30FmJV
nMFST+nx4SD2lqUOAAVXCylsH6ms6YVkgL6ZBNHBRcrRuYz99OGYasGYHWlcYXbtgA97qYwu/YBL
NoRwuyyH3WN94MK02ZJIue5wb3mbWbAHWxt2D/sFcOuWL/rLbd1uqbJfXYwtf0OcbFfzzPnJ1kj/
LTjdUI5l8z6PhtbZrFEi3ZNoFCZcaSMDAOU5Ry5dRCc9BEPoy92nqX1ft5TEPva+9ODx+F2QDDEv
KOMJgW5+o9zPh8t+1leytVjd/DtDwXLvkpoYVfkjgUgtD24bq2+RQI8/ZK6e/8u2grKLwDmEaSf8
pXoNbzCLMDQ9d4J2hr+0DEE4LtsCYDAg2T2vYfJeMDp+8BxRjcQyhaKWSoWTyT6rsVz0gbxDy3Wz
ZCw/gpMpg33zi8k9+KsTCidJijVdsmBOq+6vmrkKPSM8EvoznjYPPqllv+w4prSIASO7/wrt4r+P
FgxQym60OalyMHLaS8eYj4DH/RE79/N7QC6drnreJCZsxWUvqXkDOURaZGr47fV+cxlOVgvIs1PD
7k4HudM+HwSN0Oxd9fb44Z/re0jTFyWFMCU9pjhieroQjdquUIgBLVmjdm3F7WBmGsVhcIvYQAWl
wroPR2INTymmIdmhr3vEMjfsFSsKp2sbhO0FRygZOh8LCKDt/zruqJu2sjTY/WKfuK8Do8Q5FATK
2ZaCYnEKIYwBtUmKE9S4fN56ymmqXZjNTC/2/KAuWOdHbDsBn0iyMMkwu38rNgy0ehJoa1ce3GKO
hgtCsQy3X5MGebnv8xqZpP+U+qlPmWuWzoGVzz1PbEd2xMLCfHJiOBONL1ELkE7vGhjOocFMuKbC
x6YvxSEbL4w0LX1mvt38h0T+EVGoysoX5rlCTlWrQerqh23zLLoWJDTVdZjxFgq74Oquit2ugGMp
6VHHcrnj02hQIAXKkw0FvTPXT3iOq59qjK8DnweYqMRsiy3QSgAkhcjvvzQ9jA6Napw3C5WWI1N5
zftWKOMbiSGYXQpK4qf84sIxHS060hnUlRLgBZa5Qw2iEXNjG1eocWpacGU2L4vg6ZX/M9HtJT3N
mm5IsrY0mOnw7YirVPzmfHMCgy5di228tlDiY1UuGk4h1MLKRcMkpjJOSfOno/P37RklqWspvhz1
O8vuPecYdjtsePuCMsK6w1+gHo0moHCIDVXI+4PNpARFMq5XsysIdbWr13QC4DvRiSbW0vu2lkzl
2mbugBF/+4m70bDjODxLPy8SOBpdVbhFuSRJq48O9RRjsmUoFQyULSRwHwQv24srmhcy2h3tmP1k
wMXmF8AMnOqRXEg0u9bLIbmgO6Mhcy479tgsNHktS8Lho+7i4sgGQA2h6cgSMqom6zEw6zRb9AHA
onIoXtcpD4SeSVaDDl0Th7EKTthi+Qa55YI8NsfO0QGD1rqBlHEjuJqZThBEg1LpGi/bYhO14FEx
bGS8Nz/TxqyKDEKROIJMV4bfyHkyWYM5YXJaEhmAb1l2QqnfKBzYKSOJV5rY8mzDa8uFtbhD6bnw
t9jovQWeG9EeLTjaozwVCr5YU8s2I4eIV6cw0tNuDudovOSGkEnRmwuIjLLw0/NEP42ZPqWZwLcj
rduo0Mcz2Xi0l4mynzdsE8TsEryZkhZOZh2wlD3VK7IsPKCEf1a3Bp91Eog8sACMrnUcSakvLah6
VTkFYP09yurX9f6JtTdf53DIwVRamhUZcTRHbZGYtoZ5Z5ZwIP2eS4/9feN7zooIN+Pu4HhiM4OH
fB040xcGaX0XeKhkoGSIO7HK/7+xrIKZAVIn9ukQFV00j9gXOOft/i8LS6/hhhingTdRsv+tVJyl
tg2+mEd2hL3qHtnEwj4NMOF43hKFQA5w8Y1XMW3jXHAJelA3PCD4wAaiDOwt9l7j9GErHt8VRVCJ
XB+dXKJ65gznlS4hpZOAEpC2xN5Wj+Hj7lFLuSGk3AL1JkoSS/u/xpVnyzVJvll+Cn2KYdzsxOTA
uoKwhmodN+g7FyQHz57W5T7wpx5+smsaocaEDu5NFd2mp203EXZFJa7Tvg9AUKJ0g7Pt+8ZCASvm
dJUfksI8lsuyFxkSs/pL0Dx0Hen5H+6qBSzlNvNJvL9zOxR+1SU0pXIE5QQ8Zw+pHnh0PZzrmbdY
REaag8lz7r/HCtzoilA2I48sEusHzPBKPuiNbAFe+JvZBFmiNqF31h5rxW0gCzPnDtiQi1qNeTp2
SehLWBD7PGkIJ6HRkM2CwM+h+ntbiMOxNQN1llVRmkqnjb3XAdVR1v4qfedNqs2NuktW7+Nj+Rhw
tjv/Qg6YUzAKlp/P5fPQQOZlgF5uekcwSdIHCXlAZLk71DR+uUOzzxhlT5AHCLSNHTyurN+BKiVi
2qB2Lnzihol1RPeqBZCYnolMQ4sbsDZd9CXZGaO4ATfec1i91oMh7LxLH3zYhFTfDKaDNrroRKCg
NiGE5yc0wWumPWXoYMUTuLyKLo3JpM3HKr+QuVxCKK18u0p50BOvaKsqPly1CF0CMal6cAzaf8tI
Mlrx1FxaY45jyRYBW8UlJnR3ttE4Z2cAgAme4y3/U5XjVzBQkRZQl7e/G9Q2wswbCOwq7j0cYiO5
XvOUcLVi8St5MfG9dMTX3FsoAABwQKceQJuPjYpJnp4q49UneD31oc1uWiJpVJwjWw3kjBy0JOyP
7kQRkU4U1AXXpohmUpw0P/uC1dQ8decaoya6uDY5xBOcivKgMiBLdv4wdxPLqh6PYbkAsWoRLHvH
Jqisu1ZOXkyOK3VEoo0Mx7hzR7MaCUwgxP02lcV/9JxgboAMDzBEXODOEiB5tmUxcOJ/Qu2lYfeQ
5+FVvMrgEHpNrGPwworPfyENv6cSthJFevfIlElUyS4d6tqrNOIOGkrY+5ik4JS/5QQcxG8wQ77s
nuDjPIxVjPVcDcsDIPKgroiLfBOvmjyN6NiqwuyQGv0LjbvbnBu+TWHg2ZAeC3LjC3DhgMrJ6ifh
00k4w/hqMT1+mvR0Fg4BsjmMUHZLTrElqiZSUQ/7R11h4Q0DfBusBpnOKlPtuP2UgzdWcupT93Ib
TpOVO0pRNl9ajf/E/jcLqIDOjlNaPZ/t3u3STPQlHYWPrZz6+GxZE9ZOxE2EIzFmbYE2ARPesiAy
rl80mio7T6JKaowoWeTuBf3a7Nr0+Q0xoGfhoY2WwSH6hXbvWpluSoDPekwrxjciROUx3EhOo0Q0
tx5+zzJOYIj/dtuEKpYyNI2IQW/ozNOcPoLznrKSAvXfd62PqxMp5McfBNyz/I1yJFGFWJQGZZRS
I+XHv0lcuEQf4OrTwRPImDsHFvj/9ppYLyIFipv1fMBl8SpEbuosT7mBAeNnda4dhQaxSowsSw+a
oafFOI9voLvryLG4EB36J1al01ndbNhe2eOqyhmxu+NcQCBf2X1KewKGvGaUL2srdTqVAubsQIVP
U/2hbGx9pIVn4gen4zEuydLiz1ap0OJogpANxuI4PnYLLH2faYSin3cbMrPvxnbFAj0rnOEcfz/Y
A4fJqpT78slOnL0yJPsSJzNiBf57FxcrhARzwPM1cJbTpQePA7CHo/R2ygJa68HFC6meYy6d36k1
H82UdvKAT4+EY9cTjQyiOnDBjGIa5Krj2cx/fSiqnsSRvirduI4HdF/+RITVzWk/4vCJrumqmNpf
rkRiKwD250WX21mRL0bopwxi5R0F3yOaXBCkrN4ET025gL1IJBdgcREnOj78M3za9RcfpU1a+3oW
AiAdKwrF+WzI7VT0+0CLF6hK/E0v65TnPlAtIxO+kAZ4qZEStwL5VZdhzAcFEMwZEOhIFA667Btq
+HLDnI3Ii2N8PC2ieT3EYsOfhgdkT/jgQXpSO8uEl7wl2uucManrBDzbpk40/QGGPNlpQKAjygTb
UyXmRds94QumIuWFjqnbfmmV4LiYS00Jh3wMmNFqIHpL/FFOgfhkmSahqyizJJoDEmQeRZL9oPCg
ZRKfCJXOAKfdY9JX7oguBhdgjpTeL0fBXHj52EL+wTat4xQblktAq0laMJJVaApphEv6rGM+bzxc
EIcmz9qg0cJ/mBNY3l2S8P9kQ2SRoVm2SD1Fm4DzPad9Rch+zR97Ztj49vyFK4eSCk/pU3CzNzY2
EKWspZE4EAduz+SVHMO9BcM3Ap2SFsAwSHuxI8aqrcRvOYvg1PhxP/oDmhBK/RgCQT5FMLvMtxyi
eAbxGDsjty5GTGSiJo88YCBYcPJ9+XeSqUSxbuQFFvEMq0i7a9K1y/NZVJjaegTVUHEOpAh17RfZ
apOrhSKG18Nsqno2a8NVjmiKMI1b0WgDIj5u3xyrTUw36Nb0+LFbmI+5YR57raD9vIu3ahDqRrDz
1iG8bXXtKc0rOpSYsrHbhO19Vze3EEnvWPwByr30RDT7E0d+pmli3WWc5/xbp1dD0x5sg3wJKCky
gT5EtdsdN5uIPXECc1qiV0RndUGwLD9JPVp0uvmNlcHaokdrCWHlWK4brl88Qu1QTRWRQ/JCjHH9
nDJ2uKurwrqYa/x+LYmVZKsWxA6QOqh3O8qd4MN7Z87maDq5VactMKBZfVOVuktxQQUqhbm7d2GP
E6Ku+TnhFYLnXuPkUJBhbOuBa8K+FEmV/Of+mPSsYtEwux65fcv56ysb6rqOMVlJRKrLaZ0Q/6HR
hvo5Z4a6Yw/LmldAYtoGubWWLBzKNL/rPaSldVxKPgQCuatjXZT/4F4n8+cTMkCyov82a8T4WDn0
LG7vgNIdPPt4g3dWxttjDxmbZrkINZ53/+pS30eI2o3NL4n2qSZznif0xehIf8S550AvSzldiMXp
sk5H5BDHaRzoCnS4nphbobh4aSHMHI5j1xymJ8FSQdHdapoVZsBeiP6lVDhcxRyfohkDRe66N+8i
TQEFFJ+TBAnQEIXo2YmIrEnF6gLYIkTjnrmFkCxRjG1vuXmLjkx39JcZ2VZtDL3TlbbdcjHoR7ZR
PmK57wOd0xbKGshxPAPeP7WIVqZwP4sNIdITLrebr7i0m41AUowwIFyWfuJY0Ht084pjP5hLbh9R
ATnmzl+aGomNW3QWdqUEdTsExV3Ba/H2sfW+SV2Fr8Kl0rOd6WUDZLrgEjd0oUayryPdvngq4xeN
2JTNnT1cx6C01YLa/zcC73CFQOiPQHGZW503UOAZRw4TQQahwKje/j5BUfA0EwATgEPqdecrBXn7
giN6qakkSRPWLGhb69LKuqWCuL6Ip7qu9UMvM0/UIjIV3cX6kuU2k5MEY6r+3aWXZIsMUER5Vge2
Sxihz+Lb2eM/FeDcN6AAyUfDLRRlEQLKkS+qvrZYab98dg9UfQez8xICE5rCP8f+oKeY/h8DjhPK
ERxABV9xYXaLRnYA46jQIou7wxF4cSiiz4qTWdsAKd7YzRiLrFVlqZVMjuoe5lM1zpuGhUpB3idF
ZbKjgee0dxLY8plUdCHQSfLeQXwjeXR6WeNcMjsU1gV9yyqYz/FdqM33vs3zzWukauXnnnsPm6SL
MWNOUOLz2jP3O+OzzJkqb7J5yd6g5YqUmxK/SZZWJ47mznpMbGjKNdLD3jpTskhOdJf0wiy673TE
FIpkfqNVgL+HMM4KNDvpDr5uTo8UH111X2DwbAfiA6jc0qjQHBJw/vmm4EW/EulI9EX+VXDHl3WE
6BigzC5MDE6BKTzrwoKufKZP3WCEyBvwgiQyLWxtfMEZ+tZ0fBZZKDR8xT2WssPYWoyn3PMmmIMn
NiK7DQEnNO/gUZou4y4WdrlHI1/LYSnNdu93xl0Um2zO4zYlyXyJw58xLg48ag87a7OqLlhAxePy
1EzNwAnO1jJxMb0XTvMjE+BGRj9CMCxe+LvGiSfJT0vFN4Mkc5F1YzA+DnxNsLPW0WUkDVNPdn2r
6juq6VHj/zLyOrFxOuRxeFBe5Rz5iAO/K3MdznjRSzK0Bt/hiGZGmWLh0BZrk9l9sDIhxq7Ohhwb
S4WhO/fGvqgqZdRAfiXxPlRuY3jKD2CRL8e/GU3e6pTyxNf/zciTYxGfnbpA3bmxlGXefp/r7D20
vFZwMubmTDF52yK1CxQCTVvK3EMvx6hiAiIsdl7PAUh5qz/yiKT6UGaNG/jK1mxSvJDQ9/ulHmd7
UD3uoeRfTgsrIXvQTzTSAeclCUoLf35i2eQ9bhL8rwrT8mfzSY6srRpNNl5q3WeAhkIOJbT6Vpc7
HjwMI3xeOSd7fcgZJCYCxO7VZWOLr+mj5DCZQ6PneruZ7j1LrRdkM+dufe9vxV79g6nBtd9tJlTj
GbxNFsTQUJU1Di1dc2K1hFT/poNL29aSohbTY9M4UbRRIIiHswbHyCETZGXjLJh00d4P+pCMr4ax
ry3das/kYliKGP1DUje7exHZrjTGP8SwauLDiKhu7FCEozaHw4dU9/rChzxsQe5OR0cDDcQliOjd
x4sFFm/GZNIWKOKQ0TUFpex5bW36JhrjH48QID0GisJctg+0Ct1+waFawLooDq3ig3HtGESb+/RF
NXnsjiaEa3rcJaieMEUDBb/xDKqpN9kgBUPoFrBFcFbijaJ7DK10Fjv2FwL7DR8pfhdqbPFGCNBo
SJBLbK0k2WG8akC2njLOcN+9MtWpDdgzL0mbIKU7iVYTYQQAreDKPHW6lSj4c+xWRPAVKBEMZ4pr
TsH+KWgQNipFX4LGH79sURZ3YdqB3X97mN/v+XhwgdvBOIYBwcg6l/Mf0jDZSN+gGgcpF529nOi1
TfwvqRApa1FGcTm1TjPuf+UtSulZhHbCFsdxjZSAgTySZdD8HJj9IWeyJDhiFxlC+rgkU5H9A1Fm
WyutLyisygtig+n9JNGN8DLPo2/K/LCo/XGxvTcujQ7UBKaaOxPsU10kOGGCmK77mNp/ANNCQmtg
VFcAW/je+XPI6nuziwD3RoiS8ztCQFF1BncC2BpntwOFoAM1VAEWlSwd3aOeqaQ5UwE9H/+94drG
AmdfwjSDiTOhjoTkxfubtcs9AkLJ3bTHy+NeJ0FAyw1SFQ/jIcxr1wGxNkBBPIOY6pA7dPD0a+i5
e2hK7qtjIrm3m2rV4rjwocjCyeAMAwnk8XPvZqLXmDRl2VQu1pQvMtz/PNNErioNRvVa4T6bjUuv
l4D49lKdnmu88Xxx+hhhENa8xHgT9TiCWEssGLLS6ts/h9fUSblGIGQL1ZsV37hN+s62Itrly11/
a66bk8I1ud01Vt1q9Vhe0SAbSK2BcqAVa6KTbcEGN9XsdROV0c6/+L86TSkQeC96BZtkF1MM/YI9
90NGVD43UTTkg/FN95tnXkDB156FUxJNfkxUwQR0YP3tjY/1VOl8IVAD2EKFotylzMij/acSmCjG
M3BPk6mTO+nfY9D2Nd96+XwtDi/b5gQMbksBRT5ywouartZ95iPTxMl3/YfjESl4SsDmoy6wHwtZ
44gS0Go06VWNY/BqPGwRX9dqnP2yRCwFdx4rKdO7EH11sosbRYTifjHH5GScHNhxRBTNoM+jIpwu
ong8D/iNkwPgFwfBks0+cVdVMrrPMrQoJJDIB7j10ovQQ+8SLQ74bFvIMMs2/LA6gAkZC6ZQZNL4
NQKpE25KcMEiGB4qI/DJSxQ7U6MQiy9hqq6JmjbTEKLLuSQwYfgB5YFYN3xq+5GLUOfgzWtru1oh
K8FPUoz2SxtXZFDMezZLIlO2xXMDLe/GTnKjJuA/93lD6SRNJEMleDlpLc5V88c91rgN4HvQp0NZ
wXKOtzBx0W5CQGc8hRZ/pElbtlrz56Rrm6aUfgrKdeKWxQ54rgc1rF2cNZiuzwc6h7k91wbwYKU7
aH4WDJi5T4CDCPBYujKPquRYYbA6Rx9mX1U+gS7d/SlN/yM5pSJ2qHQ1BWP5ZB57DH5Ob8A7I09m
5OaFUa9G9rEjxDVmRYsH/cjj3IiE55B2S3hRcyL1fybvn11B6GjfyZSlxojop9tGCfJu6bn6M1Ek
m82A7zVrq6GA3a/O2SpIWvjP8+NBuH2NIbkkOhU77iHc/SyA/g0V6AWY0tTinYiuFfL1mCmASvML
J8xlukBcTj5Z4Lx33kkRy8sHkCs3iWUCxi+ImSse3Fn7rlP8LGuApJ+antfisDEFg0gSdWG0r018
eWlc4mRIb2KRJF3DverrPA3hqqE9oJ43OT8QYCJP9triaWBOTq8u2AGwfnaybkiVJUxv4xjGcn3b
oJHwuU1XQRhJjzN816g0bykGiGCLXZAsKByxq2neJhqnrSC/GS3tIhvXWTBPZUGBLEtQNSTUzCpY
GEL8723Sm710T6NWssbFvne01Bw81rzcm4qk1KILZ1uhD856UHfJyH453Wg/E0oVeYTeyPTAQpOj
Y9TAgKqntpeEAzjldhGyS7ZR6GJg/llZrFu7XYxI4mfsO/01UY6+tp6riDeon5uw6avEk12exaJB
+6x1RO4uKfH321DzuBz3SunkzlybRN8pDl3loMocyxTPJ4eSdthz9zOtO+HIrSltAo2X0avSrTll
dm50jfEbTm4eIia5+C6abr1nxZpokaUESVxdulIol3nVQBM58OhasWQMKBxH0NVS7c0MNMtIUWEU
WYBktaJm12hzV0Lks44iAQyCanFh1QayZEdRu/IK1Y5LIH4467hJKS/VON7Fq87Uqz/Nv0XkWA5t
/rDGVtqEfaVCd3iqn3F3g8ZdIUm6gSh4L1f2qFDQfjGRv3SeGXv/W07Ea43UZIzNDVkJK2hZ9nsq
j2AsAY5kg5qz7TLSLTKnshXCsYi8XvCngorr1olgUBn0GCBjgtmDHu4K8Z2HjjnRt40mJWsvVt9J
Q4OuT60Zu+R2wnPLEejQbXokG+nhtZ5dVOgpJeUyGC7k39B+d++iglyxqZnABCTYjbvKE1UuirT2
iSXuuaeUqgJk3Dcs/trjej42bdeJ2Afq4FXf6OtahdAvE4JKY3KUxopx2G4Mu4M2O48PIvRp7vEV
HfaOV9Z2rFkEuZNPbFUzexCOPY8btcdMKIop7zHcsw+dKrJpMDiUiJLcDkIOS9SdSXiaptPGvNu/
RlLX7sYJ0eKKEg4/7elrV6CcvjR9dDDG531yhuf9i6I3B4nSjxgMhFdz/jwQObrrnpQKUnZwgR6P
Qq9iGj7lByjML4Wj08n7t0nIRkihVQC8n17KnnqJbzDzREnjrlC8lnfNzqrnKW0f99peA6IO/Au6
9QNp+3Lc0qpUnYGu4rK2WivKzQTzIl5a5h7PSj4aSfopmKS4MQZR7vZomHON3Islb5uKUiaiT0iz
BBRv8E2g1QHqphGtfyg8Hh23tubJ/jp+3+ZkzLtpZ06+SMmybi4qXlbqjp2cfr4qWGRT+5OnXLpD
E31x62IQH4bdlEacfe2qh2pOAZA5msaoMD+7oFmP1xQGpbhl8U/2YUdz6vT+h+OYVv4crZ6q87Ke
UFSbknggEwFEdhN6huABvN+Q08vV6eSTNZsvZdfXoFTmrJDmpiaIqECy+b6QofNaF2yx0NFg/GuL
BH8vxPBfbFtxa9+gRdip9PzjMYTdn8H1pmGLQPcFso1pkyzrJY57uWTA2qjYFY1WSTA3ZDjEtVBf
jKTgYKBRZpF5CCWK+HKTu559+wWl/lJuuZqQPE/xKQILBJXRhlpao5GUTn/UselP6pLt4uuJl97k
BjlLXHm/+OorRQU/PNkcjN6tYXFnP8RzHVdFK7PwAOONWtLAz/PjxTADDi/YXeqqC4wXAligwh55
ub//n35DwlMsHG8s7bKN171fQn3vFyQ2iE3bsSsxzz6VB2yyGeTSfKp5GabXcw7DoSzA5ZbZgT0V
rvhIItaB166iJ+nl6CZqAu3paRh/An7VVHK50K3ChFjMBHqx1d9z9AlpHySa9RhT19PQq14LAcZb
8mrVjxCVit1dCRbc650LjyppqbGXOLYm98337nfuys0c3XvRNyd3HDSYz6VaHUnxoIeTeF+TaV+N
iAZ4XigSKFpMDq17X74VAfpAQHhffa7gkrLdkbv6SEmAvWGb506WTS9gfFw4XpHz9YV9oJhLOlSC
MCnitq4mZhEoBHrXApARCQpDUBgUCHz5MqaAwnTWx+lIXAd44ji0TOpOXgfhmH8xEW8q7J7HOoSq
bdoB/CB3MabUUvK69H5DWn/56WSrKUSIDBy5AIGeOpe7h8bspMibVX5ksZDdWBVVPzEOHYS/TTXH
84xRM9h4f/Lijnyvb/cDSjiNsSl14I5hVcGs/O3lSDNIRtVMn7OJ2z+e0ZN/vXY67g501Z3dcTK8
N66Rxin9f9DaSDRzqyPF9P//SEUmA1ARWMwZiEij8mg2NCPdMLmeOeifZNH59vRj6gnPYHY9lFCQ
yaX2nEFYZdn9eIlCtqyeH0VyeecVSvSuzKpesuI4yWQrcNwT8rYpLiZXbtQbBfJEdR4tMoffjiAn
xeZ36PxpaCv62Afr/LxrIBc4iP0WGFykIyX+NLsx1IpLwb22/Ud/k4pfhpsv40RuINzULNOOVgih
BItJE+IWFLbqS74hCwATSDgYcLs3GVZKAyHoHL0FViY47+AvQotxDlYBZ3Tse3W9p2eLpUQS/hxP
5aERll9sjd+E46JcJxKFHwPZfVmg4I8j+CoSOv+Jo724GeK2guSIaJcHEWoMHjgtf9NwHDdumUr1
1ED/5xTVUZRDAUc9Bn4/5h34cowfXwR4k4xfLXOvbtdEjqAEWIPS2D1eKYpGNt859InaCTilTDjN
S7iNMGfkUA9jqjOryRWXbP7FXFffalO652Bw3BIZCAyETLAym7qRdeLnkWoTI3p7IsaL0lbbnxZO
x2Ns6vd4Rl3/T8qhDsY8zqk5gj6d8Hfxd7vms88A33/kqSatGR0dKPxZBFBw1n9gWwe2zqiAzRnN
smJBw5rxd84y2NHHUgIo6TCOJ4LuaGS2tRqfFjFu/R9Dfoe8VQmmgOq34Mf2vT6fjV7w1xArxnEQ
KEOc5sMMd5BnO6TOO1xorvknp3/gAGaS/WkzlW5A5ZJn6UFyo/kjmhqs9CYa3ZT84oL+p9rRbJbB
1hW1lAPh+897POwLcOFSal1D7JztSwhRtjtjnZXIg5zqU23HH8yKYa1n8mSjnpFZ/6hVi5JLhC1A
NK9HUi9pAXb/ot4rNIiIABbDWCZ2SE4XWpLrGwVF7MeLIr4c4tV6nGDl7IIomgS92pgzs8dxS+19
fX1paKVhH356osodoazuPkYNT+5m5V9NGEfQd23zvSov1fS2vYthziTvh6ysQw1AnCuedJoopEa8
rMnJcBlh3+uH25CKxCPCStT1fCkVUYxTTaZ7RdBqdMq5EfDlDY7D/Ki0BnSf2vN2tm9FufcVRZTO
hQIodVIJPXbseXusocxwrzOWYzGCxDVpkm85ig4wP28sCB3mgmB7PXP7MMWwoLh8hTNukEMYyGZD
n36KYV9b4FbcKVo4gLbEpbM61cguufME6w7Tj88Hur7uQw/1ng6b6F+e1cPS3ga3nP4AEV7FtdyS
sZNu/5olBf57iUl6TZwagGfm83dZNzqqazgW5pFJ2hfsBcvXuyiMrbhu1JFsc6UmLizfQ3hXnHH1
ovT20fWh7QcCDUon+78orJtfxu5sqVpsHCYELfPRYwS50tXbMeP9tTqrVqlcMqhLHoa3bqR8YMPI
fa0f5qZVViIRXnNkFkRrdhdCGrwnemDS/BFZyMIveiSM36022kfQCJ2gnA2yiXj/U3v6K0W7KjE6
1a35FYd7KPh2DVrLMUIE0Ul466uF85YO8QNQcQSzj+c84FGjxgSYahIbxvfgG6tvYQgI0IR68oDm
0h4WBXqTlO+omCpwDdX2KZrndCAkFxoeNsxx7pXOhheSqDtiUKlXJyelCcmhyqEfmIOhhtFTnto9
w+wbxvMR0chilwLYvW+9wCR7gojqUEQHLQnBKhmbzKFp7mqgmafd41hnmdUQ2XDv0rSrQiTiKA38
mEIMU7dN6a6yVAuQVT5zTcx7LCwEI1eZbCu4RmPcdRmnFaWGRMxVJJFKNOOf+RtRDwN+IcBlf7of
2VKBnPk61ArsbvXa0mvKywV7FFlsT++BS2sxHhfe7evtlo3SKGKmlKeN7fPy2NkoDg0sGy9zUo+3
GQjQnzRIBRqocbxhXM2qiTflrBDBRfDWhIvF9ljETQWG/jroH4KyuybhwHocfibAHN2Og78WQz3i
lSVwg5KLi6uH/SJOcNRPhWqWGvs8T90i+ggQou0JkCIMfDPfiRWfmXnfu6zSNGyqOU1q8V3znYYS
zNxoPpzYkjheThIuyqBYzOscd/dO1lyjSfpEhRN6Yb+69q8W/aul5kLlJliIk7vTGVwY2LtZV4Fn
R0Xg+pf5PBCBpbKAhVixzobUHL5i6RxhcT8spay7AUimFzY50cWcbgbl2Dvc2rlcsWNgE/ZIga8o
AZJZ4THUmL2hzAxDAMrvgjx/9sox/waEgjmPil4xt87VLp4NsRuh9ElLlW+lBK3w2seTcCQktARP
Sg8tobV4dHas6sfx+1q9QdkQqtaDi+VhBtonKqKL8aulRZ9kWs8IH5t9TiRnqduhshpgEqGR//QP
T87n4yoVln9FgjSDX+n828L6nlWWZZ1MBzcHZJdhZ3SWDANPiswjx1e+z9zZTGCKGTSlpX1ricUy
fdCZGGsRXyTxYOMGE52jSY+EUxM7ipsqwLwfhP3yV/ndEPFSrB5sq+3lGiRXZDjgWfNTsF38JTki
MSUofdBKWIKUdcBQVnUkhkW7p7Jy4BN5iLvTBf6n+yCvXGEFj4iH664WqlQ99MEFe+V0xa6LLUo9
bccd4MnSAPDV6kxtuse97vkQ7+BsmPVovKt/M1Mw+6KJTnKMnnnFfM7VcsA6FpG7Q+G8rLGR4Mo5
J4hnXyHAIiocXznhR2Lqjvro3r6wQ07bdFesPveczRQ1HxKj/5sHt7y9LqiYyv7/UUCmFsEELoa1
Uin6Fs9gAraVjvOHkU0hF++3pTXwMSprpNQLzap05X1C5OFEB2k47LgEHxQX9KQdUtIn4nmjLVop
MJe0AKo4fxPEcO9S0WIvQ9SIiWYaXHsdKuUv+MLZTfqc2hB0p4qQi/oPnDv7rAIdeZSgMfaTxwkN
x6LP/rEoZYQH3Q1Tj0toq3CHE67UrHAYmnuiaod9MvUfGR8Y8NpVMKoZIBc/UCy5bptCJwuQS4M5
VAyi2orABIhwg7a6Sl8aaCWq1wzHF53B82kx1mVs3S6tJNSapY+1d5yalHTABr/c3Rx49b1iq8JT
B/BSgj504Rs7Ki8vDzby5CETqS8hMckPbGrv8ZNLgYVAqJMr07VnvlL0ULPYYSyxLfgQyPPkhJW/
6iFAVubiIFJrEq4xlnzx3Y+Ij+4ntvF6va4HctcWqUTrR4o4sebLLRhw8i54hpBfgFSo3l0h0XzR
B9YJPMYZQ3QEHhqqcPzsfJKkyrnKkyonuKD/sVFwmxW1j57ZTWrDvMfdoFZlPjl/ZiZtC4LACA+1
FPXfZyjVmTarZw4ngCHKOeZuHoEatYv6Q1IyrxxbZxkTfdqEMFqeG1nV/QeXb/NIc0Gv9JBs3oyL
HiuV0szQZ19GpAUdKlxFqlzFY0cCWSDU+3awsvp2nRDLk0YQXrRr8y2toDLvM/4tFLSQ18TUqzZC
P3cezW9uccotnMB9pFjmmeajcwTtrlR8f7pWwPB8Rse83My9O8wOca+k5eMNR9daAK3QBnVqxJV3
u+xT3UCieDXdsgH/Jj0o2MvcCMhCC0DyE9+0NDFWTdLDKcMnPLlx/t0d4rdFjuDHUyexQxxNS5SD
OwCdZcExpXcsxQT4JmM61ubPkSsvvlWcrCqv0omWT3FPvT+PJ8Bs/P6SM2y9mF+g7+xta1RBc0L6
7E/uraxl7pOGdOICESSNInl0XPnHh4kvaSs235xYX1a+VELxm6OvfCM2U3d0Op5t4q4Rn1PDWR5i
LLD5RJ76Isp+DfGfNqpz+8Hf84k//U2KDd1bliSZbiQ0fUclR/MS55BZvGJwWZTMnLcAB/kxVCXn
JDEQ/Y6YOTRuwPSpBhcpmGRq038Gepzhat5f5N332ACZUIq4GxlYTybQx8lc4o0N4w2qcUF9PKHe
Z4/n/flXF3omO+1ZUzWciI3zfb3O5qDKPA+cv4isXuOoEwuRlis+I5v6Tqe1vzVsW0iVzhLP7Zvv
wRlhOHtA4IJAH1FXvEDDs2ZDQtwJjhuLtSVII02SRLIA5nsUBNAD0lYyviMEOCr38R96pDHtfmDG
xVP0jX9q1LwS8Qfywza3xpIQx08qhKdhQkmSTzdg2tMPBPd4dAUpVyr21EdTcssAi6UnA8agnMxs
TehqBDscY/npZJBtVu54y/COB4X+G+fQn8woF5rWe/ixLulutbGG0fgdroSTgasdeyKQ4FrxQ0tt
CoO2OvV2Uk9iPpKoVtbZ9G6Rc5dLDW3v/6CYkDJK/u/xfl5GvtuMFjS5Ub+pLBsqAYZC+UVoRIH/
wz8C5x9emN2Qs70FPh9hVJflzgE8Yzv2KvkY1PAkc6Gszg3IXcZoE9SXl6AKV+XoeeQvfwcQ8KTI
NfLQsb05KdNt2ixy3yeqCy6vTbY0jTRUwXUpzH+c0R4il1kv+GAKA3Iy+zdcRuNbuTQ10RMHPJPH
WLpTQ9WPUANdCBafVysm19bXyLnV6o4PJMRXDhGVGm11oqqBaqrgJqobZjoOkMlLTRUvdWus099v
RgIud/tA71BxyDRg/k5xrz+csUCSDgj6XErSImV5SwUei0Fj5x9ZJncRRHcI0qM+J64HK+UFnQjg
MTZcQNI2w9y2Km4xiBy51JbnP3sR+AHNJnFQYdkQUyLR4IJn6HDKzz0K25+lbwDp3h0ZavfylWJK
JwlX4TgGU8EEeGvgrQX8ZaLSb+DcfkPVx2lja3n51dzK52/UY0WgFrWwfASMTqCx3mSXK6KbkJYs
2lPNcQQdnBveR7l+3hADt+9KsIYI1gXykJ2BJX1Za1dJO31mleFy2BFTqYgMYUHkQ9BUALUbVUKA
Hw7sqMitzd5lNgnghvmeprq9FGovb9LcseProYpOqQwd+cq0+2Na/tVi5MdR1IdPn0lcs51yaZRm
YlaoXn1njsibMv4WiG+zePoAjvecW0amceuXFJXvCtQq9JQ+WSqaLJ5IGuC2ZGkFHpCjRjr3l3bH
0lruNRYwfqroYD4sbrv01X84tzkWtiw2rHr7B612+9ULpbUAjFM1gGKJHAN0GaXXxuf3k51W36Eq
96GPHjY6aWH6nDdFwnjz1Aec7fE3YLHFzO4KtMd6KO5swTSIDIVxAirdNyQ4A8xyur+2hjr5k9HX
sQ+GXu4F9H0VWBpe6Usf70fiBWHAUOH+ubUXZubjF+hzjXT6X/gDUP6a/NdcY4PmWQfIH4FOVUph
qImHrhdQKezgvU/QJxV5SFzcEPznV2LvHqY3zmOLM6pRN4mlzFfVgsrjgKNeUavotZtoKAoaZ8Gj
bkSNP2FJ7nEUwVfwYqgJYG/hx9ss/He0AeKMWjwtdCJmT9z9PdWl0EvWgOVuOqb7jmY/r8J79wGq
4wa/eIStBdnlFi75CPZ1HXoiHJAfsvL/VaHHMtqKD9hdLZBuB0WY40GnotHpnGawJL/1bIpu3Pu0
x38SNociJaU4p2XbkDHsbJ/PAD71JuogFWNUQz9K13EBsVPoDo6vhNPCMqES+FYcmqzk9fWrk9hA
qc30bvnYveGT/VUtSOAWMzo2uVN8C2kmzljhSCiT+dikFeoq5SEfsh9XCBKkhtJCtUrXYrt3N6tz
2yAgCAvvlY+8L4TEumXZi7PQf0ejPmz0shi9SQUCyhFQ8B9/LL+oy23WqWg29z6dylWcgR2iX4pC
gAeWLtVXXj64LzhJFrV+2K0uA1+RQJWhgdDY+vgWs4N8sou0/BPVNFdE9iwJt+wQqZc41NoYZnqK
hZvmz9ARZzX65zym8BPYv2NerTzDMuoeHe3jplfWLeLyYEKLD/EBDSgn6roq2aiC49Y9yczkUnea
LBaejDzdbGfS28vz8eEW9+NTshu3tMskb57v29Cq0GnmKA6T3FLx616lC6q3Qx3C/LBg3Mco9VQ5
5cv53LSkofBpvnAvEE5qrhVeD3bpz3oT5+SSZxe1nncNujQ8ALKXEucRiK4i7NUSryLlAuFhJCKX
HyXmuPxeW4rKr3kuwTASVOzEtWQH/zumCCHBlQueRdVqUpJN/xKu8UIDO4cQe7D9ApWeHMoGJ/+k
uwMFfIKiJYG87ZtE4ttpHNeLD7drKpuUijmC7ORnNtK79mjJXywxSAX/pvDLlDJO4UqL0HN548xU
rYor7rfDAKF/Vz1WdEMqZ25WKMUKgJknwCriZj1AHNGopPVXCR+WrIQBP9TiBl3tQEab4bUbVYd7
QYhZkwkKpJWnNZ9BjEz5mLfE9/3YJot617lxbofhGwj0ot1yCkHEz0z5Tk/Y+lJhb5yUaM9SoJnT
9nDecVp1MDunlhXfqJ7xbHa2ywQgozkFHDd9GDD1wJdA2svq/Ug/kprvyxYvQVgiaHiGcm70uFJU
0V1afsxq6faaZ/yXi9VCCmX0CK8LUvcM2biBbKLQXpmuuABy5OMA5GKfnuV5w5vosPz+989vlQS6
eVIMhsIhTMPaUqDeaqUs1UxCHLMGX46aozWXaVv8KyK8hXE7eIJktl6Dl7rOonWFFAfCv0mUQ85H
b0HEV5aAd7zefGx2wL1XdIuyi5XDtO+CCttf+l9pBJeeDP2Xgzo7+t5BS5RAfbZlBPmLoRyEATn8
+yTpujARZsV4gs298TakXHHyqe/Lu0bLdViGUOD0BsuJQEVkMBZVzPbFZ3EybrEupxfKGxTGDFcO
lt4xCLlwVQOU30/+G6W4KDoyVMtpdRESbOBDBV2ORvojOWdZD5ugqh4l6b9dgZggrCE3XJNAaTRt
lG8f8hyosq+YVTasdmeupCaWLvqEdXxnglxighpGS6Wplyr/Fl7cSZVfNJRgtX3otiCJoH3tmC1U
uqtbzdA9HTH2fqq+Ou4Ug4REbFrwGy6tgKNbx43s2XZf7bJIKD9qO+BcnA7Z3mhFcGv0SMlINONm
BkKOpuE5sb2Kpfdb1y8bwPtFdVZIV3b/DYD5oE6DuI1aFLxRkjrjr5rW3vdUev3+GFdyEy5PM7UK
UniAJ9TT5SNgw5r+CcAUmgxo8Th+zMB/w56zukdz01NRjS1aH2VbD5CjXM4IHez53wycq0LmJmTv
Yhk1PUQvikCjFB0ctNTK+xB17XMPupU9TQAuxZbEuXm6dv5EnOPAGJTJR759rywCLwL9GzgIvq9u
DDvnYzb+mEB55Fr9zz+b5YAvv1rW2KE486bsV9h5QY1rHxICNHj2iCwGyLKjCKI6f72UBwtvn3Ty
0fZ65H1EsOMJUJ6pFrkAdjzcnkGLqzumQVX8H+U5BHtf1BZ1zwJ41WBoh8ee7ISHmkh3DJg8QM2+
1SvEKfo8PaS7QpODBQteMzELY3oy0ybk+jW8kOxNV2/MZ3C5FI6a0TWWqrxCqeySgciyp09StJNU
sNVtX95Y+OnLQbDFfzG45FyvzxhmDbo7smyahrAMYeXrtwL4hGp9CzJ7MQ9OVdSIstJVWypQG0gH
2nZZEmC9UWumiZzugYOyhVdme3yJ/2FJ+ckHsEyTh7vxpVTDPzkN3KjvMuFeAEfvydlcSSa321GB
rXA7ILEAGBFaZ5sIV2CFVzY/rYf/dFNHXXKUe7shMyDmoiW8Ff38Fd9W+dsQioBamffgH07TeJ7S
ZQSzLYOMzisIhOtUUEY1G7tvX0iCBhsAylOEr5RUlwY/hU6OmuE6xXaLQCbE9mZDDWDU4LLC41SV
fw0ax6+5KaPIIU2jWG5/p7SlUCI0Yxr3k9Tj/1xSsiwIkIWcGaUIqq9OEGNf4Lf3+JOzgqWAhe/V
m1sg8KZQEOjGXQjEWg6ZeK3UylgHDHFEF5Cf7vz2Rn5ygYQkDV/dGe8hrvp5GizqakojblrVhXqC
LLw2Xyb1R5PNZgnsUTcNgXa20FB3/j+F9UORfgcEQgGmSM8lRrh0/Gf9yViYdqiHw0KJMDc0NiMk
VbGvpS/yh5B3dbz9nkhXE7lH/v94vgYUgT8TWEoo/PSho+B8VVSgeBVMz/JdcCPLDuiQtPcnQp5r
MFb3+ucm3aQHF4HOZ2vBKmuRZakkdxs2IaWepGFSUW2GcUGOAuZ57WPwULB7alW5ogVBtolrBnXb
iaZkcbCYhkeferehO/NG4m35/qW6uJ9sGw5gAIlagw7KHUsy52gtBObzBLjAhXJEWekfp/0F9J2n
VfUTHhNrOdaaD13xRB1ZUNdZcYFwajTuJDPvhRTiMNhF5TBGCovZfaF6nXAj43adhbT6SZEXnxx1
7aneKd1fzaLh+RxF4gzu6DDbLyPhiKbZ0kT1t3NootQVl4629t648v60BigDBYVsTPHXL0NOzuQP
DwhY/oOGplQk28cUsLRnWqfkm3eWy+kASvIrZLCJ94NXwZdS8KpD4U1xR6GAPDPzscxiGi1lMmzu
UzCZPtqWDVIllqtQNpul977kvPClzF8uYkamX3YKew/zaDWbPJGbuDJo5OIE8phQTojqdC0rq2Y7
g8VdU+VGkQEXjWXGeGdFhwmOJE8iU6l8NtPU7FpfjgmovPf11y4RB7NWnGotoFafYDnGuZoZWE30
8N9JC7PMn9Rq+XlE/P5gNbKSsjIxPl5yptvVKRb3Kl1Fs+FFEawfwKSB1a/oDhH9kO+dAIFZ2fWE
ILW04j4uMWUu/l6lE2QMcdDdCinH/X4mP9rFjAGgHt+brt/xbZwFEAe5gIR2d5t09DAQgyHt/rVG
JgrokflVogGG6TqthXV1XMUmMlZGlc9G8TdedQJArA9WEwq/RX3RdFHGTPQ4/mtstqiQb/XkiKaf
LkZVRGW41ELmh3qCvXGXkfvGDAVypknqkIyvFkSkN6Tmp33DrwKBlhgM6XM8XX9RVcSf7fkdeFBz
jSX8doFVbH0iYihllb7CAeEcz2MoyrptPq3r0nlt8I7Jj8OjHnkCjWe9qQ5kzeZ1hP4nmn/23SXH
yIUrYDJjA/MJ/QFAH8aL/gCOLovdpq+DZGb16CMvi2Z+Ol9jlZHfZ/JfhdWDzr2pmL+iLyBPPHRz
ULhbSCYgZ4A3bYwLpF2zpvdsvxK56xETXEUUmIqNX0RPmhiLCv9s9es7g3ABDmmJoC/bMq+u5JNM
s8jVQIZpUeXR2g6qlX4tRXuXaU8S7EpGl/IbCkhIxXxcoKZJKounJbrEr+nnladYSDIFg2wQoCAk
7PnfxJt1jI0wnrcqZW6voWyM9dcLk3n+N0k3BnQrsoLTp4AQDbPSf03h0XwPy/53auzJluTOYbXZ
bTcd/p/8SAayfgeUZESHKkXbYrq9wjxs0x8g4gA2Ke2oXgDSVZpyySfYI+LbtCUTo08/MiXQNJZZ
npMtODRbIB+x/ifo7CrUT09OZWymQXJ5lDE9LL+6F+0DKyFYxeU1snCUaOHq5V2LuCFN8gELy6pw
RWps57pVYO8HoZzUFD99gKhvFMEk2L2iPyuUph05eZ0ZrgG+RRKTmEQJPh4gDS1iJJ46HS0oFbWH
lXPak3F0qFSE2uk2HYKmjqQcLaRm6zM5TijF+W6YekMLVg62fyVbItHToXdTC8ATmxgmctD5eVrb
75wf475jvAIjVJaVPFDuoh8+bXgQ9mr1EYcfweEg5KnZ/bCeLsM5FHG4GJXeAhzoWwT5r3eCOW/y
PjcKCJ5oETLE5Ru+ZpbSTWAEjFWR0fEfAFS2JRKGI9gkoKEQvHJX/5bcOo+mgqn/+jaC8Ile0vSR
rFb3ufGHh8uLjdfqUHoPeKOv51xilP3qCFlTLJzFlD+hNZGcd8PyrY1L97Lfgf4UW9X2OvE5IzGc
a0liF99aMiv6LJztoUYZmD4jorsp3gBrKSdBDMSsDWOX4ahaLF19Ts05ceKlr/bwv1hJCcMhXqyk
0twbpknCISTmrnZVvfzIT8PJGouPlSJjGh4kHyVUOq3v6iAvCFQZKtT1C+FSXuzbdptJaFFlrkEU
bjqlTQKLqgeKPO7UtGXmz3l+wXeUNEmkAJaPCYWHT7kIzFBxeW43No03TCypwtvcSREjBJfTdiKZ
cH+8xtW3Ds9pPtf3Pt8x1Zf3BS1ijcG0gyKX65OBKsLfeNTfDBfaQ1Vfh+2wnArczu4ZASw5aOav
gqAkUq7qzLsazGd6/7BTQZ6sSj0VFjIO51C4JPg8sDuRbVBRup49H7085gbW5geau5okftCuj/Mm
hQjjMfuBkA2TDBhnaIZAny/xCcp+7SKZhh1EQrNDGZ1pVJnnIm+L1uWtzjG6BTrZpaiyyeE/ps+2
vhp2AGCrgjuOPCu7Jbs9a7oiFZHk2p+4Fp07pU7wGF2i29qmFjBpq2nxRcS0kDQUKe/IQMUXIVos
SYb6QzpkZOyjdCOMRqXHICwGvdNYoBFMTTnhuhVCw2uUmuSawYtRLEWt9AFAmMd9Eca78MJ1nyby
iCt3zUov2Z6uo3BCl2VldftJj/nBmDbDOvoeFZ2N7uanUqtKHLt7UKSZsdSvAa2zouY7/kUHqXdq
8a8uK6EWeOdTcQlfciKcXOlcpilBibsVnh3lQ7hCdlTFsD6duYpl7jUo3reAo3EKxgBxZo9wzB7d
MzOoaR4x+n+jPk+UVJ35IJZRbmNtMcYm9BwvjzVOKxBDO0aZV07AsXsYTWYw8w4I1OdZqiuBRsU9
ZilxP9dTGYiGnsbkdwwVETt/2V1rmtIWvn4HucjiZxByxoPzc8icG04VjeVIL1ONsgxPu0eyo12f
MAj6Zmd0h+vLuobvQQahOhSJw2YAKtVb8lP0fNBfAnwQRO4Kjg0iTE3MxVtCcIe5LP333CE2w2fS
wpAUsG2UXp5Da5LxGl/oigp7zWq9xK5lkwdf3aZj9ZVskJOggW8Fwj9VilAa70JORUEXMLAgxbR2
lBYZxIVob1K03r0UdycqC+gehnLPaVySh1Qw1AteEHs+6qOBD4rO5gh36aE0AtGQxJuvu30fJK/h
p7vo31hZOCn0n9Z1WWIYb+djKQOwp9JCWD48BAd2t0WTB3V7v6n2DMkGU98C8qOctFpID4piWpb3
Qct5ct78lMkUdAQcBu/tQSc0/XFfrNQYrv8v9eDjkAWixGA4PmOjpLNQMrLyv+12t56+2VFnEMTr
VR8TMmfPXyyhmT1rNLqCyZr3r9p/DhzuWhiObpxDwSulj6tI/FlNdQsCLDeDLlbJtKmvsA2qMUrv
qP+EYABdKUJVebxODLWN7bGLJkqofYkVnxBNV4miBEQusM+gb1m3fmep0TSO8R+A9Ad2NbBB855c
UH1OhGAFQ7HVQl+GQ0b7uCNNwml1Ticbdr3xOdP0CLnygpJw9gTB29V7aZiIiYtw6mnh+HM+KMwq
0tnJhUx9Omsekdf/os+dmFzgUjsNJfzXu8f8VZv+ajo1H6FtUYv5Hk19ZSFkEmlgmMiyLpwE1Re+
YkjIJGBDlZZLKuimcrfmm/2WRwg6puIsrh6gHzkKkbwueVETgOZkoA4+te7YLgYPR9fkiYy4PnN0
Woz+YxN4nO3qfYFXeH/vZ421j1HNxa6ZSiNgeKIhvcgKIi8trzauZXTX9IU3wfMq0+SkJD5zkm9p
uoI2+ak/5kjAlb+Mxzc/NSrqIOzLlB9QFiFn62PbQXEMxhZE8FusYrai9oTerf7CW2JeFilQ92yH
ptZbfjUbStAmGkcsR5+l8NXiv0ycJUtGYKqxqrA1G2MJnweBQNeKV19ZnYOFIDBG/VfAJBwofs0F
e0aOjsElawemw9Tx9gzljl0QSBa3IoguyGlVae1n0GGEV7UhshEOwIKgKiMgZXvC7WTp1JhI20qs
h0vJzh3oQtD6dai2kOQWjLuCdn8Gg9B+IrqsAfp1Ft4ye2rAur779wv0arMxWYHjEGsK/FIBP5W6
rjW6O0HBKGEezJOYmiauH9n/SXBISyfIMvgOT0pdwbjTLjqUszHPMl3X+IxcTum2iPzwG+2Xa5Jy
y6RHmtKinKQulEdSVmThLwC+5w1o4ilMrRSAyzxlIuAJRyxWoxV86JmZ4fnu5lxuQztxGXwm6bRV
A+XKwKdjSSnfFBTTlJhAOCvwzP7pEoIheyi57iH30hS8YxEDdAG3OnbXaxr2GARNVzvp+yuGgPYg
+MkU3QpEt2vaRhV0yiN5z+BRceHF3UC5XUoPJBA0cxIRgWNjNI0pZYnuhqMd92xYT3cUyl29pnrs
gs8YJKEKBj1fKdyIPhguz1d9AYTYeNdb4heXfYcIMI7Jg+MuSA+VRElzJfWxpcyuknc3ZckJ4ajs
1Ll4SBjs62i38yAgElFnJiev4xgWFE4gkUSIKI31PezjL4tfxrVd5lqf0rwHF4kWQcJnKhP9/euP
UwSgECnrpe8jhAYvDu7mbY1T38VEHDS6naD7y8FL+PqzFV3/NPtmuWDbMFlrzcz/IqVYDcYlkbMJ
tqdE+Nb7gYhnXYA3gIq5her/gZACqh/we4r2c53USpmy7VGPRVVIBBFP6VOwtksKEKQ29jOik0V+
Ar8C1T3DJ5nqzLQigc34zi/71KB76ffMaIadZycVHx2yA4QgeMjZEYRXmXtOhE2ZNgFxtjsR4McU
Jjx7Jg3OFGLo0vpwekHTGLdWvPLhk1SSn+4MPrVSScQSHba1e+66JouQSNNWX4HmrVK1TdwEQQ9R
zc4fkMD1kJGkr6ageV2DIgpEZts/vqHuwbjrg3WWaWO1pPTfsW0806EnbpTQ5D4WPiMp5Yz3+iDh
rlBotGBWWk/R+Kl+XqYY25+dW5QZCZ65wzuxAMZfqFaCjEQYoojD+QeJtSULJ22Hbq/ral4HoILA
ctKPgfZ4h2yaRaxcjYeayqHu6YZBBkA97mSLKJ23r1T4X6S6UtCXBY5X8kuyZBoTrsnnORrCcnTk
7ctv4yD3Af/CbkO4Kyha86jF6vsC5jqYfEkIT+REXPZwLo/Z5UbMgIs/8oAmGyrGB/OYmWSmlLMy
aIFmtYsiFU8IYlR1fYcKKqqILsSvqlsUTmz0WQBK+o1rZe7Qmbwwe9w9mXxDHJkpZGHrwDRHVqL/
lYlzTKMKDwimJ1p5Hu6rspyEkyIekoeM5vWpfKg9cFEcXChtg7GwGyie/2cDr06gnO3kOad/QAeM
M00eo3+wyQ/fNtmrv3EQP0LlPh6jwXrUj7XcWJlGvhDKVHJta07WFnspKDjD/cf0EdnW/2tuNJ4z
6Y0r0rXuIwnJ6FzMR8gDbPrj7Nj7Qxy+Qkvzi/lwDgTbYppxftqQqqigsu8qwh7RxSDIlyOacrtX
cwgiTaOHFOyk8f/xsW+S3rAsVD1ThoUC9qIETn2BVlGMg9AR2YB+wj3rpawDkzlc9S3lSFPGKh81
XpGyHtRSDmr3eKMxPGYu4WPXr+o3fIItyucgTUcbAv/0XC+KufEWIq3ZcKmsJyzTThnuwDE6+MNh
AOeBDp5eNlfb+AUyhGY3oCJK3ZHMsI+uTA8z4+eRN9H41Yq7OGSqNOGL8FVUk6X0rrcMB9UMv6Gn
OyKu+zr6brjpemk3GsBHUI2yEtfD3CTODY9RwT86G+d0hu7h4vsO2NQqMQuWx4Z+Ya+Txtukt3Ck
7SHUMgLUihRbgrCePCT3RBcabey+DFb4KmEYBmUQOlJ4Pw+Wbo7D9uXWys1vGx1i0ttrB/Ou1QOr
2zEs+6/lgf9IHlr0lp3dF3/XuADh3hITxN0BMxG8n7W57Mscp6jttjUs0uWiXPdlKxVWJH5DJJYA
l9V2iOuLOBPT0Bp1hosfxmlz6EoESPNDJo81e+u/kBG1DmPXViX79rkN14UkIvisx2UM+xmMICUr
xqoMKg9crKfhA4Ilopjuxw8aZaEhPU0Qeyk+fNAR5F+F/kHqBpB65C1TJppT7D0JVMyFgOxY9up6
CkwMeOr/zUGU0EnkTAXlAqTqglmKGA5crSz++fSr4Tq3v8GINjv2FfUYwut7KYwQA6XayuTMo0k4
aAbJGZh/Io0eJoszLbh2zT438OdxX8iQ+JFLaAaksTnCWpTRDD2MN1RpHHadm9PtKDENUfXd0VLO
2Q73tkcPjsWN8but4s74n94gSRdfC/jcGiwm2JYJ+gQeZS/JrdlYLqMx99koM6SDvVnGey8ZIQMc
Uug/WJ0RxF6n1VGK47mxXU22/tB9B8nvfjbajnEH5W4ecvndobltGiS2Ahan3haSeVgAZk58bjeR
g5SBZLgEe4P2Fe4t74QPNSWthaTQgHRP2W9wHMN/00vXUJXHcOqyT7SFl3pVgwLC0IM9hQ0Paoky
R6irdXQ1fF1YCfF9sjicdG+IVRhSBD7hsF1WyP6Hr9bADbhmWltkvchtytb06ZT5COC1iSimXCXI
8u9jwrgxOzNs8qiSsNU390l9A+I3XikFx0EiZDKDv60U4A0pw3DHvML5TXguvlVg9gWA5Yoci167
usGFNSsGsq/Pr5hlX2cO41ROXY0F3K12WbK8HTGN58LgUFgITg9KyLdp/iLYWZVdyZXU/4DTEGht
vuIx6RXjEahkg5Wn0dij34K7gQl+5qyUmy6ah48lXVHL/wQCH7aBxZjutl6HO1HulwFSVToa150l
GvPMr00x5NjFsLeBTyc57p5yriVUW9b4anByFI4krhn0j2JnMmZLX5cgTlW82AZnA7vWiM/UJMfO
Yzsc3PhmXDbwI8bFObn4MRa4XF1bYkSHtfuSg/EILOoVvMiA+bf7ZJwzlI/HwUZi7j8RvmG0i4K1
O9tPgxsFjoi1TU3+XzfxlZ3NjsfdfsMB3YtpKb9uHL97LZiAPGpa7j7fmePAYJSp0MbZodSU+CJl
3TFlMz5dlZ0Ibd29uua5qDuktOzwB0i95IyL3pvZA7hUsHOERKiz7PUAgheKjRHKyH0gPPd4C2P7
9KluU4UK/d6+nwOglbta70SoolUzfJORtDmaMdehQj+pfmba/M42V8UqVTBCiWX5TjhUeywjae2o
Rrjuglkn6jY73HF+Sg+DnFh8PikfU8+XvU/NKs47rV9WQcCMkKTXHQopfdYFMg1Ms/uI12ONwbfr
jTwYylxMl3uyTADNcyRapTw+BhZhD31fVH5FzozUQXsdDgYFlT0IhMl1trb4fjRVjass7eCeZY/s
rtKIq/fgNjcYRZKNxX1AtVH8N/02llMCLfeR0uLTi5xHYHDb3hebyxN5kkGRXGd5VccKvTIMGT3O
5RAoy34Q8cpfIPWxFe1rv9Gz+9VC8840mDlzm4mVVgeUB4q/2YSTHm4XTYhrfcWTnUJMm1LcqdhF
idhLf/tSAs5lvNfk+Kbpr0x5FghBe1nAnlqqZVV3KaTKbcsU3k+d7RX4w8+9phql6nqu0/vQAPtN
OIDX6zyXjTfZy1Wc1fBw6bORnOZ92qIqQ9txcoRxkCZsjavpmp4IQtuM66MtSnX5eRPrLDKb5lem
fFJa+dJYZ8k8j8Opd7Dkeruc2l2KGqx78Bp9vwPj1tiTj0k9ssckPNC8Yex1qVpB8eqKw0aTnxQW
ymUpf2EcJ5YQmsZyBB8O97692OkczvPnfehN+0y48NjJXEsGeXW7gSnfhscKR5t5cfzG++jeOdoy
i8i12R7RXvvFn36b2YW9oaxnF7iHdtSQtmSiL1rcPcXZ7L0f9e31/4s5ZHt0NUX0xgHk5hyMhsOV
KEM+46NNnGcFqLJPne4wr0ugFBi4YqwTrA1s0wmjxB5WXddj5W4yTuiuUv01KaeXdwWecRzSoCzh
D4XrZL1L1D61Fh4byPJvpV+frn9tauYYcZLIV19A9c2hBGY3PKYcPLbkX73mFGLmMhhZNYb5k8MV
L4ATd7FaqNky8M8ApeyMaoE2srRSOJWO5H/u9ugAtyUnxQY5dqGu0ZTMhom4j1Nl5KzxmxplVIxm
xVop/24lV/NgZaZ5WGe5fcUiFIckAB3aD65h7Ntv1AS80k3zaCpEGH9CpEwvyWoLOfkgf8XOf5T9
QNxV6ssujnSXd0hfCj89oi4FcXbUsNsvY7YjEGbDVg8XDyAMx35CUSfklEe35TP7+AW+mJ+s53r8
T268MFS/hFIH76SOiMXYEZo4cxjuClqMcCpu2cLb3Fxz27iWGLkwPIStbYR2QGnpbNbJ/B6txzbv
kuFocUtVcFDmb8kMDTSoCs1jJkcggRykkp+p90v0fU5zC4rccpsZ99TTubdid7UqM+OttYFmdCGf
mN0yGYuMC8EQhvUNq2coQgLVjRfztBRbj2FshDLZyfgFI885FuAz6wu5dpVqVOyuLfeqLX///se3
udBwGPD1mGtMFlL3yAx/ND/4nmrwtevpBBwAW5OS66fuTw/qLNELvMKnv4JYcpdKpmgAchcMpELA
6ui7UXp2iAehKKHGyuGB4+hTi9KWGwQjhFxdf4ZaTRv3vLnGTniNw95ZrW39LmmBnk22S4+Fgvrq
RcSSS23BWwP86gAd/a6kJWesD23OUk+oN5dKoDpMnfgHen2mVgOSwreFi2wifkn5l91UvIED1o1M
aReZHMP2qLmULprsWqg7uuJXzdBVmZcUaNGx1hDU5Z0POyhFlX1X8sEe+jYsYYUIriHG9C8DdFi0
JVBERv9rWNxSxpQbnLtVl3mQKfW7T2cR2M2XzlbPyf35k4VfagnVd6QZ72FW3f8msj29i0usCHce
sHltoSqNVH9XXgwSRzS4d85g0WV3AZzDq+SJjWqoVUM/4q0+cG455vkUesYocSTZqr7TzVQV4zjO
TAkaMNspFU+b/8Ha3abz1r2S9z6v9kgJXQTiyPPiBvR98pZlokdYiCFic3ES5eqqVBubnDfi+Dj/
ffH5rPfVkEicAZFXQHc64sYES2SWobsXszoPLan6b1nqQ/0tZJws23JTI0n+yw8Ytj2nSlIpU/bP
XuY/aZNCfQgKSVA0Gbc0khSo/q4Cgj/cgyW4hHvB+fnoVc9E7FxPKss+jJh+KGvxWl4gcSvE+j/Y
ATSxdXUWD1b+vHcJY5wyVh4VsspR5A8Q6YJXEANsi3fujC2FpBfT8ORDbfqOphPEedU//IPj4aqj
InZpkJEJ680sGs/qcyziiTFiBGvIVIQ/p2YiD8inQhpWftQXunSAKdZAU12qA13WIf/w/Uw11qI3
18w73jhapLqvTI2iyEUTFQBM45zCBWTkL4aEt564kjYJp0oMLOe0Ui/NHohg5tA2gYU6jbZeVNrb
LmRHQMxVbZmdC62yLYqF/fIp4gDm5Cbi/yeGhtDq7+jbVElcbnXezRObeQ3Q5F0tni5JD8YzpRIG
en2b+gkCJ7ThuVgHPCQ6js/BmkTwANM9SatgugDX4ZrRXsYIeGhfIAiLo23CrGk3ckgf9LPl2DsI
c3eOyfUn9+MSbZ9F0wQG9tAq0I2JLljrns5zqvPNgGdxM9AvHe4aTB7wKTSfdhkie1QHFrs77Lbn
6D28fnapBt8kqNPKGkUarP5y33GB5jUrCjxRVZI/2sGvqHOX5OKOrSGJdYNb/SYRyz5aI+A77uDD
peG6XIjv2ubvEP9aCFECA+GCONmBPirP7rnBfRqVqXaB447KyKOLB5GycLR6cng9uqGGGqyiw8tI
JJfqTlq5cPsN4DYNYPkWrJAreFPciNLtrINfL4qcseZpqCp9c6c/mUi7LzaIKv/Dt8hMucrF6N/q
yvNDRZonNnvc4dqTRfA6abq0L+FQpQtrBsxSQ+mjhBypuIvjQBFK02bBJEY6Rx6+/4L2xZBSFBxo
7/YScrasBs5NuUhtM/9SlOWQHIyvs4mvO5lxOJGfLGmQf5+equnxeotbsgY5Ex9Av/tpGDhtxtKZ
1vtAx85VSw8BgIV/+3oABqvQ4DNEnAa1KhXIfLg5NpsCvYlm9VOobYZsFICxNqOLjRtWl3XGxblg
j+PsWBu6Sfzmawwyt0KuE+szTsVV9J20NhZVSyBf4rF5sEPsP2d5x0RBrOISNIjmapxYyQ45qHrs
1XVM5JZn9r93kzx9cKUHxoHIbjNL2ao9wcz/eGhpUPSh6tcZCCqbY527bydaxk2J7RqzmdsxWHtd
soCaYcUGPayP68bDiaxI8GbyF7ox1nxbh/iosH54bDiUd9qgtMqlmgVo+Zi36Qu97d+iPlAMNt8b
kk7TrT0LngazjFjotIaGYzWh/TrLaGNVDD3jJ4D750nOwdfFrBqtUL82Myi7zWvkH07y29bPM4nQ
GN5uQy/QFse5YYNKfVm4cOnLG761D0GRZ4Gm4mHtpEJc/pOCxvOdxmEyQgl+jTxmXB++2KmBD+6X
L8R8QRhTk9KB9ENjyeMp66DtbDc4YiOI/pzsutGC334jyE1mxGetJRglNGrc7yuxG6lpQPHyjFj4
1s7MobE31xAsVom8r3oVaRmEYAzaOcvkgJnBq6+ygDuuPBmL94v5MsNRgf9acOekQ0lfT4KiXipY
k2YdBPgJ8pqriRl5l2mmd5nNHZtjt0HdQ06SmO7Cm9GA/7feDVRVhepcxc1LSnV141nNvh+Y9gBV
S3O8j1amaE9mNqWtOUplOuoVoCPHqI/c6szbdEAYa7SEJ+shvpbG4hwvGTAyKT71datI8t0kOGFh
SiIhZhs1xnUI8JtpqdHoTvvpk3BWjRPzZb81Hh9LtIjBKPFm9MM8v4+1hPVLfpdEV4P3bLOPEYl9
iKzvCFYHdJTMVeeBKgEDK2E1DTXy2/AyLtOFosiAeFq/MS+ib4LHaNxkE1WWgWCj8Wfvtbcv2dse
DcfSLrcI/I0sR+skwNrQq9Ap7oPcW8qUQOjVIrxDutDvbelH/oogqCbXGMgATt/saxAkeIFmF+r4
6tYN1JF3dMGvsYjZT5VA6h9nbFtRSFrIH+Ct3Na0C8sEuaDg0Uapj6VAuDnmXTn28uPmbl1T1u00
4G0J8nTd1RW5AvdolpGeq1khfNUmZOrXiSEG+D2gF8XsKZq3pvjCmrCQ6bzIcQEO5FEoBPb8+K5V
YLWaLkSg8uwDhGFPod1MJoqnHOAAhFgsehNkVkk3Gpej84+yV/RWzy0+GYGsZT8eP4iY2lKl1w/5
CAJRozGl2jmoq60uN49MzOh2WujZneBO3guY2pzQKzaY/VyALk3ofxb0SZp+aCz+VRS0B1akH5a3
nFWXUSNq9+sNL6RJLx1zwvi4us87dPEjtF4vr58xOP6NAbQHfw1Vs3NcJJJNYlT0sT/NZu3aPWDm
vdZORzGDuFRNWmd9IY3mOoVZzfjDwZf6InHwgD9bqZX/4CJAg7Z1Hu65cajEifVqfFbMd574MU4f
uxgXH1PFPR18NyatoI+gbzbHHsDzJNCcJAH0rt06jKT8h+DF2d2eQuNUxGiOp171DHYALpxWYnLn
SuBShVYMQ/bpX8LRI9G6vngQhdOpcqlOdz4WvLPJLtckaBNUc+HUiUlO1xIQv3zSUUeI/zfmJecQ
86HqfYhkwg7beh++luh0INZsQvNAWZJaaWLv1HZkMRQCM2rjmiIeJDE56axlP67MGiRhN3nVo0vE
lX8J/CSgVBJRhcE9i/Bdp6EmIG9NLkqdx1slV2xGur56X50vFpTLYByGur4R+7004rRvwCcjAJWX
8PY2fajNsjS3cWTmSOwwu/dN+e91yVFSE9/EVMaZj9pNBdHq7D8ahCPuom5y3r3AQRk3Lb6VV6fI
iFunmn9sp2Mf12JNypcj9mry4WqGWOoqE+M3vPh0f8CilQiuLNfQjE2FE6cvZk+G13ifctv2tkf5
S6g8+dBFl/CsmLoSVXRFsRfKRqZZpx1qGWlW7roKyE5fw6xFoSQRaWjuhYEAK8FCeoUlHWTjNalt
2Tuoqp3pE0h/toio6dAwYl5+cuWkO6+0n/AdYExiLeDz6yf2/ucSXH1o1LgxuDox4OQfDEWoqVjI
CJ3/EWzwfrDjEobsICZ75V0ZyU4JgY+UhmjFaO0ysgEf0Soiq2hjxTxoi29QjN0cMus4B00tNz7e
+9rx4PqunhrmAM0c1eWRdwLqM7E28M+FCM5rcK2gFyKSa6NwVzylMMAzMjrRjw+sW+iCQmm0lvbO
OJ7/zIQ1lgMzRCoASiDQmBaZIfcgeIFNU55Pt6e9WkGCDBBTeeVOTahZjR+MvNLUJrVkyUh3XCXh
oxU7DihW5yhbkVfiQ+Y4TP1ZagZHYV0HuW1W8yOANRKW5fycLd3P7Z729+a5UK9GdCHYBvzsES9/
aQRjkFCJx5sFlw6+7nlOy+PU/bSr9fnw972x1SmkzblZ/eO5ns6ir8iKDniGaAuUdFhz6a5L1CUq
w8b81B33iWZ9DSW9T7yaukJiBwXSZyGyDgapTGHfnxFYHe9KokJxfG2zhKlXPOaYinHuTZlwpSZS
KyBa7Yfivi7gkrA1u+oWuJuwuB7oEp7g+qvU66GAJmJwcS+GpjSXMSaE77+Zu3wm3QPw7If7Hqfq
q6oWdCALmL1r4LEuJpvhZfKixk2ZIgjpoT8YCOIjvywkGb67MEw7w6pL+hkgsv1TXA6HjO1Ir5wE
9/Trt0WsDcfu0KAP5mG+2m5dNdjcNt9FbQTpE+S8JbGNLihkCKa2I9oDFI6NBXlsnAxov1hHIsD9
DSr5LYeo/aYhQ0ohe+6P9Pi0Ms81pFrtClk+KqvAzPEJpk6X3QQDrsQDU0qjzTXZU9cKKTBxEYqW
vjjoEcOH276uc+L8YxuPuo8xHulXWScbQnhnSPsf00wYrfsW3KwTgBPKgy/EIpAWkqyNdJQhMPTr
OEv0y0ImhOsFdTr+JbpQiC4gg5NOXVILg6F6B3iz2FIh57Sj54jU5Nd0O5ZxBY/oVBEcvpVkeC20
1gm/SBjT9eOY1QhO2OkvHEZ/yE5qzMcWg3p4OKySR2Da9F58V+e55wAkbT3jx8u32rwdKyrlPowA
eD/DkNFNhlYOsDfUh4nPAPsXcdacY7ATOdzWCz1YPcghpqzIbKQ3IlbkQGcnANSMFBrJ2U0YayIb
9gz2emzbPbBhcUEtdEpdoULlF5Yrl5Foku+JxqsurOigU2LfaN6g4UuuQjJLVF7AbAsWxKPW0y9b
jFRBhlav0Zoo7y4MQi4pCKt6/AiO57y4ooMP8sdjpML/JKfRHgaJFy84BhSBV+jLxYp24jXdEJRt
Q28vXPEL55xWc9iRQ4zcipF5LVMt6K8RA6Bp1d9T3ijcq/Zo8oNkM/t25LSltxskmk5UfkfizERF
drdYCAflX8eWr2dy9olAKBK89duW7WYC1Fj5p4sn8nrWLT0jpYWNJH/3VSPMEWIACO6deiQH3HU0
3jO7Qybi3+9MgwmbIkufwBXOwvtM4tqiZcIYNbt1NSyx78G2DXOBl13ZzwOFUYZFuN0tktsm1cip
jotdECaEP9TWDmlvqx+i1rFAY5FFCiIWGomEiSnaJWWWUGf5OXNOm338hFzxcfpytd95S0dfdov1
g9WX+H5lrwuKwBW0qqq+VO3DDWY2kh2KvPcnDtXn4I1zci8R59DqIXwB4tKkBxWQRDgnA+K2zq4W
5FDiwkBxmfPMt8USYoaTnkY55MiSAu1dc5s3cTuSk6kBCEK9v3PjzxKDanpliECP773QiA+E6rOk
WMH5WpzcQWBL4lODQArfwJ6w6tK4IX9WSrEmPLBCOuxtu2n8BdEtDWw9U9MdIApYlbW5tU1xN8fq
RG3P7xt1qq1vkUxRXTf5ywL8MvPJPK+YjjOT5Kbm6uxHgb5dxyVVjiwJsh/Kyj13YrtotorKeL1h
CMQokYE5IaErCngvBjra+/qeUqd1/O4sNjO1Lv+J0EIAqi3/VYk1G5z/1Yf0uz8ZwPUcqzQiWMU6
Kel0j4ORnohRnxEMzGOYF4l+FHIV9xAJH+orBSioiNLc0a0Xp5HUZEkV4Gr+9a/UNrvFMrdegShM
WCBor9oIsDeBU1OIGy5GBvVbkJW2bOxheRxbHInVIhAdQrfMXmAUt+vCmaHNALHv/TTVs3uuP6D4
F2irnDxakD2l6SiI2UbVE25x9l64P8OsKIMBGLCHY2+sm8zM4iBClrdhZNqXGl6bqA43AVOcx8l8
CZrTTZaoMXlcxp5lRKhXzkxPYFu3bolK6aeoP4XL534DFbXA2JeI43MN0OPh/9X3W5pfD6iByXFT
VPPbZcR9QkthqCK5BC908v+3TqVGBOOW0P2tdSa4wWOngJ2D7lRaULzw9rllmp74yHd6xXQFKmCK
v4+nB+SSgxVeSnFZRVavd/66WiNzQ9/gLunjtega/M7QYOeGlrF0kRlCB7gWN8xV7/bCZHWKoT3f
GYGC3ckV4llydxjvX96Ua7f/6gZxRUHIuvpC89aYxUYNYuADweD3TzWwcQhy1czVrReMO0O/rbUA
cDRm4GDe2oeQ0ePkg9Ul8J9DT3HRGwm2Jq2xjHWI5HudlyIDCc3yPPF0AQuTcVJYkdEQd/8cNmcI
RhM0goBhBrOcl2VGiYJo2btAyuf1PRJ/iXtRCoMfrOYi2+2uAXZI+0og5WecHmiD5RIPL7V9wdeG
9/4Vyd6ZSvhoMxca77qLMvTOXn3IZxr9By69J2waIQVne37qub3yKkVL1JbXU+l70aTvyz2yUYYn
J3K/fWKe1fALRnD9orGrPPHGga3UlJ7yo74RfiMlArX7c0oBtcGXtgg3EFQcG5mZSEsGQ6tcUzpj
+KJCYBzbQK9Z+g8SOl8w6vJ/pQc5gbaMs7WE5aEBuePtXggRVGL0qktiGezIyth3bWZPydQ0Uy/w
597JyjbRacqlgAoK6o7A/CyPb1NIjpsn660VRhYJMqrcbWdVhJCFM+Jw025eq7vE4feuDYYR0itk
Ua604SnWEErf0ZxrXLRaNQusD4krrhUJVKq/w6CCs+XS+i0/OVNIhBP+QDfmiHAz0k3czWplPh7W
IFbQO1YOd3DvoMtmBMm2gc0gop/ihT/sdSVcMfmaWbH/4sz05bTHj7g9h4HIsgSicMxoSDZ0qTCa
xOD8nL6g07lVTVEo1suSd7skyPRv0IkSLPYparMjyvHDHqhEDXdonmMo8q7PVI1FsHgvTTcTdDAK
GaznpTsMX7bYwh76B9LiHG9qSW/PGVMFaDNG4lWR6ip91l6L9W/LV13QKLm7RDn1PoqFUiaSkWC1
KSnE8KQ70L0ORuXcQ+8eiQ8MVX+vaJQppcUToUgnURpVUORr+dDKRYlp5ibUW16VrUiiW8w/1xRB
suWpbZ+h94H9MhsWNs0X6VI/foxvS0JQIEgvG5M+R1pYt74vLLGBz+Keq0g7OgfNplVe2q4uoEvN
WJcwfUj/sn/sn82LHUCIECfPACivFHQb4m9XZMRt0/5UK7w5QNvp1YaDRkCL/VlfzyFPT6iX3+7l
5x6ieRFGvatJ494whpqNihvz9TAGjgYlDM4TBo4EB9wtMx9Xdr0hVmq40gz3K0+DRRoWNglTpy4C
7wcq1jFZKheDON60H2ueEYycWIQK0NpJUDCw5zz4Z32Nc7FeE6sj7oahh3GvPC+zl6KKClq9DfgZ
ZNNkR43dySwbgeBlhK1QG7VBVgpGe+xy7XflVJhohQx+0OMuSSojym3GbUuuOlr+knzvizsF7gD2
8Ve75aNAq//xRXCDoc5h8reUskGLAVsA/NuYF+oAkX8zbYYEAwVnL7VBuSgBnNc+zQvJYu8LXyVg
aPhsJWluztik5T4CDRj2B2oNaKSJFXK/qeC0RPvQ+RsrZOSeVyvZXRk6LOhSaHIRbZlmo8PNQpAg
/Kn0VPufGpgutO9K9gvnj08PosC2xeGtl7vu6AOso+qvIz0Q438T2asae8nJvmwBPHtHnHZG4n2o
AqA5OvSMVp0isbfbAEwmKAs2vbo+59QoMZpXSG9EIOMFmlRZ6CEVUF5w1tedzIt2BqhMl5/JCfoU
yKVN0eInFQbcyNd+pzmgAK8B4dHeAdRSeHyQ6R1B05lw6hEBqFeDQoDDHlSKsJnVaMXSVbzPv/uQ
OE54pON8t02Ke2IKTHQ+O52RbcNx/8lTP+7KsNFOolNLvaLHQkM3IPdecoiEUufKPttsLISBwV7u
DysBQ51HEyfCcg+QpPT5gVPES574EudkULTJ9RYWSIP3SihECVvcVQEWdTMjGJ+/hBI6U9XUfotm
DOmnc3RH3u6Nwoueo+Indoz8FP5s9ME6NxR9/6seVoprRtOxKhYASeD1jsVDIEpmgi4HpkHBYSDD
3ST3GI0kIp5HLplwd3Lw7bWjmPrew1HqsQ/oWU5LWgPUj21vXmFDZPE0YEVCIgVF6TcZEdtd1Juv
ssXqRE6R9ZHGOQrksf1BEvZ6PQIv4htYiEdehUKkWMtf1LuviELKnpHNLnyqzhfoRxii6I4px+aL
p0wgQmDkdCgK796fOBvap7/HgyC6oyyjkynYMPaNgyWbmYE8v/9clRehNhdr6wWsfLaTMBVXKtUM
omV3UeGS2FBa1CVZ+HjxJq1XHAfpd9sCrBdxIpvjscOgy/17YsTUhJlkLdhEbP8BaUmKPlrVetlW
Q9lK8Uru5jTj3oQSSh5j5gUgUTotYZ7Urqn9tMcHNfaDK1+w/VcvGLKZsfNfq09ovVHcg5krpmhb
4tWVLHVroW3vKT0srEfME4uEceiSGjqOLnwTMZGTIOjGyq67913v0q4Vber2VbH7M0Pt8Y6jb+DS
1BLf2xEHQ/tBe91zbh8joeZzXQnzsZ2bWYop4prNkjetcB28tYsrDfw65P2rYWjiB/1O0scFTZDR
zGFlAZjP/PZFezmwRTVDDmrABPKdy7RRKAUVT8JWkVUX18No1qU1r89zeFGMms+fKjxsq2PxcmJm
pltFe8qCSkGba8OSc9HXVC5hCLy2IwF9FmcUxHD8zTjWqrJyeBkAKdGIXMjuhZssqkNd2Z/Y4ovV
IQ0hByCJVkmFB676FITeyFbc4HnK3AUd0YT27711+ZnwyYduTJwly8I/iknNvRL730PiJKtOqo54
rI4SYRL4itO7DWHHf2tNlMKyaBluIKSJfb9WaSP8eKp8KCx1VG/vpXtei1mlU6J+zYBd1g/dwKSK
VXvYM6P7BlNmLgqaDXPJehImdBfv3fzEMnIp0MNLmAJl7j0O591tj3qdolbWjwfKmphq0oYBp97e
/vkqcouRoOtcMzJCg22yAnunm3qcllFFmUqYeFjA5uhI228HQENCx4ZZoIyZgYvf1wVils9oow2S
j1fZL+kIx2E5d3XxjaOdfUdzMS0WcV2YsW8GmGNMq02lNvSDG/8NB+WcSEsgE8+Aesre13JcQNTy
mietQu1xz4ABLaPQRsxtQQcHIK2+vElSBQelEyOTWDpl/7cyczDRSvuvu1i3OMvaMXiFBu78B+I9
G68UoYn8aQeFrJYFmxziEzScFW4cjzxC3MP4S+ZuTit+neWXGXTlrriAWX7YiWYDb5pVCPg5KIzy
qxdaZ+wQKEc6c7wFjx8E8Vgj51itX/FyI6inJqjlDkVURcQg5vQHd2MrWMCVdJjE3RikN6vcY+d7
93HQjAaBtX4L5qaBkMVAwpXCIrKL1n93FO7h/mjFOcR6s28ZOb62pTDm+YQJbrvbjwgRdv79P7J9
gUjYhJnV212ysOC2+9STFyhqc3BS7bSJBnQaa9Cs+ss4ICVU7EToqvr+fiEh0y3vPK4L9RQyAZZ8
a4ToohoB93FzNj5CE9hQ2NnW8429Fz4/O0f6MZCQcMxZRqz54Oloi9au2AcXkJrWMfSmmrmsWsaX
XWvP9bIqctnSRdb2eNoJflsLC/LZJA8JIF3qOiN09kNyM/ls0Mcg8w3PiMBikMgmOKrxiSUoO2R3
RDTFdZ0TN4CmJ8SVLi35zFYC1/A4BlNyLNFZCTJRwuX31px89nbasY+HeaY4lKxEVr4pFluknIQI
2wgCue2AlsMMwmAL0EtGgyhU8/vU5/AIjuYlYK8DF+BaAw/a6XdfsX62Hy/52K/i4RrAkBwIEGo8
UgMbpBqkXTK5IWc67SwCQVeq+3whZ60q66zEntq7x7F5wdI7f4GyzWkOqGKMqCdNw7Y7iEyiQmto
NZ65Kstpu4uochWbCD3En9XabBTTQU90dg3w0d7M3r2NgZcraoIA/Jm7gp8VZVcLe5nDRtvKx3mV
wj+1mUu08wYCYxKNllwmAEoFu11d99t5Laosv/Js32KsAs1wFQwF1CHx6PGlfmieAVlIi/fb4QsQ
yjylPN9aJu1HmxrSd8mcIyp39jeGJ6CHaKnF5mYQrbt5UGQMFWr/fEIG0I4rKGD6D9WVGRJFyM6h
RybdaqwoRzho+v7LHcNcDU7XZR3vZ+C7Ei0nrOegGykQCCt/vijdwtWaLW3RYUb0taca43bWoNGS
D1ZbhYao7MGrjfA4pGcyqWwJ2zX7gQf5ivMoMzhAFAItr1e5HkWsnhnYpGO//mzaYpisKx5bbUNJ
99c35xmd2dCvhM/aiUW3l4jo2gS00b8VL7Ri+IPazHOG0cv2h2n8N2v6jwP6RuW27I04LZW3ngZo
oAhBnoW7T1nvLPtRfPKUaqx6k7v1EL33Oy83LtDWN4zAD2plWRn6wASGABinWRxhZAQOPNpL9X/E
KHaBmBGR59+a5WGnG++CPE+4my1sTnk91f10LJZ2clCkO4ykXJQa1SyuM7roQ0GHjObEmJ1A0HEL
y69cl/a4jx07H8ZEZLuSIIIA+jAnRyy086IP4N/Gmwp7erv1is0jWDx5fMbHzUGuqe75f+Jc9xLn
GevfM9aNkNhs/yJ74laACn5hwX+4eL/CBGjFugpth17A5ky1F99dkwcZ4kktVTdvoycVbzr6vfLC
Zp64j0Nyr+gUGfuSR6lNkz5RbCz6ePzIlMmKZspG5Ymr//PLMzaodLUVFYWTYguawOtwXKWJI3yF
3VOc+aECpiSQea/eY0tQk9l7kFUJip9cE3bw3v0Ozwpkv38mFPolLVDrYf54Vm8N+N7q5/SpSlpr
6VW/D9ymJrFEqiz8lcNm3kCYFAXO1OtUqk50yiBtocpPdmZ6V+7XwKTFxhu8WZG9YS+8yqsivdmJ
9BbiRB6RliWTNFSeVWrHcn8OOSaSxk9wSA4nhQm38AJbv5ofvI0CWgH/8Ua11W2Z33iczcKLeWtc
i7dQdH2HyP6Wr08XLp0J1tgv81DCYvolpT9FkvzKYSFAA49uBjysSdySj5alBJOIIxXvIeQBiGJ1
N2KFTuwnX2/ZMgLISco/ixsVwaJ0sYvYc9yBhlDooK906m7yg+90JokefeQykSNIQ3axuOyYcknC
pbukk4lfdzcvJD1gppDhzsELJjJlBVfi/+r4IBgaNs1xWXD+Q48RzfOryteCCJZ5CuvhwtTFSYBq
5AMXbltRBTbkICZAbtvRrpJERRfo9fhFNzlTvXE33CFYdjNLaNfRT6VG6pMLoyM4+wPpc3ZD86iv
twRZetYW0fHcFFYyD0PW30yAXcKwvmBXg1C24zK9JYWd6NDxvN+Gn3r22H7/1UwApFYrSO78Lsqg
gt7qitbVrNFpTucLbCWXn12mS5gvWL/Mys1wS8YmZuFG2QtAx7eeJ58hf9I9McaMG0PAQMCWwWa+
pm9t+en+9KnQGKjGLU52EtZGiVreCvkktmm1mwdAWqdaSGCGqTCUm5x3d8TpafoF1Zbp3Gx1+GqM
Tzayq+xI38F/OFmT/V+gaF9yd+Qym91/S9F3Mj7kQQWG5Ikb5chxVuKKqzDXH/aNmg5H7XV5NZDi
308bQ2gIMIIqrCz1mt06FBiaXpyWkBJ1QQtOkWEz/MOr97N00RnJQ3V6HBew3OkE+vEdHHPQ7B48
BLcJUEXJmg0zoDvevd0wLAKIulMDbMuC26NLDa4YzA/X/1zpf7T2pXv41lAb4+JV4SfohqrHj7h4
xwtAC6Jwdsu3cPNNMcRBh1HzdUsLsDjsHx3S3d7Zms2a/DCPNLBUqYsXrzbvsVUiHoCAIvP9HL4M
WcFQMcktayDJo8qiNbRgxL+c+GnvIbXnsoAa7TScBmIadCI5pVLfVTPIhBWs1SX3dLVi8rvegAFT
5NgCtyJPz1Wfb+AOzWCEjQOULP8t9RpwblExgkKR+jOq9DU9BEWJ9sFDjyZSpn+6nN57tSsqhHNp
OlnauZJbii2hop0P3REplB4fUQ/JUOhLtgwOWkSxvu8asurCR+bH9IIg7I01aoOGvs5bBnRwsqCy
I7bBqxGiJkck5jqga+flnW/zTM/izExhZ8+pZZxxh0UZWu7jhM2umeUGY4MA65qHarTI87w2PA/c
yCxpa8SEBOOrc/1h5nuK4auEkWQSkWeS/iNHqC26R2SN48Zu5q/BKaFUXGRtV4gHBNdCj8YUu61c
vzLKBy23H0bLNeYXG0JJtki1HjcgciyXDaOI/5yjZmNPlJ/yf2OA6k+AMtwQnc5QZ6wpCIXXJ2zj
HEMIZ9vD2Kmt2AfF2TFg2RNnl9zKLl8A8/SDEcqer+SRn4JGjIqyTt4vQ8aY+uaDEHAgjcDeGYxo
lzE7i3G5ABIW+8hvMDG6ufFjm1ggBGAhwZfWRJRwC4rxj9Xf+69WpPlnjiR70UYi6p4/n2jktPcV
QoQSw4OTUApQl1zze8OWej1Gr7nFZ1oJoapMPSJeHQpfNk0jOR0Q2V/EagX28uOhNZv6TqZAXtqn
u62NPbSuycvlLi1EvrNizpZxLtHP3b1+YhZkCcpAi9tEnzRfLrLVNEGBVd+rHtq1CfsRiz9kGRN/
SgndraNZXNp0FwYfJEnLHpJoO74uZERxpEXhxfPbWbOqcfTZjru8S9j6Y1F9htqvEdG7Z47VLVdh
PR485sfNut2sUU9a0CLeYONu0qZmyZ3+D7Yyxm7qZc+u607ClsuX3V/Fddea7N6/R6QphwhIQdtr
I6mWe1/7F2aFO5e2iGf54kuS4LkRgVcY2CZj5pQIWecsSHc3iH274AUtBZCPgV9hmNYrUcaLJYXf
P2esfhi0MqEbSchZ2Rz+IGlbrlN48abqey0D4ELTWVV5tAemloRffk7lc/z8U8xT9GTkf58KXXuV
C/rRSFBwawzWXpd+LjnML55G/x6h4l5UPX72FD2jV47uZ3ekZdr+hyvksEbpBpzRW2lQbm2WfqmN
24ZPHEPeTp/Gc0rRTBXwIh6qIZSGJOYORVbs4j/128a37HwuH+sFOS+FrIeA51EvrN96E1c/uSXq
aUUkYyweBg2ziKusNGyZIGmYkX1a+7FNKfalWdeh3CPZNCyMHGGPhMgoxOPwErv0y7hXo/27nbIY
TjWt8SwSq80XNH/hxHK8AorENbCxKtvHSuvr7p9G5xc92LamMrySvTnnJ4CuOSWNQ2ou2Z20H8aK
FsFQQIR7zxDiXk+tojC7vO8maJBGR88s8O5Qc/ezuvdNPJSctpCIEWz5sJUgz7ixQe82qRcLFJel
Cdd9sULx9jBJrrePsf13kZDN/nVYim7i4r1PDnZ+ND4RXnrvgIsDL2Y+MA6y2dq1OlQq3lsnKqer
SRyrhcuOAP1VW1misjKm2qYt6wUQmZPmM+C78RPikPXlHIiBInZ+zCxdqcsN6t+vSA63M32i65Ie
UOYidCOod5UywyGtBgp00YmprJV2cEg3aGn7tX0RrMBvn6zRfQrK/5Pk8PXVzx6AqMHkSymNWL4+
2sTKV8y2oeyMYwNFl2xnA4Ms/W8RZ7ijPZVnLbiNEzTKahkMlseg2x4aOw1FE44KkrMvVxASuGow
MEMKUnKmAgMjv+UCqFoYDzc/DvaR1kV2XN4fngzfNGZSFoCrGyFB0pasQa+3d6qBxDA4AfCFIcC2
EHj79eGjMP49kOLyl7gn07hmwSOHthW2QPcROirGu2mDGXf4N7WT6YhjhTlb4hh07ZyBNKWhjH/w
hqBl5frFwSatIS/DblW7qt6zX8XqMhx/AklRl+vtWXvUjLgf0kkXfIcTxI+P2/nYN5UTlr2GGHk6
V8kScDJgDSR87BsN29/ZNrUxFUbfpdUl6sbHUCmhQO2L1559SdFxYC/POY7yEAstIFBPORTUlPqe
qkSgMoZeWvU+NByeQ1Smm0Drxb2g1ILjTq66hrQsCxwtrC7Gggg+cguURMHmxJYRInce+sbON3hl
FDmR0IPHI1SaU2KBjKBylyKX364oE3Cb3al6TVVN5L+7fMi5GI0DWajhAD1HrQ9O9cTDM8UdUjrt
kjbg5QuoXIs8mCaEb63c6ydS5BuMsw0Ug/+A5iLCAEzK9xG3Wnd0XUUXV/Q3poL9frgh4iM3jOUV
SkSVHbRO3k1QAbEjYYC+ho4lDvygcSDOAXd1nOlRHADBSRvSHJCRaVFU4gMe0Xwo741bqHKFJdfw
NgJNKMsthR+Z6ZHPPfpMel/GUkorpnYEk/42yHb5JpqnmO3IIaodsa7q6/8Tw6mDXKQzHMfXLdGB
CwjPlCECgjjUI9TLYqJ1BtDm89UvJTxKmzHSCFeIPnDIj+hbLJ6yveiPqUdmTn376tIp+Ntq73GG
Elk2rdSXA7W2pAjrcR6u37lXwlAuzkWZ/BTBH1CDxQvDcIE/KthQciDhnKt05wZ4ovgPZjg/BplL
ViGdkpbcTjMO3St9fusTfAohdQItMoADyvAiX8bwh/cf40Lvux1F+o2swi2rqWcum4SM3sK0MqbM
fi/2eEs+vC7AtjhSE4soRnk/Aa+EalojRNWXG0vz9ctTuTE/3UDMj7f3lTjfcUtEl3gTB7PYzE1X
ocFFkniBFcb53Stf4yP5Cx7txuVzyfZd1WtKi/z6PYXJOQfecBalmb0utBhzlDcOvWTYK8dqn6NN
L5M8rVzd/gHuwhoWUNiOhwBnKc2eYdAt6JnGHZ9hM0LzKD+OTWfUezJ71CiaMEMz7+9rXKuxmdkQ
AkOPXvVc0506+4QePYrpflDo4x8L1co0bnxTzhxNsJKLtUs9AN4QuihCo+Ef5MT1jWN4HSjxNjXh
I+mSBh1yymclVDQBz6to1+pb322fVAvxGCzSoIIv8KmZTQAD0FuP0SKT8z822yZFjpf/WGePNMip
HPr+uFatCyZlJYHb+BUvSCMLpyuQV9WfATk93YOM2SdPqblRKEakAQpVoibP+fHFNVnG7F3IooUX
01bX/7jruIyvh6IKe27vJdWN9sjXI4S7RqyTsgb9sbQCjwnkaUCdelRbUlepGA/3g/proiEuUpUr
kcmgnU+9ojx3C/YqMXqf1NYFEQR5RCpmdGC1Rp8840wI30TY+9hzbL7Ra841Y6MR8XNCz+UP2fDt
/fNzd0cqw6RdtvMbFSBOMxRQzLc16F1UdgRtJ1MB+Ks2XSH+IzaXaA1IBhXb17DIKdEsmGMe7ZUU
USj/pCO6ogbI0AmxCzhK95xQs0iVwlObKDZrFTnabZiUjAWzgPuCkTQM9AK3Sn088UZ9CpTuzpAr
bPxA5Jml3IMk9EuSJqROlz1zHgT6Z2kIYGfOKxRyd3r4ctnOa/MD1wYt6OyNicnOawTbQ0eDmOGB
oql9YUipDMeHzCbWYBbA+AMVCN+EElGoH1egR2EzKBkXqqMlgyQT/zxqptKKPtydO5WkhBISWxzZ
oGFprNCIRzEgfuP6xTi9jUcBkpYQGLf5r+FaihyCa5csneicNGFBdr3V1y04soyH6+WZlToL0kLK
P7ZJ6UIGavsD5fACo0XLh+fuNV3yPiIvKAVg9UQwQWgb+MnI5Cc3ZnCTehqv5oWdM7lxwwD+8TEQ
iXJJavXIadOOYdAnao81/88LAyV85mczJIYem9CZEnhCJJpJXZ2HbklK3b2v/OJO3tfAV7JJ0qvk
8KhCEa/0BrIn2ehJkF6kWyptBKPQchSwrw3382GiNOTH4u7rypFV0KRsp57slhwnPQdm6KXqM80b
fagkWQDeJlcWfyIwQXMFb3iLTOSimKyvMGGp1xgu0h0IOIR7vzHpqpTx+WBmjEe8cYmEEL35wHMS
Fl9ZA3zkT86Dd8NlucWHJBYKoXwyO+vg81H5JnzT3qleV2GtImEJdLrMjsA635wStbGCv9/dOxv9
232UiqU9iyHWdYgIwka9kzZi1KF+ZODzVsQgMBx5CxiQtgfM8+GxBVuUxHY8PeGkuDS3rrb29Njs
9oieVZ10aQQ6PHlWgaJ23obpo89bjUi2LA+5GI9XMmdApjSxKZmQde+Tu6zQCSTghTTB5THKh87m
iK+fJEThtvo5KLXoWSdFUHP45GPt9a0JcUMDsuhZ6ABTZvc+cGYzEt+bDROjJ2ASQ7NDxuDOtHty
LTjq7d7WTnZ0+yAtww+7hfeUw8PJn1T7tvSGgRIV7ET8PQn0BCKfz+AxfOmgWKDa1mAcWJrZsINp
S9ySSwnRPTs1diWjqXdBhUKvolzgqLElSKHO2RLCSHI729qg1RqOZ/vvTOP0gAoDr2wor7ZHkOa5
7+1waoR+WKOmRh1seZ9L/hyhN7wDoh5VXz2+1QFozzZoEOAGwjsH625eilAbQLvsvG40EFi/cWsJ
GxTWT19/E6HThDFx3CaGkO2vRunmcZEG/NZeEr2JPkhjsfz774vqG7wzzG9f/pZKS5TMDx8zTqmc
+//11J9ITkJXd+JhPb5+ASOdwqta8HJT7/OMSC1lvRKeR3xNmQKJnqF6dTwCy3E6IMYrSa0KXjF+
K0zdxLw+UH3GiJmm5moNnDiL/+AcuCWuKoMtbHtAOyZtu8+EEpozlb5Hjv1H9Tn7q74T64MMXM2r
dmmPL+BaseuaVvfmwY62ZEHI8lUcbMIKWb0T2+obq1MvEEIKxkY5lSdcNY+3QVpZFr3VMKWeg56e
jaLAil2KrIegJsAG5t7RvnxoWyCsR8oeVAbdIHcJUbwpSw9/+KhMKLw7Um3wsyTGTJRvKvujItpy
tR4IYKENJ48+tnSQL6YsBpCnA7UBZJ6ZVDhIOrBlAotZgmWHIP5csbS6AyWJbp1NtALE/75IWKV5
KA3x593Za5Mj+J4FVo+cwvnMbJdhicVR/ywH5s7WHZAUq1OkIZCSEs1HBgidV/imwyPWm0GdGlN2
oLggly75IjWoTk0cBHn7vWNGD2UTt9K/1Xwr0ICkNc+qbY0pjvx4VVwY8XZ3p5WHjRei79pRB5Xi
1Fk4Om/UpvKeq7/LTz0/9g21fNjRh6cuy3i98ewi3YYiTSLX2LGPmX/JB4q1XDFKuf/rYcnlHgwD
OKjUYf/jWkI8QIJP9/rYmAQxiSxwWTghTrFvENi5vPFk85sHRWkI7sfbM/6Do7TeXRIPs/F8A+qQ
E1nArPc1MHubiV8AbrAMwspiAVYdnYJPx/wOIUxIMPfvYJQJJME08EGzrw9u7dXaGWiU5uEJrVPU
+vfKsrgUg/Z3Hfa8ab2lmqtrlQ0R+kH6c9uA5LRnPbruBAxYwtxVTLK9SK2ZtKuMSGLktoXf+4ka
W4eoJGHu2Kegl0kTsr9VSfjr/j3po9t8BXpTPXxFAnWjvvNBKgWxbS+DO/cZNE9CA9wEfP4+J9lE
m137QmG85MpOxQwXYdVt1JycY12PecAa1Tl+42bV59i41COKk4MW8+8bYyzge0FcljXXbsZ55HWE
vHgEEqQkYb9gOKMjYDGWb21AihipUfrbORH2slHAeq5YHE2oNG/2nPG2Ss+On9QG8fPuTW3hEDI1
vl9d77NhCLGd3TpTtJwfLXMnZ7ThTXGqm3DddARcygv+XLOPvZFkOh2VEMQoBLNNFdLmNXVlnqdJ
05xsssUkQ2VuUH+iJropLiNQgxIpVK7jxW9o1lf6PWY+YOtpCMJosDVnYLcP1a0RTNVL38Pw/wZw
4uSbwVt2Se7norayFuscpa7gZ16dlIyS+i6SDeS1foFrR6nV771Vzfz2iMmv2v25xlolGD8rqvtU
n+uhtpDB4h71CUe4pL+1YW+3RMf/SNINfhnWeoxZZ5FlpfBKCklay1mXmgL/kgzWd8hKt539OSOu
YPXrkVwOf/I7TOWnpx10F0kLi8AraOYPQX8g9/Tnoh6yDenFp9GCG6x7kgv0bh/jj6njLq1AiTjy
Y0x6luo/+u8rYalomkGEgd5Cx75TGdJ7f1Gz5rNAjhlB+F+jpJO4fXtzSB68YhwqKDji4T1TH0GY
WfDh/WZldmIka/YC3u9VWpKmSAstf8Ljo+vuImRm7F5A27fsJXL8UuWbpAdHnaJEN6WOyu/R8mR0
lzwan3zBbdE2pTCZqOYZ70pk9Gcq8HfXLq9DwxZeCXaBJIFt2oLsLcx9WScmspzHKDg5XiK83286
f3UPFswdg2gzduPUw3KD1P5TFEpsbeFH50LWjfWJogTtCBE3b5/Jo5Z89Q7oHaDdVb1X5fOUfhcw
FmlI/VbBFBbDpYPvoHLmrLKSj8wm6IaKra+mvPOwkEg0qLjWRIcd+ex8qhJxsiWlXDLASNssG1bX
be0V8YI5kPu6v7EMRJQb16vHNSxK3cfWPzNz9xwB41qIiCDmwxtZGQmtMqEMgaAJk4vIpCIVAkoQ
BdjoFoZKDUwN4I0OIGRw2sH6V9awdCYQPL/Tok3J/STXsXlR5rJaF63QX/XKc7ZFMnJYztYDPCy2
Sz4R5918CeaUzI3OHL4pTkNd2wAupROlwP6w3ULrjUkcTbNNsDWKZZjREN8+7yHHF8ABqvhJXNbq
mBNCB5Yg7hcoGJQu2tbYkZJBYSgEfoIPXLRUF91Xvulhm5D0hcbl8Vav4vaABDwwvQTvS4fqm9Se
CP9W0hL3xzteHHATKMf8axKS2QU4bMb0lQHmT5bWox6xYUvGtXPwaRWMpxKN/N/cVdLAQiS9KQkD
zUl0g4Q8+RQPYy5VdyPHbqVd/y74LKeoUBAwE4pKA5cyA+JbkM9NlkzXscbf6KvxCosFxiF1mU0g
TuoI3qwJYMPOJef0EqC8pBdLgKpRfqn6/xQcw0AoX5k5x+5PBvngxQN1wrrFlUaHXQp6uc4kj/im
qLIO1xNrvpnEpRx9mPS0jxrWc4/Ddb43xfrRcEHtS/3JZDKoPO9PvksiAx7Y+Vgs7+S6Y+YAytZ2
9DGaZA5Tl/O3XrGlWdNnDFuBIEsR73vjge7KPGb1bYo8pKP1iaitW3aJj2eMnK4BiN4HFJ0XMF6W
f0VoukQCUYzeDVdgR0RtAqqHba9CMGd1Q0D34sm2pUhxCL1q2TvzEYYqDSxjJ+EfeRMph/MwD2OX
lAvzsfz5PtslxdLlgF1o3j1Rq72z+jXvRAFk+9P3jYJHOf0tuEKBTFC33v1iuWJVcIDfhb1d8HYL
y53O8kd7XLZZmrn+GbhYbibYYq0fxEwnBtXM4hplOpTc2NjnbGD+5hYsfsX5Aaar3K7KNnQy0IaL
uE+ZDwJ+GrRsLuwCskdusXeWHErr/9qekr50lxfOjnJyUKHBZv2VooN129M2Jee6GvQNgFeHvrP9
LblfRcMZNnUEDw6nFiw5g9pBPl3V4G8LC6tkhZSOnZM7s2H8PhmCG9ZAWLZmjl72NKohj4VrHUOm
IQaOVRR0riED78J1WrGV9KFixt7aMPQnCcjCeciyIn5FTb1kPbkYCSoTeZ8BkSnp+/V98w+32I6x
6P/3rxcaew6OGuxhcVs4pDfOMJSQDa1EMwJApYh7JZuX/JYDEw2i245WQXn8ij+3VS2vVOSK5H83
J/7b7RhHCjzd6xfSQMZQFSWNdLKIoub1epZI6I/S3BvDH4UyNjRZRL++5iv1y/aehB+F/yjFKlos
JZEEBoYEkwGEphNpdxGgQYgnlupfZxZWGteM4Xwl90r3E4kxzHxAehnlfz454yXlTXUHiMiySBkQ
jEe1BESZUAjVKTJ7KsHo0MbHI9yQg2WvKv13+0vNDWI9ts3vDwqCLiA3KdPahtSDE/AOxEyMiOr9
6zMDqf3E35M0TUWUjERRIVte6vESN5TuKf3Hab3nRFvXQWhIt8yD+PKITYLqUvg2vudx8RZQ0sCO
25ZPWL8lDhJVAlMTDbS8Zh1a8/WMINk0nS6UM+N5A7YHTti4JBKNskXbTVEDav8qHOjPwRJWQl/d
UmeWRIEPXZr4EUvz/AQKzmLT0Tsv/hyowjdLCrgdcspchdLWWL4RfMAYaRLScGrWsl53aSjq0MmX
WZvFrJw6WHE6psR51ajkgvVGdch8z0Hb9sliGT32/o/QilDKqkqXpgkKWEECAnTRyeIpRANjjUSi
bNr9oIZnRIckcss/Mp74htNFq7sLc9rsC8nroCU0KamHewrM5VVc7mpvovRbC7P72M3fMMxxPgak
EWbnvyXjOPNa3Rru2kHzrBOXXeZQks0wvKW87R+MWbjAuFulcerVqWlerKEc3dLCy7uwQzY9jk6+
KeOPyVWsAKEN+Jw+fjzMxoMmqEfa2VnweB/H9izmNYqP85+4Yi8G8AFjApUPrPgDzoj03cjvexe9
FMPqqLqePXbDAyWbTWwYlerCL4aIC0Qf5VX492Bbmqh59WIXlkejhzJgxkiHPO/p2ynroWD+Z2zm
/IeeUQrCTSKjFfPjekHfT4HRxWPeLlrPivg5ePEbaVOg32F/O3YmOgPXek+wkEduTjcveRHdjDRV
sPe2N2Y10GTF/ijYKpZ9uihvFY+Y43zinK2YnbpMSQS3ZbzPDQpumxEhjGVHDcEns129FMf6va0d
JdnfzoaKoISDk6FveE4qhdEilQYYWLCEjb/LMkO9xcaUI7X8zcNHkZYc2hN0dYkcKOMwJfeFeKRl
7oTwziYnhTbvykJrrvq+/aEKMftOwGHzfArB3WYl/Nwn+43cXwLsTUGsj02PL63ql+TCaAizry8m
3drv7tdRAi+0/MTuIQhwrIv/SDkrDYtjWO6xy2f5vVVMSz/1FDTguHBnmPJe5SKKFemkzhYsxbo8
R+JGBjfHW6kRkLtScBdsVn5K0PXMnbgkN8Xw4+9Ct6mylNaur9fLhUmj3P5h/U6XNypjpqnnnDJg
n+GIRNx67WmL2bxQx18ehybf6eQOnRQPqrVOIFibRTm0FFIzZxbS3CLUObIY8lNdo6ka9QC9bLhV
0xwzPT5hJEzpXA12MRq9Rk2m3MRjy7GGtxkB7hFzYDWz4C9z5hCLhNW7bPhrdzSEL3cLWZ8gUNN8
+H9/hLwmlaxQbeZsPQx1f8cKcI6qw1dgnA82VMXzVpRCeOt10Jq7RxzuXpVivT33U04gWmb1rihK
Hzk1VtvnCx13RO5mA7yNAtSPg/0rFBxL79Ddv+VJQu9syyiIgpiZn37/28Xt80TUgLFJFSYNSrYS
lLv2oNjV5oNazo78ydyfEslgr1FUCibcF/YU8RM3TMVV2QcDxXDUFhbrvedHOT5sdeqpvkdqaocv
QpayJQuiqxnB4Q6yQOugIasnsGYaCxqClSsc0eWjWDmj2NJmyoiPUyhNBkVRVcUsLhezLtpiRyiL
U1568JY4LWj9kT98iR+Dkwq9x70dEB6IxXYewwwqibF6UQdlvCvgQzN7TpOwdHiU/MaFZz6szI8y
NgF/2dAZ/84gNHlpYMeyQ5oCN90qx/C/ITk7ad7KqrGYIGcH1luLrdSoT6rBssj9+TT7cHDSIchk
xq7qdPrqtRhsfeX1qlnIsH9p2J1N04YZiFYqmZr6CSZUlJZ4G0h08dPf+8OKvLUclOW9ppHm3E5r
aRK79YHjeXMS62qYeV3gniwVCvUw5EcEZ/i/sEkhbxvXD4A0qa2DyrF7rBEID1p7CgsnnhhQ1pw3
4oueIjzSqsDqXToGDKGshnrn/98o+BjDlVq+k6GauHj79NZXYTs3NhC9ZiEWHNez6Eh34WB1LFBe
4/fcvp5hBtFvpLGnF/Bplfl2dpxQWdvPjnWgZNjc5Rd3QUj4jN3v+Dfgo4n49cFjziWu2jS5yMfQ
6ahm9ogq9Xi7vc4uZjzm7TKqSdpVQ93ov7anhbTGeZw0qOe40fMrAdj7XjWA4s+5YZBA7AU3eVbz
Ol4Z/bsnzM2HE7O3OYWn0iJuAJZMcjpHOTcgpG+eSAVi27E/M/kfw50q8VthdmLIloLOQ6qkm7aA
M6tdw6TzWrRI7WEfl7HjaKCOKmAsnjGYzSgEcg5ePJvryKKRBe05hHwY8x65pUZK7n/7XWbOoZTj
IKxLKgsekYHsi3fDYumn0pgpyReA6IjFsLReaGpqiCaygHKlsuETRqPvJVzS34xtUguHEaF4mtPy
X9bAgfta4Jt7h+UwQFDTbcgRBx6LP8XPZzNR9iwiCkzKURc60Q7pmaTk3MvQQOIMDMV/x8V7gdaN
Rq5hmECW9IGInY03XZt2/j95d6NTJAT3h9IxIOwf2Fq+qP+mtXNN0FKbgUVL5YOK1h1jszIbwdzb
oc6DSYYTrF77Bbhj5H3O1Tx1IBY1783uQ6IO0foYt23E5CN2LrAmIL9wH3JS2g7kAo6VTFmOCzDS
z6TGZ6QcKz66DOT5LHqhM4dvL6FRo0zWOp5phrrU/ch+k5mr0Hac/6DXk0pzkN3bNtU+PKuHfgxn
fVIFyM4CM5oDmOIEt1B4Re5YPtGboo+/MPf+U8wt6S8wv/9mIMr9QsSFPe1xKocT5aqn1AqzV1Pg
gxi0ni/eh9eTBS/kIlZX78OGqPmxllZhAYU+BjtSarIYodLD2nX/ncAdgF6X5n7iPbz/e2TnB271
/m/ppv+Cjf82f0dYRZGy1aYlOBV5GNFhjiHcU0YVgA1wLbyWbySxKWCFaOL86M9kRUuHv9uWh/FK
NFSEUrX7iRESS9L+iXHp1LSOxJonZBFsHMhYgnAoO8GO9XPRZGeD/1wt/ArTUli4kXsbfjKWqXmS
a9LDqzrlnDCy9kdKgzLXqccizDoY7csKbovWFHnKWqviRE9RLdjaa/WoOkXHBbadZnaAzzuyh8Nc
tDVZ8i50l0VnTD5jU9Lu7wcXAhXC5ttZ4FdaMDEHAhMwNw00m3l371mcQtnVpKhi00A5te4fcBMb
SmCsZZRRnry0FKsaCmWb2emc0SnIWdUFMWXdKONh0xD0nXOBrI7AJYx3cDJ1+m61woMY29yoqp+I
SDZjf7Y/rbDHBFw8wXx0F0DpRmCGJ0tLfj8Dxyi00/VuQG47uUfKR/eNQInOoX48qaL4b7q2M26m
XLOR4OPpul2/8MxFnfwt6nQ8iqJeZH1CoTW8Xcjd/X8EiwrREc+qYdaM4qbPnoLY+F3ktpU/U5Wd
rKOy0yCV17RzLxKgV4GpSnFtUMrmkyXeWHFrLHlhJYNR3kpQDz9s34D9SiazxQXEeZbj2rZlRJ6N
FqR6A6VETaChnohmypHzy4+N6THNTeUpjs46QeTRPMA29dpebhXs9IteL3mUpTcl+ib3Jy86OkQr
pOIuVKYArE4ts6oEyp5RVDzZ2e7jWe9A+ugzJ4RazK1FVoiMrz7RX1e8FdTbla6TOugt2/gqhNqj
nE/JT4hgHSb3gSAjN9OqIne1/J/KTn3o6yeRIQinwZ/NW7gKGJ9uMIhonRQDm6TsJfLvG1MRlDO7
zgzTUefFOH5hV63bAZB+1xbd5/qdJV+Z93TSYlpKGdWY32NZ4YeEjgvt6gH4d1+ZwG76q9cnf7m8
EDMXHiK254ReFMpXl+yLEFenomfwFfVnyq3PubnMODC3FS6cMp3NXy0W4R6987+/OwOPhZCUR4Q8
SZDevSwy1OAP8WMYszfzRRCrZvxwocc04FvviEuIjC4lYir+9oOQDt72V+9xqw63Ore6lzYnU7mJ
9hRQuVtlZH6iBKmBousbdWhcqJgAYKhZcbQU/nioS0wwSYLgRenGpswhbLlHAh1n8wyi0Il0yy60
HRx08B96FJzbDw9ovLqW1z/SdLqRuNsh4vGoOnDgkFrZZG4ic6Bjfu6+2PrVeH3wip7w6B/XveMP
TmwpX2/ymP+NYLDf8GotMKv0qWb8xSoZ8GnD2SHz/ueo5GDRtPFlrz5wrJi+RlQIQA6snLNI+3qx
IUE6NXUbgW1+zNGiXzh0aHVqSr+8675ojwxJaPUnFxYgMd+u1doGWmqQYz2FvSLNlFmkunx/+oGg
EY0EwUPHe82gjX+XYRZkQScC66/zg8yfrg3CViIcuPsROPJnATdHofjqvR3cl16/69moszwB8R9Z
wIYOx3rR1CYD2GiTwmL0aoCVr2lZOnXrikqT3qWRd/HCYl+BFt6YlyX3AlutjveNzQWddnUIjnjp
eP9wlDdyo3iwSclpu4rqAPfaxidTta5LQAno/RTB8nRYdIKo5MllXPfw76MJmr19FrnsOggU704+
M+E28Iw4zu7vjj32dvp5W2T8AOoTkPuS61jT/O8J3p4goHqfIZN4RIZ29TK1lMXd+OpENH7e6Nj4
VxYdssPhO4lwMX8y9JUkUWd+pRneaMeQdEBga11BKyi/OjZNRQMV6IUagz2wp6W2QYIfnJvIUxAm
iprKVmFHtyP8W5mAoAB8ccg13S22kaCghYSx2f1Az61E0mFtSyYcbawb8ZAeaDcdo9LVnQ8suhWQ
W2/47qI7UMGWzjDhM8CxKl1bXE2DdJAk7AQiExIgIF4wWT47CEdVwsgFo+W4glc4/VVX64kPB77/
2aE/cdNBPn9ve1Kr3Ut6NaDjRdzl3pu9Somg1gVxf2XDgdSN6l27CX2RX9J0JMhb4UiEVTNje48W
iG8XH9jIrtBZvCFc0hteyKgWDvCqLVsotwhEh0FTmZwXs/TQh5Ui4xN4uh7+GY7e5nMp18fjMGe/
guoAvNo70N94YjH5+NMCrFdWWPWO+Wx73ui9a1F2CuMmFOupsGvnBTlufULTYVAZrVyz08UbiAdh
1ypd6JcfNS42TskagrSI2NdcBkk/Ng4dLZ8ZtQyjtnHAgK/0rPWeHt2e30gTr0K4G9yC098axqul
JMR54DnMK6GGiLIhnzKQiHBSHDg71+VCk4SkPfd/bQC/j8RIRSlYG2ahi/xz1qYGiW1TrF47gBti
uWlf5zG71qrZvBjTowCtvlRt7apg4q8enyOUorSw4txklWpwY8rOOy/APCor71qjBXWXprWuYlaG
299gnYZXzlqJaqmbyuZxxLYGYI1ICedGD4fO+YZnnFXwYn5AhF9WrtTddb7vfO5ClH5f6YvIte6H
uZtZJfagyvqxby63+31mQ0IkvhroykpfchkzJ5QEQFIw5GaErvejgQ7COho4rhlxLYObHr4ZrDRH
FpY7aOcUxYZz0077Zy4hEsWrwKahYorRPsDfnkHdyaWvMrKarJiH7jCU+eEWO2bIcXkp2eJDNibF
428ankwVBkzLgcoRclU9vdtPetOpmqGoYt88YiPCF84HXDCHujgCThgtLZYGb8gnzOQ2e3Ei/SPb
ue5ZUA39t2RxDBScNVUW0h6C4Dx1a8L82uvKa9TK8rKUaXWXVBbHXNAS+NGe381qEHfjYxLR3ef9
IJ0WfGbBQa7sVg2VPd9Tg5kUr833zprilZJWVmeT7WzcjeH3CLjuesVtxYF/qRMRWw3VAQJApzOG
K0cRHD1V3U442ZNofoQY5NH9fKtoVj0bLz0RCdN0MCTQSKaB6qwoMAK3BpN77qXpbGh4wjqIhodR
I0d3iknIXx1f4gKYuw7YNKKK4Qs1N7n5e/kj6gutsgWDrx0Y4sh3Scvw+ebcwWyYx4qPGPjzJSJH
gV/SVa5+7RUOCAnGMacEdKzZpLWyl2hFZv9M9+Xag94KhhOFgKO6m4MjdLJgtSZYISqAMVOo3F2O
U7ZD4B9O776F0svPSfn/9sx1KD5EylC3JcgerPLv/PeBkbWwm6WFs6L7o5ZL8ZvyQC/lPIhX/W4H
xyaH8hey2yGD7sxbvG2xw1p+5f/y/iQftnrEyMi+Mrk+uflPqfZfbdnkXl1a+LwRuAgFwyGSCvpX
ooC6rcjBa8V75e5nH+tbhGxZYAXuTg6enhgvd6k0WVXBms8zTzEibYuSGZPRmodsvZg520fGtFa/
WivN6igSRdDbdyrkoTwdLQz7SuY17xrrX2VKpUivvvrI7RrOT+EE19NtO5KbhpPHa+5TQVZ7KZv1
wrn83cLfBsZxWeWDNwTw6cEqNCPIBRD16JI/9fNFauwS3e1G6kQs6jmKcpmw1eAF6UhT83eYASFq
NixEK6k0MYscr8fC+VFPVBB3X37oFNHoRjlE26jyXukwsOhBv79DZvCbYDvZdKu3DJmlE6hmBHX0
5lbXrtcZwxLtmMvnNbgsUdAhmNcmDXNEFYa3ufrdvtsQdndJkWAzDxT99XctoI2QxEvwoTS5s2+F
Xx0sRq92e9yPustk+2v9JtV9crifuBjUvTA/oE63EfLkZnwBN01tdpht1ne54rj69BZGEj26leR2
woLW70nHbssR8/q0EfeNmuQff9/G/m3L/FIXjPXbCFq5bEWI3N/yg4XV77kVa4DhA2QWZbe5ZMrH
1snTtsoNJif/UvsM2s0QPhgM7HCLBnGb5FIjt4hJEh2+fNrUKkw5u1O+Kgkw76L1EiQ6jSXEJLWP
s/o8vfv8/fC/tax6NIO3aEgtgHEijA2uViZKKMB20Af5VHJphHonzZjDnDRRyR1IeQZ1Xx4bqwOq
+VuyU/iXWziI3eGMCm1PsUOCxIrp8cAPnJ2rLxTd4g2R7wmHHr6D6DMehGr7iLz6GwkMn4Bn5ypY
EJYvk+UPDQzg5v9EYVREmrqSRhTmXC0U4MLaidzJ2S7tfP5ASMiN0A0cWdRiWLR9EWYOnn0hFYn7
+9NFXWsKeMwgVddQV7qJqO5lS5bsNqkwFffgqvZlCXXBhHerUHuV3hh/FlWqHN0VYkztdJTR9kwK
VsNHLGoesRcvHoiR7njdDgdyGu/9eOJO20eZgPB+AIaVP08+zb+HL6uut+OCPyAbExvY2HKsyS3M
E6MUcar46hFgGNGO9XSu+xAkLXeBSj0EZS7gQ3hU3JnoTzTa9hyA6dOWA0UAdzqNZ3MUjwhiIX9E
KdM5yCOlYMlsuuEdsYbAg+ca/AVJe/WBewlI8vk4Zy+2dSgoPNHAiCS+7ntKOW71qOyQJdihXdz3
epvSyU4ehsszAoIQbtW6Xgse12oMSGBxvrRwDNcKsatUf7DoakfRZMWKyyNm56CLvttzcF1pIQ76
KVw3wgtn5O43FbzICy3YkmtWWe/0tv35OS9veGOOC1NianNk4MMr372G+Zm6rYu6m1h/xSex9/oQ
X8gKXWnSrcsR2Wr3wpbOwubSlWGVwKH6jscKqddRD13IYjGDMw8VWKTGxpIZTU35Y4o3YJqz1WU/
tHui9nWkgXxJhH1kQXRw+CMEAqP87ibadflhpXkgaa81lnYckEEuUGtkDIefZKd7LeZ5YURoS9ds
7U47HRC8WP35ye7Gjs8djKOJivVjIbLVG3Spo7oxoobzb0gXw6GNa+QiYghwGX42s6uiLMbdvrXZ
9pjFIFzW+COretMZEik2aQNyeVBKXZDW03S1qdZOJnn3dYgFs0cPyXhW9KiiFJYZSvqMj1QBIYet
a5L7l5ju5Z9UzJLwsDNrn6Wkgt8N3ULiC3Pjlx0tHHVXBr0KyxgaJ0WZjdai1kqNXCiArMKnfDou
C4oitMctXsYRqpjn3ySB9eGeXyxaqusFzVPubB0mkiEORF0dXpDwAMT1Xe92bNibxVPXs5ahNXBR
crUw/LkBV6OCtt/MpeqVpNhaXbHH3+48bw9RFEqplxPpJokuvmXldk7IJAk3nmsM4m3G0nEhzgCF
Rmueq9XLwRuIZqA6j4HEoPv6OLUruU8ZEKTOi3i/mfhEl/NTGUHetdLiV+Tj+TUx0kbsyWg0Ro7x
91L7svC2wLJZ5VbQXUK5SbHCRLF/GhHVUtk5G8g2fNH7H/FQue3ozb8sHzKyPTDsObW5bS6mHWkU
QL2Kv+A/9DieqH6OAm+r+uqsA/2QYVmu0MtaAwIBHFtt93OjCbhpeSwjaEU0EBrPNb1itMPbe7gK
+tabPkr/UBohS9L4AgQDgx/xS2BL8slfFVS1+mgkMQxvpR6a4AtSEGj4j4+1ZZ6uZzQI0sdOMfBd
PlHke937lAH251Bkdn/Qt6g7xm5lOqVHq9IsDwSpcOB3oMez4RiBgTyYs8K9h8hF0bmxnItpgmvL
XysirGeRDfytcWYNdr//65k8RGc9x5QtG92Ggp5l6SB74X3RMPS5zxGY7Ij1/AvrRzQedEcHgdeq
DR1iI9RMUyXaVEDKELKCQnGzVeeBSIv45a6FdM0f8wMD4XZbnmVH1uXiX8YUEqOFFv7iFzZ4ZZs8
GxHPX3lZd50WiHsw43De0D6pSwKowo9y/qD0OfvyiaJEccEpar7RsRzGZIOVcjQFY/r/b3zZbGpZ
Rd0PZKOFMvoym6Zv40fwpIiYA8ViE5bTfpDeOlMsXoaaF1DrO/RfLCmE7/LmANS8O8oX/OCAfoxa
WdVx1qHODYdLvjRARnX/6RcleLNR99TbUVJY6ETqRo0cV0HL4Xg4mlQ/AtLWjkCrI4YYBOCjoxwG
EsUMY/Z5UviiyJ/enEJByfy0CJ4OhxpBGwLKs8TjaRvT4zPjGeQ6fZK1erygjv40BLPSvW5qur2h
4SO6JEp2CDE90r2KDwST3KuRRbtFNKqMmtAbhLCghqDOkZaO8ojK+PXnqlJggWx06OG2Qrgt1sut
icJioHxn8CIvwQdoRw5dfSaJj5+C5pejzS3gbQYYQlJrMgKGbuUGYoAYMXs4+O1xLKobgLe5hWXK
I2vtqEssTqE9iQAo7Cp9fRSU5xrGpWDVVDEnjfNjaD8o3feI1AlpN3Tx6NsmKME4S9h666AG6PJ7
SP5mW8MdhM1VaNZ+z52E1/V0aaxW8XuviZoL//kOZu68sD79zbReitO+tS6J0nN8envx/c1PAHDE
loKx67AsmzqCpe2kID6lkhEtRI6wxRHTn7fTEXsWcgVV09NcP2dyhNT5HWFH16RUyW0Z/etWFVWO
1JYi2Ll2nu68/LdBSOml4f0II/+Ri37QT5qKPXmsxdBSRdkuC7bBfZE7hg9Af4XT1yZZo1WvjMKt
g7HfSAjC0en65LZD3/kIAVldAzTok+VkGWEDmAhYgiAhsCnaMKkeRk3oTZ9OhyLCcDDZct+cP+Pj
U3lVabmrwk2vb0od/fOPTsWBUMCegtHeUhp2WP7AQlEaGsWvk1yeepttkpmjUnzCHP3BoigiWsno
aiymIWrksF1ZZADB1TfJVwIQXfOX+ocMOA7Brvp8+vgmQxQsSwgu3rpQhKhHD1vThHQF+tQhcKWU
boaQBPwvN1ThXXgcsUCwusdUg3m/71tREtRFlEP4tVcc6LyE4I5pkiJ5zqlM1fDeIrl0lPURFMe/
DXCldDK3rpNiOpB+K8LWNs+mGjqOpE4Xw5meUEtA58KR5Yab7WFngREpOeTFl9oIn0F7VJO1jI1k
5frdrTV2U1ZPZE54uUUPY3e0nsKp6FHT8oXCmV4UOt/73hsyZ+CbjAmGaFXnULXdTAz/3s4sMdqk
6CnJzK4LXsyo2pm2Yt+LfjyviapZdr5SUPxo+u2ql3SxlvpOIvUrv8c0wsL/YdoMwvV6+AE491Kf
jAcGPtB5qAQ/tlTvnD0HIa//WG5kg8jLiljiYs0xVx3gbF4PPCOAvqXN+HI82eB1IRe+gltrJl8L
NqOwPfg39d15ajh63iBv+lGPAyYmWq0cy28pGKE0+v3D7h6hWUdAXi0aQ5/Gu3ni3kmohbB3WpXj
0b3YzwST603ojwxkpo8AkFeAqn/vDT1X/W1GW+MHbv17Ch20V0C+ggn26qBwO8Jryd5hQ/f+PGP8
HlTEIYIaAWrTq/JFYs4FCqr9bxgShGZpX3oiuh+IdI3f7MYnMzSdpYZrL4p/lpMeT0tjznMDkHeA
5YBe0+GJMZxvKUpOtsXHuAC6dQCJ0SiPyiE2z+TEtH6J3y7dG9zN5V27y93TnX9SQ1HxlkO5dydd
mOLQt+Jk7y9FMPOwk6ZVeH23ZSq5I8FCjoUD+gkRTtN3J9waq7lPJeYzJRGdNftyAMUq3kNMBn2c
UYSFNsf2S08Kv3dv1Mxg87Y7APY9Se6WQyd4FW8i1hC2SWTqCjuq7VYD4WzYYIVrmJopfWugBoS5
6gUj3ZW/1QvYQRcSJcGPGq4rRpxWWlp3E++1r5DI4vB1Xo3bZLaIez3MVql0CNxJ02PucAu9R0BB
5e70E3NjMwhQMO6F0P7QzDr9ZhjiStyqxtQKd35+vf85jTFHqTrUNekm8m9C2+VU/olYa8Y6lRct
lJwFBMMDfo9qQQUzYLW9fNAgmhiwZUPAcXk0lh7LZf8v2lpZdF9FiPdMQI1wp72IFFQVyjxZE/wY
pxra1nI4+E9KAAyypeaQoAYwcWUo1ZgzzyysFwHuO41L01gnec4JPTii5y0XfHrym65Vy/YI+0Wn
+7Jj98FwrmfxjJEDGn4kZqA3UjtYxMliOFNP6DYETOK1HZSyBcxZo870F3JKGzAZhyZCvyVlH0Ug
sQmIkZFxI/c9nKcrdyJ63B481NH3+0OHqjcohVc+q8oC/tNcaaCBQ9a9LHy10rLgU7qAgKOnzf3i
KPO3eJsMdOhgldtGnT1cwO17f98VRlXTiwLC7QjhywFo990alNv0+EAmOtZ7pw/Pj2ux3s/90joG
SgKVmEZ1yVdbpj9NZbmLM8oYKBzZQcuPlaHQrMFK8gSdDhGkhZuVp1IfZCLWMfT3zcOido+zzbma
+H+ZXIySh7HgcF2F1KqmHehUn1MFnx9wOKEs4y3cypl/TUCAMvGuz9g0AV09++nrZrPaT4GTMGhL
WTiZRD6F6bivnR/WSgcPTO3EkifaywS0+J5XHjWsQJ0OS9TqQIXx8uOKOSBUqMJGg4rHjqa0k5ua
Gpbe4voxrfoea7AfiWSFNoMV60XFa3IX/zNskWMdxtLYph/h/3mcJAUfOCehDImVDr4I/460J77W
fx6VofojJ/MET/ewv3+L2xFfAxH6qDmP2HSrzpps+auc0+hDCrqSuEJY6HTwdEovDHREaMBK/A2F
miJp9yry9YPb7Ypq/vi4VNql2fHPEKtWV1FQs3vFJxfQ8A89Gzjmft4ETtr/fsMcY8tX12Bblcwu
GqQfYPzglPHKw7g1WuuT2QWm/iW7D/R08zg/eE2yQIcNSw+iWD43uP5GRqbf2qEUp61Kg0J55fbv
kVXUZ4c1wCTC6ANVCiDTszKsm3Ibft+XfToATNql/4F6JTIMchhH2791LdyRUGg0QToarKlmTErt
UfaEwts7B1qTn0FcX8sLSN4V7LA7o7QR1urX7HYHSdO56vccoItlTMPoXz3kk5xfaQN6gbMmb5lj
+cZ+U7vHkFoJfEd5Om4fxIXl0EjpSMqs5DXpx3+4q3PiUBTA1TlshdBnM9G9M9ZPHxKn+zMjTs01
BmlsJrUkOp8YBvBgCtr7+Erux4Sf1faKVtGPuBbVztcaT0Q/Z+tRHfOXKbly0PxJgYZ5wGTHijXV
7Y4LycdWGrDLg78j7y+395Yq7x1LsdruVbf6LT9m6w+KGjtdLYQmzZSe2gjY1kYD8FxNJP3TfxEE
ujiw7NdK+Sfi+uZwAmnrQcrp5pzKWni+G9MjWd86uISas96uAgkXEwr6v1vkThMjFQFR3eyaiGJs
yROxMZANV0yoEl0ELznQ3Ju+nU1mIduKtII7844QxaviOliJSwpvGrdemNqATB3KmhKmldQcBUwl
eJuKdcHW7WodTE5uuYsyPJe+EenKHYcDdS3XDmXJZWEkxaJdA/dxP8PtQRwp2Oc6lcDacS+juk9d
yc4+EPhe2yA1paqajc6fArQsELD4YJ5Kn8mlaVm74WXRbM4hajT+z92sRowT0T864iRXuR42CVMD
L9dF7A4slYU9cYuC+OeZ3A5cnepZ4Iwd7cF/80H2FOp1brTcDiMNQTS/Xo7RmjEcNaWjFuKIigPk
CV/c8O2x4rolWQ23NGtxaOFNHcM95ZWOATVEG7CJ/to01tM7Zmul5/cSQEQje0TiS2IQTYhefnHD
fdxFwhm2+arAmohsI0+IWu64DGraHNL+AV7ZrkPuq+xB+8qx5+nrFhX/WIaG367kpDmKRUELM+bC
k5XoInxk/nvDaj9ulpqHcvIPkmbPcTo08ajV66J4BRZohjnsxwoh06yCd7WUkMOEfz8gKkuqO/Yg
Z6cAHWBbZrD2ezevQ/N8m69xYS9FapedXU2KW3FwQXXpB+LFHBAZVlO0h2CVurJYvChxMOy78Oe4
i/bZ5ZxqOlHbPir0N2aR1WkZB8MX2Ss3mzqv5fnBZbr8cfE7IVRWnzfFi4Y011w72gYzFcgCWZwY
Tnhs6PKPxSlEYKrQrEJGMMJrhZMEj8bKgt2uqUZKs46CgDBwUUgE2WkSi3FOhQc2qjq1/FSjk+xj
DlTm2aV0YNRNHmBsEHzR7KjpNeSua6RYBKdzGymA6zMHgR/Tx3vJ5iqziltc38vAK6+JunObN2Nx
dRFF7hM6phUCViQDgS7WB7Cx/fSE+1EJ52+ThdKJtQgibB5tua2MXZdn54LltW42S3/2j1+NDoaj
oq9ft4kQT55bv3yify8c7UouFPcZh2UfAxtvufzeP8xhDqmjOiHVoybb2ToISRQhIvteQh4yl9NA
np9L38fqT8tH3vo1gjpwqpagnpmD6G7YLTQv2Oa5BTWlR1xyMM1X7Wv/hk2hnUXjRV/hKV+z5EVg
hnuAtbkABZ1QLLuI+JeHe544ts06frR21pdIU46C1Lu/rTa+WK8piydSddC6RqqE+cWrZ9nSVnO5
MWFbqckGSEYApwPFaTMntN+LhH8tZsQpbDxRmvmiXfke5RfcOMwjYV+Y7RI1qZvksh8ekphEHD83
gGEHE6uMjxBbtwg0G+m392VIaRZmIW5uz6WXSISwZczhPL923OcGbG6MHXFBLlHZj8h8jCwuY3Xi
PVjcmVcw2/boI4ui8EACFYYCDlOtur2DOI2L5NVt+XWTIo0xNIk5EH03DOlHcHoC/tvGN+13ggq7
FDHtM3EG4QSVih/nuU6FlIt9Ez+ku2F57wJRda2eKFQlnbxv/wgCWPVY5/PeCLlFha6QgcPXQgD0
qO+J5yFCGyK/LvODdQMOOsxWdGIINL37cncEI6AokPQzK5pKGPLbk+4GrfVtvfF6iI4uvGkIvFg7
/2bjBh7z52Zu+PmBTAdMhh0T0iTmj0MzIlh0UYGBXKUNUX6KFmpvrwsge3UYqaLcKu4qiDmi6lb4
pJ3OqEghyuztZdx7/4FYOvLJDUmymMMy8QklWZUnRp6BgZ8NeMTigTcaOaV4TOOQ+SfQCm+G1w4F
Oy1gQgXylOvxj7hroUd9PLIxr7OJ+yNIzoz9nnQ89UNaOysRYzKD9up3HlWZuIPc06ZwnjNZejEa
f6HxaieVWvhNvUds8MBT6q+4G1j3MKtLf3N8hOAjTc/pDkC81gRa+SWzzwXr0BJRE1DHGRr77Mo0
PuJSq4XKsp/QqfWR7XT114MLHvi9bTXukl2jyqyGadAIcHB/5Yp5Zy5Oqf4cDXNw14h38JdNnwTz
uHhrPGbFGBf7UNjdEyT9Y9qrgojb5ZJ+SH0YSgRKJ7GUSba6gFCeBQPOEW5VRIm1CJXPXJapPBT+
bjuOu9GZoByyurKY57YczYA3PnIQra3NgdK8YSzVFH2FgkuOKakAIOKbdmNQbYuHWTKQaP9gk4bz
fz82h8A7nVzkLARDC4QgM+CaRkbWjM/HlgwW/9xvf9IadMzLbqp5Xfvm8j6QL0Vgd3Wf6Paiv0AE
UPraOPnICrPaS4YYrOp5sNpvBQZOPwj3u7xpbLMOFxYddftjMnTKQ8Y6Q/M7fF223TTLB7KAB1DX
5DRrh4KNgZPFzYpT9sOqFlJcDSRY52TcJVOXiKk7lh9yojVud9veUteH9SvurvN5uLFl9c8cDLQl
1CpgAPd0t8jCXYzngfqTe8GSbpoPCItJqIBl5epkTAJwaLpzSqk3rfb0SB9cbSN7dy+sQvkXFV3U
2Ho9HwDFOm3vJqy+phRrOZeSX6YdPdQHTahbY5isB2Ut5AdwWsyLbkZCXOitfUUf8O95rGC8ytco
8LpQUCtO+MIcbvjxoz7ylIX2vN50lH/D0P9u9KTGLlj1HWw1l1OxD9ZiDX89NfRGy60HL7I98poI
FjAGXqMNLieTf0KqwNJ4KZf7dGHENHe6Jmiqc+TREDsO4Bx/xpVpeOBjr6ZCUW5A4K1xhzJfzUpF
RfNIPI7E+BGra4sjocXyrx0Ctveo67g0k+7a9TUYDo6FntqkqJKEd72GKYrp0I5goNFrfa8sAdRq
RKcDBo6w6f+gPDYfawA7+aD5GLt6enX/smv0URDPG/D86JPG93nC/828uA0qk760h+7coVg4bpDp
B2Cf/n/YeTYG/eXF3K//mY7uu3b32353shtZXl3PH6RVxbN9fKCIbDCebpqi+8oE2ZBbSSsntUAU
tnr+9Bs4GL19VWHvtZWsvtct0C1u/eWGVvsN+TzbfyNhECWkyuPqbWuXq/z4DSfSoQLElk7IL1Eu
K2z5awZkNkvK03Zi/VFh4aC3N1NupSseySdvBhLwdwLg/3E1wmCWf9v1TGKtB/o/j1FeEKUjtvvR
+FqOLsBcKdGO9rznMN4t6n+JDfmeJj+6ezXfSCXZ32USZ2YRhDrQ3eZyp+IB/MQi5prZoLfjClTt
qfY9UIhm5wEgecM/sT3gYXfqu6Mq1CciKRHwi1rh
`protect end_protected
