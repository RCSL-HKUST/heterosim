`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b2Kv4L8DtlmMpJWsZsFI5/tqEbxQl5x430SVGXzPAZ9nFXv9Dd9fp7Xo6tMN3Q4R8CSm3TdZZLjln6dY8uDDQA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gtWcQNrG4Xh30ok0hwABRm5RWPX155JN19vkeLFk7m3f3CAONNvLylswH2xlnM3UYKP8NMlMFghFChetHm97SPFP3vRrOsneRHwov8E/eT3yBTJPuMlZs9GNM4JZ0l6KIBnV090jASj2hxtr+oRd8IGXGt/6k8NoDnQUhdpY8JI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cLMLF5kt8ux1Y5uF8uq5js3GoonSH2YqoqxXFNHksB7rHqVhNvzvtmlzwCY4fxMhQ87JnDO7vRdspsveHT1mBnXmj8EJxEA89+wkf9LsQDof0HEK0porFf5e3XrH2QIYBrVRGIz2z2hzV1GwhxMBMUEV2gVh83T7yyAZ9yo5CMZqEbKsrmRvnX+C0kWuZdg6lQSSZhxIl1jFzeuK3f/ZsYvRTe9ggNOZ2z+BgbyK4f46Db36pK5JSqqlYjzoFruHhdl+3jWP8p0743QWuVQklKtoDMElbmKyOphu2CZYXE/Z2m4OffrnegjgmJazlXvEYt9CidcuM91zeXwGrtcyHg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hN2X4jGOsefMSwGwHiHWuxiiuyYsaGhMwOUHFufVbPYrIqR8Ul5ZjAGqCAU3zXB28CNmZC6cW+dsM3cyvPvGKDVSEup9SIm3W/PgS5anhBK3iN4Cr5n65DEDjq9ZaKXwkRY+X7f2lP1lUV7/X5YTpBgzGSxNNr/aZPUieDKM6IY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZN0tCJWohGyfV+jkANna+ueNhaasrR0griUyB1YY5gcqBtB6gnAYicsa4uG36DkitBdIrQ+sNhNHSAWGLtb9C/ZJwzwbzYy7XK4cg+BPEfeeRLlIXYyYjD80nupUZLmyYL2R1AJq9k4tl+gEfzHs/hhuwpA0nIMUjHFx4KGvexGQsL7OYKfe0exx+Y5DELC34hZXs0+D/4fOye0xeo13ZhNAq+MDdtz5iiN3cdJRV/JQO1bK/zf2fNu7nmElkR19KMGo9Wh3Pcl2xYD8w1ZAoT1DqvjU0dggCVIFFD+zxk4zWlNeAWRc53mmCpJGSIDACdeIwzrXIgHogmz0A2FJPw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15253)
`protect data_block
gmW8lFmYN1UbMhyrdLfAUIE9yPM6fqlVYo7H3m3T9BkP06lf8SU4dSZCeun1Q4wbWWOKy0u7AHTS
2ayyfzMfJsAJ1lcDt9Bvc+wP1kBQFjuILosnRFm5a7U2OFOXbw6mWsg4TRmZil8yqCVUrMW3ZSb2
ryjlxHqucthnCti5rtcoBt7vKcaFLWKsOOmWXpwESHU8OnTliCgb5TOa+0CM5WgGMbMWL9iLfjKo
9OSxYOp5U/eq93IYhYZmDlKC3GAzotD2dGhepY6zwrU3Z/mHRBVRi0xPOMl4FIsnUZRdzw4OltdD
ilP6IncU/XvMdbu4EzZlwwoFm9JNrdRUUdgNDwGITP18AKJ3hPrxHRLnaRt+0X1tjBkO4xK6R7L9
rKa2OI5OyPx+fY0fHdVd8SwWPEfn9rQBPt+ua6KL4T4XEaJEVrIR1wrgzfplANf54PICpgwzHgT8
M6f/u5jocH+SOzfimgpThnQBPH0SpSgvrH7XWU5Yo/ieAtiUKFo/Wb/VVcFEdKcDqeUUpUFXK0wn
ddSiPt9eblbD8Kg1NoddB+s0mUq5+9kp6hF6sjyP+RtraYUEaiLI/X3TVI0gVBPBbfpXUyPKbgf3
czoI3q/tvMRGcMLASGp+f60zs2dBrlKafielVW99GD6s3qLaPyAmw+GaOfi7szxHf7iy7oFk1Jf8
vZnfvj+wb+0lpYXcBH8yjRl3R/MxbZVzS7n07zTlOfV0t3MPSNagcwVNoXvpoif607LYboyOi1aH
TjvSIPAe78VPqXab6qNaHuf0scbgsHQ2OE723v2yaorknOKUssO4S4xfikR2tvDXS0YMuCPXD7Ai
JQvIY94+AyU6APxm6uMeQvD0kxjNLc2ujfcXFcZYfX2uCgVIKCafFeu6ecj2vKZiGPJyGngg4k5A
hF1TqipbW2REpxGf8arWo5Dp95/MdTdw5jONg3WhSnSsl9I37IWy4fyqyb7aCtP73DgQgagXs2dc
iaGNrIDcK926MpfUnfp94OkT8W2JsQ1qJAYqgycVpoQ4ikC/4XsgDb+PnyY9xmrVchv5XDE6/X6T
78rW/NPcT5IwifPn/vcEkOIIn0JWH1rCeJYttbGQELzSiOops3ZOEfm3NvzP58yxBB+IatzhVUcZ
U/hC4ftWGsEntxhv44t+8tbhOUdqFTMgo4RZQToIP8J/GOcmp6FSEHfPRMIhPO07iCnMFtS32JLP
6uO83aB5phnDYBvkJqCVjJmjA3FgULsuUvuUjytfDqjdVRHrYxpgs5kSg/knWstIInIRLCFZPX3s
bgsSYMHQqtagXUH3vlLyHew2pelYtX68WYi67L4eVYouARZokDW/BlhuDPorQXu9ZC3c7yLCJNvM
OGNkMU3YmiMIsv5Q1UQnmMuhceO1BdZ6XeN6y/tqu6ChFYFZNXkGU08Jx0HATBbvxYqB9DrcuCX4
OeCJ/zRfXEG2s7sJlMQz2A55CQCgFxlz7zwQbeyCZyloawizZD4tSqHCqiqTd2FTi6hOuV4MLFsH
a5h2Q7e63iVWTvIeFQepA9tC46UATZgnC1WVy34KlleBvdnIp2Khk/ixFgQw4UNCllPL1a4pZJDW
TGuGcyF7C/3zNOnTXruGuVFFPzhb3a8+qevwaNA1jcD4LAhp6d6AtGFZkFxeIqd5Z6VDD6wSEzXw
g2ZBZd8AL27ow640OF5beYd1CdOYN/ay51Oo/Fo4chRJAjrowkA2ZM241W+OENzj+BDETKLGNsOT
u6e4xpGY4RIsPn/3ukRIv5HJz2OaeLeFj/KECufrq13dUuXBmZYTuu4myzw+ChxfXncFqFi/b8ZC
ooW9P86EtUwrRdQevcniamFoexHQXR55bjpSS93+ygKSwiQUviZLGQV0SKcXKP97ad0YMrBXnzUl
UM8v37FnSGMS11/KlvH7VNfJG8AB3pLTC0VZNfiIgdXD2GxbhIWwMCnIEhioFRo2EhBkYVWOC3Iv
qKiP5GmvPwzFjMPsSd0O34TyPq0PJASJDYTDDYPCDDZmo9889sMJDA7YrmXoZi7qimbP/PMVU1/h
pyy6nNFFOfu9Q/XwobdaEPKdS1yVLPS2rCDdUCJghFmCFdxtoGg0gea5x2p3RQ590mIriZ69AAXS
GSKHYRUhvX/FFlQ/BwvVE0S5JyXt+HOKaeLhI7o9NPW0tTHSlaCwj5TlZQ1ub8AvscSH8lHkGePp
ggth+Xzpq468Qdxch4CQxu8q/Yyf2D8f+WpD/rYuBmbaLP4VClRCxjkIScnXaT591v/+DmLqZsOe
QO5ZcpUR0B0pufYFrbbGEvBThWjucu1lT7pnCVi4Bk4bPH+YWL96W1+mM6Xa7uXPL4sL80ihSL5R
prLn/yQ93MT0LorALFna6wYHontEjIsmvvPDhOuMyPPDWdrg6fF+c28Q0FvQc8D8uZ3fon0yJz4c
a3pMa3xR7+D9WYeo6Uca/6/UrZJmnFmoPtn5AjpFtwxSvFSWvUDInULWDDVOZEmDEaokxUc5y4fS
IvONBDO68I89Pq46Q6hCVHZH1p79jdKiklBNxMZqIgW2S0zoyyypUNvs96xsiMeRa1eDQB5DJ17Z
wIdiUMpwaXhlS1J73yWKXqJudVtOn7kvy0FCAWvdRj6Oy5CKjBUpiV+0DqEuAb4sSc10OnxRTjKh
g4NMouYNXnqjKLLohqzlINEQevPoYezkj8dZtX44P1Zqg/L/3Xgkq4PXHaukYDXq978CJ8RNozhg
OH86dtq6vPwwSeDwni1KZktSuBvcxFNPhmhtP6HHAvROXAibl6NpiIChXOJ4io9eKRBbP6reQI50
8ge2DE23liZcxdiGI8J9UoMeRQN7qRvCyqmiA0Ohk7CmqNfL0+U8Uuv6RfvTtdUcsEdF7Hwi1sFq
wpaLTR73VWoL0Qm3602FLh7HzjH3nW8vlUC0zL0WL+I23UBqzcYwelkc+Z2OyTvraOv7/WJVVhjU
JydDKe8087Jxk9c1chZzWTfeYVDZmti/dmMK3tQhoU+rgMYOMcJ2gjxH1PBtkDzdyR3IpthJJ+PB
st+eWXZV7shtzn/J6zMmsxi9oNeJFAqXMjvJUajnPDd5lRFUpxIE5zRXHWFFUB1wvmw3m8wUv7S9
jgi80M1U60LTUTlDscKr5iqD0WjHZQrIBu5Mj5cXIapN11F/VUkJ59kME/wcX3tGtXCbrVCJHaMW
W0mCLV5sVbEr1ONIHyz5lLrQjFMZsQjn25ENqmCy5jriyVrUvjEYXW6OtlnJlAZGbJAuUdxLLTzN
Q6q0RnbjOKh7ncgJurahO3NfCxqDe88wWx3vbxTfVVZ5C5qmGaRg8+qkghvsGqvE7Y6h0Ub9AcFk
K46g4a3bWy4UkCPPjumgTxMPQHuYm2TNi4fWU99OBWwlxVGUoJ3HADY2ffuENYRfwdBwfJocTo1/
wazKMNvquP1r66ujcZPgUXlYXztM//HLY3GZsM6RXJBntuQZAzlFTiXdMYhPXGdC8M14lTsBI3hm
2ExhpX2Y0E2LfkZ9RmO4BA7g8Hn+RF9khv611DNj9emZpb239O4JjjlzHRnWNJEPc7fiAYn1Urz0
mOCv51gKiYayA1QKy7gVzgNp/V+heJLruWDeYLun+OHIrgpWG1kkz2jm0UriJBwnJDvysu4tUGVI
3fuyJwBqTotiMPmhBOIYGKHI9zte3t9FFAsdsQ31aGA6ajsVcIIyD0QLHXE0EoyOd7AbeW9xWYbK
0lwru3BaDq6JiJrmvu9H6Mi4WDczN5UY56iMCX8t01dnBBnhZYL8Zud/B6FSHSN48UeMM+xq4RW8
2I/v9gutwPmBZVztGLEarQt15np0bfOmQd4H2lUDhBcwIiqd2fbmHm193e5e5xc/Xqqw+pURFEkh
80bAY4b6vLFTjUQA2/QbHeetVH+stb/VjN1QxhyfKHW0ximteju9yrTNdH7gsDuCqqBXv3FvOdH5
3Ah+/ij/FvtcdEyGMuNH6ryAJ6Z8oMfh2EdPY9sQ4N0AMJnX99IN6GeLmGo4zn4a2jN6kgXH/lcJ
VanWT8YJR+j2Xoe7U4rTY3ogsrWSqgTVhYc56dqvLwqiWoHq5vNKhU/NQXqjXi/UxWhC6m5dNFHO
dbB5W7BBJqtT7amWF6voprDCLs92S5V7UvrYofud0yFZtG8HQb3LqkWdO3j2fpHGp6qcbnZIa/ty
ENsBJ9FMPDT2ey0nwuaWUhMkkw0nEoZryXfGDl4twg5oCmsxT+fCL+dEj83HAL+TcP6K5nJqvlHl
8zB7uMsFX5/XuujnBLlnQeWrtIG0LSSbiG+rarZuhnYllNiURPCrP++/LGkLZq3v1yTA1T7o6H/i
JhOyk1soTd+hkImaLXHAjanw+GLfUJyVjf9coVJEBkMsPxBxtX6V4dq+MKV02DAGqlKjTqCIM4ET
8ynS0laeA38pJLnrmFR6dydxiUzkk2MEILuGyZC2STNum0ERcmy8/FRYIf6VABXYatC9PdC8nFpb
Om+9mJCVRdllgNWNSjcVpNfN/8BYQzhNB0jAMzbHx866qXTRtJ9+5h6Q6r9AfXGlc1msz8I+sNYF
LmLzPk9+CK9RJk0akJi0qENw89FNH6yutWoHuvNLVlk59IXr2u03Qmsdx39sWhChGbKiIV5Yye4U
NsH0tS18EoYVzMXIyRUlfjxGl8BIkspGajVbMehUPCaMssM6oPbnI5H9af1UkYkts4hzVKQkAgfx
LgWdoYRRBcnR7XpG+0ecWYgA/Y6ydIDd5vghPCpVZhbyU4odb5H3lQM0qYsh0+skXg5HZN6PWNxT
/cP09vMK7DzMrewffz29iaTYQpaezDMP5FOvIziPLo958GAnMtNIC/vsYKugo37Yh1yRrSXJtm88
JJzIR+n+ADkUMQk7xZ6qvV7R/Y76hvXFpZB/FGNf4Sm356Ddv13JtvSAUYE87E0YKya5s1OlQhDF
5o6LTxq9knULrLxdhLTZRvxYN718lciGGHJ9rXKYZNuAgJgrKuqRQaz3w9veo580Q061foXpsoxz
IastCwM7xZD9jWwI7QzBkQa2dqpgQ7iO3GdvD7vQimfXLITB63iG35/ZZVa/fVGtVQMf71oiFgVe
TiA18+hyheLaJZblCo54YbPCE1/pSi/vz+T0XRQrIwsxvkG/T3X+GQHkTF779p+TOwY59AZGRmr8
prj9xkWu3iGbOdXClTm0yt5+P78UsOYwKijSFXPm6BtxxSIxDkX/K8V2mouqZNHMAgIAn1u9q6lV
a2tKKL4LfV9FbAKhGOBGIyiyCKDLDuXIi7A7em070h+3eZHS5WqM5hO3HZG7IXfTAuOMR3+Heb7q
rpPw2mw50xHsZdS3PA/osiCvp4xOFOHwgM4wifEMumqw5MhTSm2Ryg09DEwfq0mg3MeUjbrZzxjb
BvKm7izfiN0hiKGSeaJ2fCveDp5BpMmK6UKMBUYzB7GwjWQGANZIT9XravxTfAgXKV1t5DBR9hlY
8kMUOLzCjwxEo84DRJNISE9YXfNwF6Q25zsqxmDSl/Mu4vx2WRW1tVDVWxbPN4MUFttiCYNqb1ug
rYjPwtLuc9aY7Z3VyujItPCj08BgpdtC28LxZu/w9rzl28TLqM1jQvVZhjtFMeXRlR13Ssy2naKW
Zl+2b36g1nmGBX9LXyk7QoDBAc/GVyzTI12ovzRnsD2GECICSHK+FHtxGXq+qI9XjJ+g8tBoNgPM
OVyqzzHg6uMBcASihz7L1e9zvo8AWB2ZMGrpyknjURmbigGwtGrOgy8XYW5WA+fqhs9SayYWsDB6
HLUt0P6q7T/Tz/xKuf142+1lpbbhc5BiQcBWJ/HLrWkphj7abtFkS00axf2FXcXSkzn2Sg6yIySp
W7w+xuXz6JIf3po9tem3WdqY9yVgT5tnqJ6bJ9TzqeZVELI+CEjL6wh2JoCxpk3IdiBIwiFZ26L6
qaGSp3qIqNG3tmqTu0IqjTQ+yyaohLT/kCwwCC/Jdwm0j/B5xmbjsNWlqqiMcWq9+Bv/oOk8psAo
0+HRS4j0P3JfgV8+T5eLwHiwYeVimC5CDFATrnPoKZSqL5insWkHJydzCrA7p/iBTFLAe1RlhdOg
kgWi5CAmeHBy5f1d43Clx/LPCjPFA4L80YUtuST281g2O0u4YDGvhj4xaDZUiDwEsgti8mpgrwTp
OxNUAhGF7vjfX75v6oWE5XUx7de1QFppytUZZg05V0+yiBHZbnXpCFhMyv2SNsIULxW43V6mh5/i
tkUr29jhYgG5aSSjutX3L+U1CJCvagw4po9SoUCq4ijCLtYxDNJjYuy60RvjCCwCMphZ8XZJ03Dt
pS2XvaYSXtYaJ1bYLK6shvJurAdDJ+UpjmR4YB066nAiByOK4QnEE6JyMvQ963WupcpI/NVD+roL
3e6/JlINWXhWCj91BvLbPOjRQwTLQTB0/zm5wKvtwZflTsT02b7qBlxeFDq/A8X3kdq4CRDPHaem
Bh5wvo/UbSGDzUXDrR3jcW//wcfu6EAsJtDC0/SoywFjDXk1BfbrCmMz9aHw2AD1svG20qEZg4Y3
apLHP3pfTC2muwuujjBBQ7OgWt1W3clrbkQlDY+uaqICGFtv/+aGcS59ZN5leqTv+TXp0M5wgvvc
dLEzABgnXpnhiX3uO0N8jJjDxqWOe1rfCMSETkAFnGigVI5n63ETrzSrrGO5mb5DBRRn+Xuayn7n
Zdmrie70D1klVU8nXR+6URYj13cdh2DqFzGcd8jf0CBySNwrmJl3ycOhkxzsat6mMty9AKyWiaBZ
5F198/PdNiFgIJR7gza4iATe5yxjeZWi1fArZLyoPFy35qbJCPT04XVk7BV3KdrXk14hAtqfkjXI
orSuBATZb6w4XFRIh/TOdeWspYvQSB33iW7jUVQZBA02MevCx+rc9rBSSNnHl1Us41Ub2egiyI+y
sZbUpQ1aKSYVpTV1/5eclXZl7hjazBQBcEglt6j6wVu5oG4hl1VK8f6y+LkiifT83V6AdZ6TLavN
fXWgGjU1Zty33NTjLutNaL0Flcd3JXmdoeYyzdL9vFI0+fNu5xC0A/X1MWTi16CHHzUc3sKfzDz3
GBiSIqcY6sfwjz7FaudzzAIvw5QCaSAvx0hzuSThbn5CfvMLtPuAGEzYi3/pgVwBoTNYr1YU3J3O
m2MsVh2l8ZT1Sxzg9uEnK41H/DOj0LZVrkpI5SR8Et/p7gAH9HSiUUU4rMQeWj4luiCPc+SfIezZ
xdJBCo84E2/so0qAdIj4nVQxx8ZxWFH8WsrZYqsZyFjxh1BICHEi4ClifKf95Q+9q/ytq9panmig
FOC2OD0i23OE5PK7rxLNd6kzPBbuc+rr26ND020FsZ41ddyQnq4Z/WRmmJ1Hkow1d6DhPFf42rsO
55IYMK4Oq6uawwIfm3W14KBboZ9rskEoF2FaQCt2ex1JXHhC1iep6k124biJEgYbLd+SnpjV5ugt
6qjubmtc9xdkWX9oQI0pCY2gSGKcWFxuU0DUAk8QYTgvpsghzJPcmUDDaIGWZxOkx5PneDIelMta
jgDp2CLxJt3JbcIZeslY3N/sNorSsWk1JsDhypFO/0XBwnBqP389sqgZ9e5gAsTJaJy0ERtDNGd3
eI79hypUlw6hBTYonNf+OGl+KQ5hhKLWbq0SPgsLfcu6nm8F3KcSiB4neQgg4yd9DPRZrfHxSe4S
JoywrLkw2HkeT8bt9qDv5CHzFIXm0k/DItoKi7115dGGVIokz0rT9XN7kWORKJGPzOnIGxcE0cqa
nfB0BtGkAZZfEP4K9se9UWoE2ZrSXXSgg1lxUhNH4/jJKQWyCARHjxPSno/q/BE+yDCJhh+RQBRr
MPaV6pEGLaMBRkLnB2ic2YWU0eH/2NPX90nT0cIVEirOviSZpxbopI4nQHOukmCx+VrlXPxDYqVk
/+t7SUUtr4um84ippt5DvYoWS0GaYkpiNbHs8tdcxxppjmNdOVKaUT+zNCIRQ43NW3Yc3jBQgvPm
A1+Tx93nlpAQGHuQZQvgPYdoMEzCsmTnrkItDwc0R9ANX7WCSCWtLAbjlm8OU8XYOYYHQF/Wiczn
8nBRD1UlD3/opfN0cbF/GPNhukOKHaPUPFWdzuqaBXGKvJqw6ZmBcnbt/XL0su0RLYgViixwgH6E
B05i5I4hKvpty9U3nQLKdq4w5Wv+BQh5Vc4k2JL6QNwswMUOW/8k8bRKOzWSucXVkgra/EfQD6WY
Pu5vmGPZ6VtqbFnUuViG4G8MTZXAC7AwGx+vPe+VhPMsJlKG8QSXMcduAM6QlAWHF/TJQ5JVU93G
bstZt2X2rycmVp/UaYHW+3Y9X+zgJc+VYJWxXytK9MFa8A/s3bpr/1gp8CXToockTaw7lLMNhW0W
8dbhYKOHOUaipQt0p2PuNBaKd28/ITe5CqpNMyqr4Ecy6jrSoqpX2RqdOWYupezrIokcvXAupvLd
VWUyDavZ1LCF1L3sH6dgxzlUmDFIZm9/robkgGM2yTKJlpvwfczbmgK3hs7x/+jVfn+93w0Iu+Ua
yhTBrUVMieASS3JMVPcofF1kJh7YvoeFIylO6rBL2pebb5UfO/Sp7jki7cRihHpH6/gtvx4LpcHf
gKS3KVYm87JxbDsWO6Q6RNQLU5C8ODrdFcJbQxO7/bnsRkFSqQl0MNeypM2QQhDhyeCIF+9zUv4T
vr3oWhTx1L8ad2zzcwrrxrB5cc5E19dP0o310yLWG0O02qXhVv5L1weKLsxhtWDRne2kMeRda+W5
LzRHYA+AmY50gGEFoMrZuovp5Cl6DwcA/SiMuPewl4AH+shdHE4gvWyPOdc1iOhIFQnYxylHIVf6
LATri9JbYItrVbl70PveatR582oQnTZ1tM8sxF3KH+Y8O1XzgXm4mME8Gz6tJxFxBc0T1GtMqc/Q
YF7qMRdPqvZCkbfHu56sAKyYogELqGWP75iPOo58kBQRc7+1Q1XMuqEjo2HdXN7iw/68VscNwoLr
FgzK1CsKc1hkY+m11BvXNn7VRTKkumN7lKHVhLO8GpK9v9sRqkiPOfn8ioOMMhB/Mw2cWUAtEIDn
EIfaRCIRKe8DZ9iZhXciuSgQXdOQzso12kheb3z3lQiKlpnINPkwlSUvb5Rz16g+JVckfCzTaNe1
uY1RbShzuVggoAnX2r3aXgI+Sfjo2rj8/3hkOCyFtf5JK6DsFleaTgdAxKYHy3xJOk68HF4kad6X
LZBt7FLiK3nC0oo91OJnVx717kRbnp4WuuYpjPOJwwl/4fGXpsdf976k379WG+8lwxGAkxda6Ymu
aYNRsTNEED0aeEw92+o/cOKnKXaGVM+0b2SXrb0C94Monw0YrwlQl+o5xHBMxHWd6hWfj98nbGP2
AjSUyNht3M6Yx8U6QU75J1r7Y7md7IJCe7B7oljvxEQ6BruOpu4ztF4tGo1iR8c04wQcNAVBgGiY
GSQoeBhRjvBNOnmvwBkb+fDccpAqYNStIjVlsAkdUX74adeUh8wPhYLCqJvRg1Xwko6kKjN48Eka
ZCLsn+UuQ0Ue5a+iE2UKLHluXbjxxxwjcMJQZ+x4Gu+XCTDXdhrrS2JSjAnTsFeIP6qbfBOIExR2
zGrL1KHr++wuClZ90rJPhvLec1tu7NfgbvM4zFN4FYr2BA+FLm5WlClXndI94DUs2QKPQQwRS898
X8GR1G62c+vl1Fm8fwkZ0JvA8TMrNQC7UrB70sy0tJPCHmHM05nf0Ke7qOQw+7G1ySZq0c+Vm39V
tA7lywP3FV9Zwj4drVfDm/pwPjAhE0kgqqua0PtarOeWmeUialz7AHF8VkvCIjNxzJTcGiihPRsx
1jNyf86vWCPJvYZAZkptP+gF2n/MQ5OiyXCzZ0jsD0qzThmJ2fiUZFdHCS9yazgOJfDzBn1vsnhc
PgB1Z7jgGFRK1drGCz2PIw2Rn53bh3E4aGvFw2IwZKtGmiILZvMP8/gSQ93OGqlB9HrJxexZ3tk7
bSPlG8nDTmfWxT6g+O4JO5fSNxT955vR6EhQCTDDYK2zjnPMHRoFdSbQZ2j+tpTEIfA7GFLCxW14
MkPESDTyTEpLT937AUa75hcXBcXor75Fy54aL+g/WNIqNLHiVssmzbExlyeaKa+6qP04no4Wd2Rs
NMm0/0E0klsDAuisGVUHPmY8SKmgnrWz8qle9kK1rxFqMQ/NGDbL8vxAygXILXP/H9707Kd7MpgF
MS1h+/XEG24QX0f1omppikDVbP+tKdRmogPRyB8efMM0WslxsaAJH4614h+FSk3N1VKr1ii1JT53
iUilL5jciCa7oeWV0GVdNgbN13I7IkIfFklqK8r0iTuuCF/T12+8KlHbyV62ReYJHUhX4q2/mNne
U/pTOS0ihfK9o28G9jVZ15vQNSrO+ZXaQAwbLl21yWFfk8x9Vj83K83NsLJ+B87/UiMzlPE/Dq+o
Brk+FGjGrCz1R/GGitMiySuw5/GNfyh8TrEb9a2md8d2eRdJn9xr0jdJ3dIl8zf+H7rOFSxULv6N
o4ZS3upftv9XD8x9sbAr6av7l+H0WNGUO7UlzN8z+zr0EU7Zhj8WZ9Rztq9Rdh6J+RhrAtIRCBpX
B2+a5XaH2MJTt4/XMwFJ8AOdlIFuZ3fJnu4naMfq2L9k6Ucfv5k1SzohP7sLMKBqpya/IYREKG3A
P+dq9Zqn7g6gr+ibB+kJW6I5o+dFhzWnOjF/20anD5BnytdVscTR8+lWWpHp+EqCjs5iIv6FFyhf
iYworufIoF8Wu8NxqJNtJn/hAgDp0lXwEQ4ywKK1j2s7SVfuAnATi+Rnj25v1QQcdtXc9RqYlx2G
uG19feSoiNc+pP0X5VT45lKdS3keHhLKU8y7kRp3LsN/jjjP6O3bhwn67YS/gd4vg0zjMdhUTgF4
7CZgIJE04MtubZiLGnfoqdVYU8WZboGVi70oNO1KtUwwqrIWDJROpOI6DjMLeqCaM+VvYblRaQpX
Eyi2hHVk4KUCGdCHMhuvQFSQ5gfgkkR+XjrM6CAyGSIHxJWeNp5lGIOHE27q6Wv94xDRys0aTepO
+SLPBG7TfdFkdJV1bjODxeMIWUgbSmNuunvgs7dtKfFdEbfT2NsGe3JlzAx5i/FM5rj8vlYR9E1f
FuA9GVWYIgATNrXpkp4i/QuTEyAxCnAXc3D74PNgFFWzO1bzVqyyRtyWXr0MOhEElZSxU7MGIT0W
86bnnkzAALThR6YTczf2J6iqOZ0CQlRDqKQn4eqcn9HBnDIo/VnspdJFeK8cXgHUTTLeSkKcg1tI
wiqIwyH3nTW6aYhRAfltm8O37kszy0pA6+tBrvQGklJfug4mXRPJ8R4pt1pUgfhauArKPydZnOPq
gHgtvPQaTE8DxNu/on/zVJDxhKt1azi4fCNzw4UKaLGgRCFlkxhExTMqwH8BuXCIvCFZnRyJvnhK
2tCVS+cKgce9BJZS0UPn4qeFAg10akdV4p4dnZiugdFB+5wUEF5LUKce6AlSqKKllHuwxR0i5i/4
d0ov79eTc/JhSVZElULKyIhXDC1XTion5ni/Nc2WWK3IvFx5axUYAAFcUkcA74+mpkuiU8fKQSop
scw220TsxdqpGgyjFY8i4Mi73n/JnMS4YXopy9z6JufxSD4x48yI9GgnsLv0lkXCuiTbCfsma6fb
NHX9TgKeqpzHYW6W2mOyy67sSq3Q6W+yqj9Qts7aDSf8KRE0/tphSj8BHH4QMCOYxiCHoMF0OdhZ
Dg0M2a0jiNK33XOduGMA/SS94HoCt2SP5bjDKEFltg9XlYahqYqt5YNmPHm7X71iK1MvyM084pak
6kA6i6zotvD239bRkwxiZdcIoggyltdah0ZsWD+FD9p6YvYI70WCcwewh6nuPYkn4TC6V8+xLLjt
PAjSbUcBAOGahJTT6Peku5qFsnZaZdkruYJG2JKeWvJeWACHKFrUPOr65/BOx2Lzf0exGRtNsSJf
HRE+UuRc6vZTzthjDrXr5wMY55swpP4v5y6QnglHNpDf34D8i674LdepXWtSVeiLf+YGUOnT5uZR
X5sbBhtC4r3Sxt2CrtX/dq7g9mnDwf93BrlDWQNOBiLMaAzbh/MnxaS41QQSJxlAnv2lI3ot2mKn
luU3911+F21PYo7708lkF+LgibVefCISUjMAhtp5fjjiU29EGv4w1cdFJJZ7r8gCR99eAaqSRICJ
FXi0b3IybLIKrOk71+Vzlzix6QjtMH/9NiQ2SdQOGfTWeQvmRa3cXb7SHAV2f0H8/hMASqnUoMBH
qpzYH30jMMl8V4zk1xVFXIBFHHQ8Qk5QcWQa+NargX79EBVJGp/iu3bW0VwWqUna4V7VdkaX7dOk
nUwF2OwvoeFCasS1ynsJJFod872kDJFbnyRiLgoaDjikbmR1u5K5UlAHOMmBTXiHsnnrR8iBWfb5
JSZCf3kz/tJMipbUJ8ZnFtSdpcDka9Mu4nWIAT0i8ej6ob7pyHj6TLFXQ+Pmm9m9O0eYGTJlOa3m
SRn7O8qKX1KwB2v7m4BdunWPuOV3UoXcTWrPjYcVVz43aL6OAJSUF4ogsidgnkDIfBtUhZeUWCij
D/8hCJiDkn6OsrjdQ/9IsR5B7OQmFCIcOmmNC+0yiMtBBi53mMReH5p8kcSCNGoLL4HcQl9P8YQi
wGzX/JRCVgAJx9hmZmexQPcAqK2zXtX7iCYWj6heDMNpDVyFX12HsGpZUZW8R0u2XLmgoMIKU8ZN
xjbUnpxVEJ3REaKZRwH+PhsfYT3ApA1HzHV4coBVJHfRAN7oTV8GYljgS11d3Qyg+ESDZmkmpODG
VBqgZAaynoNBiAE8sRuLYVa7RccshdkzU35W8ZC9OaR/JncxfMV7NHrCFfImAx7F8U+vrPQbtZCT
8I+Nduv+lQpbQyjINPc8NlKiYA6NILgIe0bx+yCPSbkUOc1vi5FNnLaqSv8wqtNQLvTuJ007knDq
5s6Zhivn8go+UvfMCei26W1l+8MUzfFwrPvOHR9MAF1/beV6eX7+25Rv7TTWxlTP2dXTjLxI5RMv
/wmxvdhukYSEL0wsFnFMb2hNDjIZRy61VQj7gFZccdmuiX4ZVt54iDlyMxPrivy9K7gjdRhtTkqd
l1eFbXWUeHphoLnonf3hz01Pb6foAHt9Rm2LDolcsc+f/Lq+CdVPZNpEzhNnn4s18C0Rt9xestav
hOeorgUGzvdTcPXmURjrNBLkMdvdyZgbVbLsJamwHTZqsm6t1CaGR7JoRzgGPXj8t8dpq0LEJISq
nWGhVXD3PxmP9zl4aMi+onap2Ra8W3YgDf9ozhKIADfLbzFoAiziEgbDum+cp/A+sldYVsBhrkXs
Y6zKhAgfddeJQYOCRPjEyhxejcX9vmoYCZpOlUo5oGmEYDdmjzmLJxkaeh4UDfQ0qGhgmv3/grE7
QhQVfu0itQ0tuzeRCAOumwrhwCEBcAqHCL+fQGIVZbKuCoCEq4sMvKVB58nrcJkitCo5hSyRRbDV
rGIepEP6AsXuUj6ameesp1AohDUd3dpcebUou+7tFUKfXSTYi6tJ03RWMDGgrW8TknvSDViFYdvX
nCxkxri1JHDTKtvrT8rPpneWdlqJNMD8NBDsI6XAkHJ+DikTFjMnEYU5EJGlZxwgtlHFTE3h+CvF
B3W1hbNneh//saFMoglKSUdvSYIDV3rqYLlAA/iBcx94nh5jKaKIDLT3W+3vCsg9bDvg2CTvWYwn
9Ppg4hYxZQgHGTGDpKtl3QFCvRRi/ugQopMA6tGrYSPPHTTjtKPoE6agamKurhpgjJI9agr0Bt2f
Ww+8nC08CI1Xq04hrAHDT5ii8KHrEvOChehywArOa1QanPjoIpUrHxvy2xfKVAU2UqaR1zdGzFX0
WSs1nbS2i2lhUiBzwBkme9GoAGs+ZtZ2+S4YPEWH6FlyYdpXq4oZ35L4cIWFgii8+0faom/UkRGE
QxKjkUqrJ9n8TcEUpsOGREFM9RFB31iEcPFhj9zkXeddENCtnrkltIdA83lz+TX84Z9FZkZhFrEY
ihdS8GS1Wa8J5c2uWiApoyHz8RheNV43q6PxHgWVPbHd+OK3/pdIxTQp6/2j4qfwowShsfypticp
o1rDsKJNLPdv9Jp6hHRdP94ES/GzahQkkoyXp8ZSZMeIqG/2w7yXkpvB87gBRh32Fl9NYoYxjhrJ
VtOVH491ykkGOH+E18jUqzYsRHRbRbTwValDD0DUxvQcc/2HAzcc1YBUXFkinKbWsacq1ITCl9Xs
yR1njXzSTXjwpW1hYIAttnNFTCBZLRZn/jjLlJzyhMYcCNaoOMdQwRAtOQMDj+vEEAOuzOgirrWz
GCbdAO2qDLuqETw4KPdNx0bJ+lqbuKdkA3vbU4rQK4eu/043a4tVou56AklCIwxlHRh1rH+vLKag
/ztoxpTiba6rD4gvTVNM0crDz6Q5O7JqCcqGYGBpThqCaA2WRCFyOJxAnQHNDnDJMs0dkwuTRthp
ilR1c1ogoz2CBVkj6ROUyJUWK7JfWhdpHW68WRI8EtdpUbpMBZxHRApqu09B+QnALJz9UEY9xCYX
EA6WAtrG0UaKF15aVXj8sE6iW1nCtu7dCQ8sIW0lQf46VrGDCh0zco+ymQIhbRBmortLMQv1JMZx
jvkzE87G80AjnUgtFZrdKuLYJfUOdbR/F4u4x8VnHu+RrYT78rB4l7Q5J0fRNsHSj3Y1ub5MSz+3
8uMRkTW5JPkOCS+W2e1yv/zWdh5M0k9nVYRB/DUOiVJT7vvBNdGQt7YcdlUta8JVXNJti2tP97eQ
EehdwZJuRI7ePvRYemK75N87ndO5B30A6ng3T0qG9GbVDFF+uqC0djAF4d50Q8K8pRmRBO64v5lU
N4RoGAx3Uq+7/As7JJJFN37DPDVojKj9eSjGL2nKbMTNWb+ZNXtHz3ck9Xg1xXt6zGMo7rCuwrPx
6kYhSJbq9fp1TAGKARqmxbWc+BFO0MdMMBFPl+ZTLkAfpwEzTM7vlgR7jgzULoXzuXfDutSFzDQs
PJaXd2baZ99UvOLyNSFY0z/OZTR8BEeZsQ/jrclc+w6M82lR3MzwwlZTcQhtAAsr8qL+qlplpu8C
MVIX10OtaCCfg6mHFRvcOL3E3aclS0y8qFS9jxvhRob7Ff+JfUtW5kOAJKtAGHRDwcesMrkk69gX
QREclqQSBUlGo05x1w6CbT+j9Nk8lu5LZeLs+I1jXqC91EmL0en9KXyaUBKEzMdOIFhA97+oZlGJ
7B3/TcxUuQ4EA3r7cGI4bGXZ2EnOKzn0JD5847B+CFZSiELWCWj+yIWPxsPMZ129t1AzPwIKt2hl
GIy8POlHP6ORbztsyBLSmCqjL6b6QfmRFOjneizquI5HIxGDqYlYcZeamTnICMl766a/Nn/3okhq
5BYIw5FFAPGnlId26e2roWPmTSbRk4D4UjCbnThTC2knsz9Wh66hdJgiT71XDJlknPHdVBu8dqqD
tLBCam5VQM/HSf8ni9cutGfkxpeTK0LJRjwZgYXkoqz5a9FmqIHlS19Gx5hW4RmPdrIKyiYA7quh
LYLHi7s90cJHdKsSmp+TaEsJtHeEgReP64O0Fn8nbD0g8R7aOkCh3EBoSGIdROZZZHNgUWZxFxEK
mofvdJpS9MjMQ4GU7Cf2bmSz2tQ5iXQHwq9LLxN9ZtjEboCMK7M2R8q8AXubVLdVtmatRU1POsFT
+Ejdus4tNwubWkLUlBH1tlID5HnhE4l97fr3rI9wIlLc/7sfqs0l1POv6QmH01oRMyaMHTSjvymf
mhpxZmTOpzYBNfNqaLJE51Z4AzsS/iKQr5pEDpBRaGKHTb39zcWkE41XBEyn12xrajMIiH/VRg0z
MTkzWJjJvA+ZKrdGkL/ZygNwlTkxmolLAS0g1cc8eI8OSHPDogOsLCx6+4Zm2zfEsFuIEsmMRAsV
cB6YhFLDitfLm2dK8lvYRR4767gtp4KU015lWxQYm0KP94G8m5yr8vLv53S6rUw3Tw4vKoa2w/mX
Xkat9S16cZuf/JVuKhonFU1gyPa5qKIB2dQnZiPRcU9eK2bx9UoZtoaflXe2VnRnVI2UazsG5oN6
UXD/T3i7c5L3yMV/XYPsHp3zM3uQMGFbikTAP1mmaiaFN3kQZZ3Z8XfkYKXNa2alj6/H0HE/xoVj
6St/wl81ZLJLVoJQvoC9tnOK/13CRSFbicbfH8lC0qX5yX+8P1/RohZ1MLqoNnGAB96T2HjP94Sl
6dLjKJde1M9CbBsjJU309xKwlS9paj2mYtwQM+Xb1QKdW61P9+avxhFzPAPxNCbfAPb4jzbcHzm5
Xy7y+75bZnCyuMjbcrCekTlzr5HAXW8s3jM2MRM0W74R50D3tLf5c/ZJofqvOGv3pEPL+Nn0SEpt
5kyMsy+KZXNIYTvkrxCV3SbP8rFfb2+bzQdmWVgVuXSDn9JmybL1R2UK0cRrh+E+arf/ANhYRLTk
X/OT+ly6eFFQqGCXakpzY1RbgO/xXT0CjfmUMxqitBPPSZO7tmSMDgviSFNkjbhF3qrvcesbyugq
+a8uhWkO1sjTVi3XW4jkg909MOlPyZo24+85VFv+DG2/ASoJHLeJ0NrvdbCGG/KGDUAuSaWjPNFd
/BBno8F37wzct36yUixzJxtl0HISKFjzc1bTdWCFs2MmDdjS21ScQJH7nuVuBi0ePJc3vAKmZ2Hl
BK394e4HWbMT/aL0Wr9Z3J13EPTeYNTTUQ4H0v5Ch4620Y9A1HwYz0mnsZn4yjuti5NxaHwQxWv6
RcwnF3scnTAmXQRCEcSiVWJ92XXAY7+Ar6r5z4S2qF8tg5e4V/z/IKzIM8mgDwn1oDFzqeiDgzMW
IbOq24AYidW6ryA+Tc+HZhvGFvm8YmVC70TSlSjdIPFfK6VV8Q4vE03Ish4bbZVanRT4Cwh1c7AI
vcp/e7HYWpPdn1KAbXSc5FoYBl6UiUuwYVnqsxnaanjpwzir0wFRvh4Ub0ewE0MAqoEoYG+e8rw0
dg1Vaz0VWHIyhQn/i3Xl/qw2EuVW/K28e46LYashX3op99mxwdXjhY9PGCom+fXe3WCalr/5T6L3
zG7N+Xjvlei4BAitR2q1ZIAemQ6HrO3vNF+U7YSLW7asLW4yWOh+D9bqOUULV+XzSkl4ugcc6Qtm
gFOp3+umR4VmqANKtgOZ2NEF6A3eNtaP6/nTthiQqWMZUzo8BSB+f17eNbTl82IP8HoRkcjl8Ev3
sIMSyqWWlfpGOgc+HHN65SUvDTWzl6FpGa+M8kdKAsftIcEEFfP55E5ek+5UCb4lE8qOtKVt5Hlp
+XLGiiSfl1QJTYQ57CyVmnzHFTAaedsf7d/y0zBGGxxJAyYsRI3Nw2witOdNDiQkKLcEcX/2WZdb
uVPj5G+O9P3JG8WStUjUI7Is8cCDhwztsrsBBEmPfaU84NjYT3jwWDe4wo54U9wT9eFKi3XqSYZw
f0fjGs89U7iQZRZieUbulLFr5WmAUfDxbqThlDrAZFb+5Z54NBIsEG+4oKbJgElpIGHT2PuI9aVT
mQ4WpU9jAWcCwbvrJM6/ZCv826yDxHjnxUJLKixOopOf9QZVXtnpUGrqANyoqQjpIeAhZB1L1jbY
bLEOZmQT/0GWApLzEtd7+PQJ+AMN0AJ8KMhkuV+0p2uAq/NXAOoO0N9kb5M0ayZvKHxgVxzA+Yl+
pZemCBDXlqwwnD4eqGvsKIfwfembRnDVDuo0mkKOyrH6Ya6j5xxptfk8HSt4RF8r/4uITmyaiLpN
vo0LhsHcKrCKMSiq3ahXUdWHdYLDsk9BOzItCqPPkt3JdRo4i8lPvkiZXUcRmuNY/zqEamLYc0bS
TuXq8G5bHQFwlhRA/KSl8vqsDtJ/cDbmFd8RCAT/nrPo3GY8Iz0LXcnuet9p+TSDMSrPZjx9mLtr
uW2Woz/VL6t2KWPv1Zm9zEn46T1ZDxYMou7RguVAubbQ2N9sYuRfc5QbTL+yx2sig876Hfj6Yhs7
Nw/RQ3LTgmnqiuvYjHaF4lJWZ3i+8ada8/zH+8PVbr2MuEw3oJT6Hlq0Ujmf/EsoMnKyNK3kn/zQ
O9ClSxX854NcZUrmfpOS2FQ2Agy69Y9H1z4bI2/qLgzQzNUW/fPdJvwbaCNgWcpR4HyUsk87rtFD
gJDuLeR1lWBENpCzPDX2FMGA9eQ88laXnA0T9YuYTDUJo1/nBAJW8epd+TKTV84g83K5bj9Ikcfd
xRRwrakLeR62zjLUJ6qcstMjnDOxmN+1zvLjRi/fOheGASqm/3PkqQqZIZaEdMOFTvfz3MruFbaV
bk11RbM0bGltQ5qJgQNyX730RymfLOjQKSb4/7rNGMAEYDPuO/r57Pj1tXufp1ytxFAhdYZcz7to
QF9SM4uLaGNOsIroNZ/JLQT13KlD/m8v9AQPqVLlNZasm02AJbfyo6auRwTbDdXZpHme56pYYmhJ
uzteBAXlOqOkvUqrvNfRewiLb8bGJkVULPK5VnyayEPPNrNUKBaScN0iJDnrDp5Cpqn7dQhUXULd
L6zoxVkhbl0LqLDIbDjwHqnzEyJNI6PR3/4ruJEgxGSTCiaqrWiqV8C5uUjdc/tkYjxwao5HuL+U
Xv4J64LXb7h5O2skW5ro2GMvt3R/z602oiQEUSYs3bVso3ndyxu2UbA+gG2sFTKqREaJLoOcVCa7
YP5CizVgQM+5Six9NDp7L1YR8JsXwWE0MhFqOyvIRyMYz8oLRrHk184xrn7YTE0jPCLGMR+x/uwG
8Eq3bB47FC0YnCY0ldzAZ9M2MMiR4EXDz9G7U3I1dZdfnwsPkZOkE702a44f1bkBLASDhk4Q6NVu
p1avm7Etsn5A/X49VLcAc39oQHmcmd/Pa/x9vTgPURkjXLN7Ex5laEHpcW2Rl3RvZPUTTPj3ieFA
9K30+fQ4oD+sdj71tk65N6RGmSMaF7f4I1ki0i+r9dCJ/FKJinGxwh7HoBru2SnbeJvsb9/O8Tlb
GzD2RI/d4mT0t4c7q/nce7fvazzhqvLpP3ZHD/GvDE5YPRT4M/hWlIvesFqxZmXMYPH4zPwswid7
wBhikDSCqqpGJauIroPUdO+F+57BZ7fUc6Rrtl7xktQAu+wcpodxXYSaaSTbRBJR3n/V+trBsp2D
j2ApPF9CDT6Ouy9MXTCfP1dns4lrnERbuXWpjgtbSguJZJg+VNzZAJZDTCMyfkoYWdJWCZ8tAXYu
xqgEA8ys4o0TTvAF7fBqZwFtjEUHIdNFlLzcnjgFoiDwNl9L1Bc4kA+xbk+eujF1/AdA6lCcgtJx
f4a0/kJfqFx3fIWKcFAgMLCp4j1PHQWzxVLibs3LVPRKWYFw9xw4eqiv8+seQt0tsKohReVnObvn
2uQB0HUxxiJwaNXg2In+mC1ivo6/CwczERNLBpyHSWx5oFZQ7OeKyYBDZW8clBFwa2/vKZRluAt1
KDQ63f3CtPkNogEkNsWDgmhWBR4wPqeY4zvBjgrRhDwD5LML2J0900WpWk/j8Pn12chnXGsJcEoN
AuZx8FzCuuXmEtl8cT4xgHAqCgW9M/0t/XN7v9mcVCKa6Pvs6E54WW68Jkvore0R6MCxP80Ggaij
TTRT16iSMPyCWmtJ09tzCV18lGP6qHA5YdiKqArdtlF5+giQDp7jmbIh0Ni4iHf7Jt4XHirk1raR
7cSW123XJz940lXpKy8YQHD8opyX4xtD9E/IXsnydQ5o3BJbSXYUpISdaCwWFZCVAMgyGiE8Vzu/
9IJklnxqoZD6HJhhTX/AOKZi5wpiiM8gnQfIE86/Sbq/jFW2yIokJHJkAx9+M/W/ngyQ/rFKrGN2
W320pbc6njZN+VJy5Rj6MNw0R4HhF8kITGRo/jHDPZO62PwOfnyaL9BWTon1X6z+1s77mUN+WW7K
Ci0tP+71gL3YEfDem3X04LpJJ3iZ6dj6oL6SAUp7K8mEt0yJVJCU2Hp9k3Z9rweJET6sc88H8sSW
qGAEBbde0b7K/O0Pt1Lzx2dpQkbCoylwxnjsgRYFsjZOJm5Xqct2X0oufki0wxNopuXuLiSzblQf
rLUvBS7ChKknl61V/3XcT66pq22s6qQD/ImJji5gNoH2qXVexIHaXiF9Eo+bb6XJ1FX+MApVWk+X
pS4oOg8QuQk0qkCYa/BqDA3nZ5CvzyaE7Id0h/puJYVPmlPB6yq8R2TtD9IheVJ8oPFWryKgGuH8
8L75/eN6gRkEeZEEZUEaRRpS1dynG+YSY0LS+9+49EMuIBcVtxx5SHCG6/cw/ycyWdwuaVGG6Sg3
OA6v3My7HN1csPcxYaLCU1RE+LlBjvLSvSARfGi1M9/q8pv8sWfNKgX//1Ezs4jF86/e8Gz1ngzG
/poloe41Tc2YJ6vx8BuAhkI5dacNaHwF+eTDOj29qnoscw4aOjcBRIYIH49xYGpwcPISj4fZFdry
OyDHpQ==
`protect end_protected
