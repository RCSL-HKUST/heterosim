`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g0ZnWWd9McEFR0MsfDyCsHV6h8dsTUqlg5GJ+EW9S6NNsEYSYyc+PKwihNdzjF5CKJdAIpWZhDV6dij4N1T+RQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a+ccDKedn+93oXv66fLeUR5iNv/RUrVhV9c6a2eWCJthPW1pG2Sz85QOvsQ0weiO92yQl3Dqmsr54e59nj5zymSrA9crV3/I1LKjxgSJxKoD4tW/yoifl9BVUaKULvwPzzpil2T0GPQsky5UTJuiNmD6ZY33hP8BVoSmP4qIBvM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tp3sW7PsqEWhsY7fkA2/j2lqeR/zUdzhWaHAC8wObv0XQCdgcrxXmbdDmYNbcCF2DmzzNuSwXpdpNj05Puqg5AsJ6k3ouIhoQRYqyxkdj6oLGakfN+JGVPFIa7VuUqqFNKkXrMarOtDLbi9O+OWzk9QhSMmq8/XSzTNsossQoLZ5GPHC1LZQvXlxkWyE7APMJIqpzyFnJCGmTh8quCpljYtO/QmQl1tqKygRwjexDVOt7WfB3RASu/uHRLTHzpLylFrlPSWZJ9QyQRq+/WgK73xcCfnmShGwO5zyDL4/d4ofUbdvVSHat2ogAHGlCyIRColJ8Xy9vJpFpumJvGlJIA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lwHa5a5gvCLAY2870y03M2ltq+SZl8LOtLO/XUNuHk8Vs9bkHYDFUp98hOKexwDHekREsWlJcb2UbFr+CZrGUqGhXq4xoWqSq8CKOJob46IL2fIyNHOvbo+N0k5E8Mt/RnYImkJ57MWvL3s1YegHIJM5lwxBUuGQ/M3sxVim3UQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KYgGVB+Rqk1gfG2IUGlv4TBZPYusKVbvBOqL5zDqDlTBvpvXyCwwV6yn4+wTwElwMhlgTsAKU39bOVY+ep0Kcwo8u+7FJ06d4dpiVjLdIqhPXAtaSXLvWtiuleffa+LA+nTly/4l/1e5Il0mhSbmpm5hNYAI/aQ4XXHk8Bq5yUriTTdfCXiDCMX5GtOnbnGZ5YpI9+ZlVxcQBg4pbqM0VZap6dYKMpit4YFQj/66YfB6fDE4Aq5Mb2uJc+nmlGKUeYGmY+yDAG3Gw1LhAc7LNkXWtL/TkyB9+jUaKqK4qYBq7OFvV9uTbxCc6fVAt4h/M/btDCRH3kfI9WciD8d3Og==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62810)
`protect data_block
D/tF4VzP2UlQUV9CICMOWQDYWTDSplnWmxwP7sOqj76IvisrT2XjlRSNopnHvDaOOKd8oyT2jrhK
eFa63Xpv5xiL1Y5SCKZnUKKa8Cq7GM+8Cq6LpbMyVC0FGAtqCc767FCz+Gy1AxeUnhqXi0+fs7mu
be5PPWt3fvxmaIE6W2PA3CPt3nD8TFnBXGn4Bmiw2HW95eINx4Az57kwTV55P3ip+gTjcWjo+eMC
PH7SS7lkKquX+BB6DYtl7H6vPDt7xbd1RkYDLcDqSdf3R9orkUBZY0H+HMpDhoMncUfQgw2wz7JC
YkjsGTZ6/oG+YJciGtuPWMWrYGnPKWbZFKvKXcaKcE5mKyQn5Uph1tzae6Qylw5gbv4Rgub6Gs9d
Xuk9ZmKlkgKPZ4eRbWTD8/9Btb767JpAwwY4nq+ow6XnGqCmdIXFwktDINe1Qgk8qH7o9QHTkjmU
2rbD4dBSQQQm5hePrfOTV0wzF3H4wHM32TleHz/Ju0cQ6WzUAQ2g8rEBjRfiHTpETiZvYDAe3VWB
4sdRWvZKrchjD2vJ8NbWkgS2tqesUYcdLcICTsYoRuK5xJGvoG9mVMW0pSwuevOt7zObm97ovuK+
7R+R6PxSphRiAT8vSCnHdNkOY3NZkMNCpCQip7k5hwFDcvgeeDL9TMMocGAUPPuzia0RMqbvzn/l
gwTDDdxUTNmmzcA3I6z3rWu7tBYtPlPGQjNVokwy5zhgB7Xh62L/7i/ZvTFaOsbfXEb6oXQSIwxA
VusI/bx/8OvDOb8k/PS7RedEz/fK+4sXn+GM3JRZytPySYY2fGM7j8AwKbUaaq+urjnsBP2YCeDH
SxHMUBAOn19Pb0XK8xp0L1TyxqoaXnG2esP0N6jHhq4glTzK7bwwLC7SOA9JNhAcbG/+F499KeeH
84BcfjH1BPxaM+2gWw7A1Hn3XWU8qHAivU13RdU5aLNWfwloCPqbj0KF2ju4rUsc9NX5QRDSv6Yh
US1vX+EzftIDDGbEQDrUewMQZI277niwg2/7hTP7FjZpD47vMKbdVFjqNAVrIS4ba1gpTu1TJ4tp
X8VQUJnY7kAlA7/2ZR1hsXR1oeFFR5z1kzbKCw5p6PqAq/Gu7fRQzdE/lSM8oesaBLqeqIl5Zwfs
yNRZK5pPTGF8g1RFO3nG4qMmhnpArV6S9jyQAj6kKiAs/NIVfQFAh4PSyRmWZtRktJrTVnnnAXni
/TxGOexuHV99CluI1siS8bdzVvpNSKykSJvi7gGz7YlwI9ovfvRYUvH7h5b6uBpzXQ84CUJt6Deo
6gFAyjV1cakaJPXMUjo9Y/MShdxstcqgc8YHzCdPjkFzdihuN6YTvXdZOF+RrdF/lzHjq0cAAfsy
IUNpPpsoh3arVAFIsYYeuOE6zOQuDgyx+BVnJOSLPyJ18Hok1B02ULQacyucw89fZR217rXVtn6E
3Se0j09KqP7TaQnSgD9V29pRDZnA1Lc4XAB3ue+sYAWOX/sZBmCe5aMyLb9RHYVQCoyTweKuSGt8
QU08Ap+UzYO/G8jDJ6BlzB8kWZSfAGz7gcHlEDNfwdV29is3uQnk2UjQEzySwrsVnHpjYfEYZOs9
Yh803+GgxKwrYjLjEi1kdzqs0EHQeW/qQGrFeTNTmwAW3wjMHnCwEho2Geft+v2SdIqIh3AMla4E
73kg0VRKVSg6FHm11rqY9QxJQg2q+5l9pyWJqaHberpXAKc9MQF6FG7rl+udGko0qPg9rcctSAJN
fwkvNFFwTQY8JGNoKLSc0aVoRxK+4fRrbQid+xX1FIvCECC+aNwjzbe5fr0OmuFHoGhlQnH0qMDG
X39oUvy0J9IWfhssvls3Yem20xZDqVRphx7zDHzKvfWCkO30yygW/iLEgwk2NppzCCPbVc43hfth
9vilhE4Rc4yeC7s1x0DYauHwmMhnjHsRyebhJpOqMtzQDgViCPQDinhkZuY1lSzXpCvOwXUDgply
YX9OCZIfUZw0rBGOc0uFbptGdYtoHl6U5cbJalIPJfBnQAcsai8fSc+jKd53X6uyxvys9orhHMzS
8Z4lAJ7WaILp83XcSM+my1+M9IgLLHA9eGFnQnuW8EWhIxjpG6GiUnZcxmbWZIEPs3crRnOcVDwp
J38LDQFDvuFMXqIfaRtkI+gwS2vXoMfS9nyEsqanPaJC8wFY0Erq6/y256nNyRsyAVtvojiJq0LF
7ijzUY7iqj6PqtOog2qnBIgO2Dmqh2yM0HXk41+TdZcJNqPfUsnp9nW5OVqRSlFe9nHvzo9wEeXn
/r/5stfrehV+bWknucr2TTgmHqphymr+rizUmGUn2fg3wLpvfsRlAiI3TazsJjcTEHIyLmaFbu7k
a1QqeKE8Fu32TYo+j/b0GjMaZZS8mPTAIlOAU4YxPWIeX6mOeqlkiddkGZWW59aIqffNNwuEzBfu
5mTrIXLDUXJI6da4rupojs+zvSz6RshuNFWeWt9Krj3MSMC+YMwQeb9nVOk7zzg+xgQwKLv9imde
/YsrtE2s6nU1g1fJisQGSY759PCj26C2gZQcAuE1IJ5HEncF6rNYfNi5kqvT30QhJgWt2DJ4Dq1I
8IKOMzbbgvksptzbaFL2yEJAhB2fuTc3tIklID5s3uAOLSlLTWXNJog0dAGt3X04CN7whm8LlWNJ
YbRySjjI2gI4cCJiC2qmzV4TCzj2uYtw196cONBC6JAyzhW/1yZ0ZSak0nYpFQyFGtPtmsScjNW/
3bszIRfc5lA0axd28USYFPfMHZ8uMDL+wtccvrlUFda7b51QoDyH+v6IcICsF/bu4qBmmp2KW/IN
6nquPuC2QJtnMJMktNVpqG9uAVya44+/r1PQB0UkFsLpazKiokdpWTYPNwxoa5v6jhOHV/G1YT7k
MYN9MLb8/OtY0wEvZ4kQqlMYSRIy3wCa1MUwK+Jnyi/FsfFRGwCZDowP2ZbA3SbZx6YAov4G/yyG
Wx6ZQK8buV5XhXMP+m0dDz96yEU83vvSRiEuSgJo5of7E5BVthk840CaDQexcIDCSglsuZjHY/xN
1e4uSqO0z2bxjrbaDOnGgzhGYokipeppBcObIUTgLkRCqtQ8mxHWs0a0yW/Mt8cLDrqKGMbvReVF
EADEG0VC+y7z2LpQ5n57+wSUFyCfQC9YIdyI43VAUnsxl33TY6eAS7IoEEyDeAXp4ZRfDy0tOm09
dioErxNWcHO4apH22QvwSswPLIfPVhHd7tkvayKdA3qXoLdUS5mdC6WfMaLgoJhq8C4u7mbxh0jm
dD4oyDV8E9lBFD6tAsGnv1dzmVvMIaFy2ZR+/6+ygCg2MgvddggJhYGqxkmeorVAw1FL+wvcZRLq
+ZUOmRt1dGUV06tTAdaua1hrDFuENu+VDK8bQfZu7ljDKf9OADlkf8lrFsro+AuHTZSsOVKiXU/v
Ae1d5dKeZrHq6EugJoTYeGyX3Zk9ryjn8gagFvwU3dkt493o/TIthIupgsP/Ovz+k3zRTTSnPKem
ELwLZnj3fZpuutuwTtHtMVt5s0hhxqpEJLd30loMFt7j3GF7xz78KGmbGxqRpk06dhyryuhQCdIG
fPnVb2zUE43PsKrXIIRugURdoNbOhLU+Qbhw7WVmkON1Clk9j1OUNvarofOc+y/yLT4rwT5TkPLb
t+fMen5E9OF3WmlZPayxHBau6FwGy2CWHwnTwyRPj1u/Euvpcqcnaey8AEaa/PphWuX6FYdJKqMd
bEj8aWp49bm1yUyD4vXgWgxUzl56PkKPC7lmeDZoYRJX7sWd7uG5YZWojT4+RMsXj6TbinEERXX0
6jW8VHO6dj80s3LmaRmIx+6tPW+Y7T0Bv5ytgSmmYfgYhvLQGmKdoJMXlwWjSXb058Bb2FT32yZW
CnHBShmIZcM4y//XLDR0CsS7vZ8QA+cn2EJz2ejzGRDlJg/7VXG/2Wznb/zDR0GT8LWdmpJJrtWo
Jr440hQ9pNTxktiolHTlfTIklqo3HNc05eSaYUnFrJk8z4VTdRLBCUL3NtkYm32JCV1mffQOb3GW
rme4obCScOJqSf+Yh2WPW1s31UXBksvs2wfpdVguLG+xv0fGtewXQ+mGifQwGCELWhARf8eY27AJ
wxtZCHzrA/rtAdjWTDYkaTrsl8cwauvHTUK7KPs8HMzCswoeA+ILKItT0vNlyP54yvMpjbJCi1fz
Z/ngUQL0QCjGZHKp1YmSZJ95I6bbcHN/4nyj58GZHqByezl+qD0oNXYRMwNCkmOyGE1KnWU3aqpd
USfn2sbNxu5TWdodOlqA8inGspUl/f1wirh3FFVMWgT0LFVtkpShgmMy795FgDqf93AUGwczzqH2
4+yeiQ5lusQYnPySWf8G9qDijWuQplQIQiE23YLYihv/TtUycfjvAg67HxWWfme5lhwa8zFzSKNt
OyeKcxbJl3FYMYqUppk20iEGzTfr9qAsO+VQMuxWQFpR0WvouYpIsdxtDMA9wk02hhEyxnFCNuyk
UaWZ/EOcvs8viuOgfu7Em7QCuhkCjxQwkW+ztWjY7ssaqDIwv2UDOG6yKtQ9kwJVf3DCVUxG5kPk
KMXfiH82EiLCA/sWBPa0Evn7yVm4kTWa2gZm3miBHo/CCkL02T82Uya/O6nyxVQ5c1jjdJ/OlvSS
MhaiidE/hN9maThdfmelQYUxyhhZsggV8gO0yfIENhy7zT+omtMgpniGO45xqtqGg7Xfu1NDfHPo
VQAcUEgZkH5CfDBKCWANIoOnTyC5WPs5Y92SRIk25ZUGco00zo4T2w4fIlBL5lvt2Fx9vn7PQ9NY
r9NozfV11cNPXkAQwyHDu9OzIoEhO520O1vJxD8LlXObvnLN/AvmvIUOOrNG8tAIZ5xUGuorm6wr
M7lJE8peoBSKni6cTYAFE8UrHh9TuZrn6rA0OF6pAsHPP+10T38RnH6C0ROLGBxs/kUkgmCFvyFp
XPtfwZwUntTXxnXjR1+zXvE9NjRxratqmlw+p8Xv5a7uL08M5pA1IyEx0R7aOR7ZpVGut2ByR6Jc
BgI5ZHxCxQwiGZi8F1mjaotHDCn22T++lwQLFyuB9jjvFlvfaupAl+EABzP9cmvbmTR0Pn3TGAjR
lFMT3H9v0Iei7/NwMMklc9fQaxOwcFnn0cUOsgGCJ+TQCx6HQiZLSOoUfFg/G3RLmrLMWMG7gcV1
hn1X6zOVLHbPdYzvDq8tQV7cCE/LLws0L4pgFAZiGzhSRfKhPFp+uQXLHXJdWU1TW9h44WP6UXlP
YHJAGKgxw2/KbDuqtEwe3iPRauAURDqWicP84RJkb30ECksVIqkR172nfI1lGx5Q/OROzEKypowI
8xP9bypACc23QePCyNdHGQAhM5UsMdcSo3++kOZb+GQPVPg/4Y0o4K/ozWbw2o4bYkiWIRq7uoVY
uJFCgwXsanymaTHvcr9pG3cjtnnR8l9d/0xIu6Oz+9CdMy6KoBqJo90NSbV/sVXu0sfgyV9H5JXN
xrSDjJXSLOJ5qDpfT/+y5HE+Tcfl+GUMKAtD4ftF2ySQm/2MbewA1uNFXr8uVDjaBAAG/dTdZZxO
pAUA5Fu/1DjXszzV7x33t6cm/ongC3pA/FOAZCUirvZjISfI2inMaC0bEUiYvT1l/pkc6L44+k1a
dKl4ieBnzq+f9CU5fl+ELI1eOazf2GBMezyQYgI9HnY46rSwaeu8HXwjxlRo83vNaZLSL/bKPZ7y
yH+YLZ5FFYrrtCPSdMRE7SX3p+YD8jegpEtwcgQVnn5SvCmwZv45+v7xI6Jok7hi2+EzpRurbIpm
Jqelhe0K9uH9z7GhjNoIlVoB0xKjlq6PfCIQ2zxNXfG5EOASAW+iP1zyDEliTWZPIqGqcC7bbep1
3uO/Xn912SYwO8hUdVlQBxaVr7mQRekOZPx8plBgZTqYSQ28PeaqEbEZk1aL81clhfPfa1gXR/RK
gKNvJLOU2syScZ+4zw96tSwS3p2xFI4FmtYiZNvu8I2ydpM5JBmo+z1x97uGaKtp4DOzM0ryg4nX
t8jjn+sfvyi4Y++is+ZwYKiHM00b+/iUwYYInRS0+wcISJnWisBxgf+HDFB1iC2wkaDl3jugdllb
VBzTzJNpN1/aZmEAB6lHLetjc9HiAb+mxGAZpRc7G5qiOkd+PS6qpyVK378y8IJztiBOn4BsuOWE
K8359HLlSQiAhac7UzHP+0seIvAI193/GxOVi1nqveNWfSsdue+4TqnRMbEtUk6h7ttUYk4fvTFh
aN4zEL0QR9UhjZ4dTNyXJCnnt2KQUkbD4X3xe+Kr1Cu6u7JTUa7aC0YA0FeNV1oLu6c3tB05mOTb
9pGawm6MiA2tlWroPHBXGQ8ZCpcaT+H9X7Cx2VWe3Qwi12XVhbzBzctUZMp8iPRvioVAkFrCEnga
kpAQ78R9dDlLlTrW9Q9PGEVb1DykZsfrOhQWCRaH030pojzlRZvXcWXvCcYHXCVjUWo88Vd0EsKR
4RWL/ODPZUeSgOEcOepuekqz9QLBSUXtLOzW3gnOVcjzJySoXOHw7XvHNiyN34jRJTBoq6Qa3dSw
1jtVt8MqkU7cAHUKxJb4KkKI8hkDnE6ebJUAqyaPv5PzQ4aAHWhYWxeI0EIogOwuJc6VUcwSEe/K
FfmnpDRKL3XMpzbz+r9tihthQVRk97CKetABhPi0VKKmy1h9WAV/dbhBmlG9sHyWEzHbLvUMEefT
tgqyh4vlhtMpaOIlnI1Lhkejqq7alb2JW2zaCTMi281WczmflX3UN+JeL3HNe5cmhqfHuBIXIZs4
eTvFpBKj4xhot6lIzpDVbgjNnns8e4LmS6y6UaXTrPj8YO9ooAigFNAjLn74fjGylMkxLQK4HkqD
8yM6vAEuX4xqKAtv7Jek7gbAl8gbNBpqquxpe1HhNX/ZFaB6EAXjkV3Na6RkB3Acs8R0mrfW3pDi
p1BZQDqsDXmjQzyHv4ybiUnav9omEEJz0/i0Gs2G6bT7z1C9Xg7/KXORVIYML29td1VKvfRwarqu
RXK/kcdSeWV5B3I/VOSCuJgca0rHNpCUygVQrKAfCW328wNkQjiSaLATo+El7DNa41dmICXq6Npl
vkcH4yYFaF2IDR5iIlnlbrwGgM8UB1f8gGODv3iVwnQMh/9bMdTLBD6Dt3oszz36SLP9462N77sN
ghffQ+ottZOT/89F8KAGTYcz9fe7vB0RsZOnTd0wnzTcaFksraKf6YKesYIQioVRF7KMyoXYJqTx
GW0V6AzjzAkSiEKl6//Vj3ALr09AQqJ+63odMG1JakccU8zjA8RTCo4HLuriU4wE2Yk+2o67C8DE
sT09RpwP6U7DwMf+27xu5Yp3CJlGfHn6gEIpwPH8tMjHtjsbk030ysHM96dIXC2d15tFNwpoUOjY
yuVsbkismNUNurXIi6PERg05h5d+sCRBo2FsMOmabYNN+e1xuBBpSCWFkal69Ugm3BFre3Wq16Do
bYTVE3ScP2IugIOeZmfYHB6U8x+T1lxMoM58l8FDLu+vekb3uXHDTMdRkfu7q1GTUKSKLFWrbCLU
Txl9rmRua5TcD3zn10ClDqMeaHQ/wzN0sW42MJB9BYxoJ+CVpRzzLcOQAJ9UWxKyD5hRRfKqzSwz
y8U2aVyYCGzr+rHoJT/0/pKK7Bx+BSFDONjYCAgjfzjeRe/QHDxmrcPsKpqccs8nmpk2N9xNzI9y
8IQU3nHqInmtdDHWuoIyUyWIUvvEKlQ3Daq838mkAnZUG5PFkkou5vfuyxTakpF6aCZwOuCgBGWN
YrhqG+zCjt+TeuxsFUHPSqMSgKwnrwv5YAEhh7+VwDx4OU5rt6oPRHu5Tr30gpHYJDdTd+4ZmePa
B7arqGp57kuucVhmmZvu4YN3GV0JDzwa9lIUlJPo9Wu4S1HLhYnkUjEhhMoXVdCuB5IvBzzu1X9W
fG7zTGJdOQxgnKgoHErbmKNfJKPUmNn9BRvj6WehXwHWUytgcaYZFoUhEc0ZuBiBKHZQZDvLKvT0
HGrO1YYvZdMX0vkcekwN4mkXqik6RH+nJ74ZbYG5/tRk/gchmXKJEbpie0pxn7Gu1KY4obValKuc
5KTrrzyWnSVkzT+SEFvM2xwLjTem2SxhPcsC/sKNiKXj8Npkqig/knneVnexdOx6cwPg8o0R5tnJ
oldtVLwgKAazuz+/KEU59vYp66bTYROeYyRRJ3AxaZchXkZmtszlQSzUI+gYoOUsR+b0xgpQbDQk
+Wnf9zM7X/YuNR2schg2rxJGretE6T7/50PvbLXrmHxPtFPPuY4+sYNcNwG2EkvnupbjEpf72lvo
mJxBfOPvbrH76xlTPKsmXPqwqX8nGVshb7B05yIsw09Zk22r/7tbMb6/MepPSKIM+3p2eZgUQA7E
dXEeRP1XCUakk3wgU/mDgTkiZqGpitra0g2DJgwjI3EiwETzdxTB6edkJVgRnn0zQsi8hc1F/JUa
XbNeaPvBX811GOF2rza6IwmF39c8SSp5bHYll0v8+kG9xzAHQv0+TdRl5lN/GnjUYm6XUcONCcDA
BBRDkxJnE0eb68m4zKvugCAVf+e4kzqFoYO7tW/S+CrJ6YnFL3Si4XPkHeHIQT4nUaZm0/yVTIGh
Fc4yijGk9y0dYewiZDu3SYgamTYT2ya564ce/XGi3UMXs0C3kTZPIqwB2TP/Y1jC+2VvFgWkqAbe
df8EPrFMv6Lk3+ea3PRwZBF/vqcPT8Fmd79kyGqH/mqHWEgESdHZ92ylu43rF5ttVW+HNg+Ca7jh
GqQDXMn7YdkLEB+zjJQl2efNQysUJmot1vHBQ59NB+vGPCej6HxeSN/h0rOjWYLT3u9/EEs+1KRR
qKCFWCiKHdiPzMme4bVpKb6I3LmDfyT974AYxFa0KkC85zBW/kawZ0QFCWZ3wXZvOOfH3goX6/N2
TkaO6dmJ2h4D+1CrAw2Yikztg9NNP1c8H/UvqTP327+zOefT1+SVqPfKn2LqwcC7QYSzQ0mcsx9H
zIebHjQo7c6iTVdbPawFO8DobIhFQ5/DUGDT7AW33+XGzApYQS0eDhzu4Dq8NKUMSA5XN7V9BgPy
vabIx2BIB8Qq0WXav52U5NvHnz3XbODVaGW6jeHweOrMQQoIyV9f+E18j62YDYZQ6tdNHq+IphNe
DsFL/8qHpg7pVeTsCycDVB61oGxHcPmNISkCw+Q+H3fKLBwR52gY42bXbvZ/th490Gu0prJvycG5
Cn7te1HDBBtMk9F15gKJmy7RtQiCvupQVI3ZfH54xqfCObQyYC+zcyMq5NkUQ/Vf2owhAU/bihJB
RLuQ3yAfAyd6UxBtAFznggRel1oauXml3P3OXPDNGN2H5qXIhYQBXiAbCLU6Lr3ebnDDSeEnDrKf
xuZG7csL7gtT1Tz1sJIlexT+bQcB37jEapWnYQdj91YC9f/KSkJ9rqUMoxpZXNTbw9KgwPPSM8Ns
xffqpxJoH1jxRHqgjaqMSwjAii9UjCQiW3MkUhS6cStMxeoqCaeTNl+qeZzpq1lMgJjHZQwDsWgt
QXtQ0R74eh7LQ9ix2oskX8rXNjWjNqQykpKmiyHl96hKs20Ff3tLbmV4x748Cx/6EytmXSEZejxi
CFnxyL/fyXcD/08BWvZVsfD5f43TuznOd1XFaEWJ6WXYBUNL3ea16yUewg+aZHpTngFhlOi7MDJe
clJSZZSR5Y8c9LSB2A1b/wA0WaVo8gwPQwiz6AmRrf/w7Kzu6TqV45RixRWLFOw+4vcWRPv9jDTK
zTJhCYqbCm4NKp3Q0wY2CNzL0EeSG8p1ESa5R2qm06p5s8nJ/4r1OI15+fbqv02iOR2QHQJPyMB+
sSoNxDJhivUBH3QoKYlmF/QtKCHhfx/5gZYSnns0xEu+cOUybZ2TgWq2dkmr7VnkDJvlYnv1N6ps
MiTMIBKGVh/3L/M3cOv7/LLcGcFBQvn1dduTIe7rveVRBvqtiTHmq+QwH1wJJWgRqYTboD+DN7KQ
8sOFtG3tXSwn6XqY2bOzIjjaLLFqb/8uZcQZGbeIRtw91gdFH0Z+olh92No94OG4NLzt90M+At7H
YM3c7NgFNkBlOnQkCjLjmipqaiUQK+hxjlpEWl0dK/whyttRDIXGJrS9K5MZnMJNHfmez6YeW/0K
GKnoqRqyUhvF9qkHYplMhyySpsrqqOn1B/vTlA991yOhriJyD8lJiJI0yddNkqvrFoAMuWXPHjVH
74MrXTGQdUnvX6xni4ejWXsvD2sJ86lZjGvsEZGwYYhlPzo34csFrqeRFCptfQjoVU/jplNgU55o
9HrE2T1l4n/HEmoxtbqPRNjF9FM/0iMsXPv/D+3dSvU5R4zx++kpmv62xXiVSdyE8F+VgL7kkmEw
f0m8DwCNdqEL08YtQXvB1bpUem7pyNEVHDZ0PNoNQvK1RdqLWNrvAFRsz3W1+Tn1pdTUPSzUZ5WU
R7yJ+Q0pAlrK6eBlEF8CJE2jQzyJ0DtcrMouvxOcEePNRbfBOPk5EirbppAgkUMqGUhCHv4t1/NU
TFqoioGDdZfXmkVEi5SkBSbDYjnsoLP63JDoEjyQXMbd1eTQXCLYblv3m28IGa20GgRaOQMR6uMW
M3XY2THLm8leKnrtxZlojjDab+49rLVwgfSY/8RepcfilfvmrF+y5BzL+PyJiZQsYNDfu5z9PYQj
U9nyh1NGeUK26nG8uW2BIdpVR7Yw5mxn+Ai1+2/HpnZnioXZUefFdmR041eeo2Ws+Vv9/m7nneH6
vj3NBCT7zzEMGjGJohkhWdO9cdpPBVgiN3mAO70cNS1TuMm8wUI0LOzNvCD6ixk6smHL6TIo+Neb
1/yGJiqCs4AF073KyWefw3nh4uW1jKKfdaqmuaZkBUD7RRq3lYyz9EGTgxigRM4yIuCSCnRViNFP
YBmXZI+DwlldW25ZOun6W2IYbBeXCiAkg2vI2IP1t46gWSvLQ+gFbaZnuiYznv4JKTyt/HhIy5jr
IzwIPQ1hVc+immXDSUVs8K9+wdy3TXqPqkWV5+fJFL3Mdm3fbflbtVmiSy1kxj08kJ9B6QcbzRWc
Inon+rE2NBT7KYCfRyS+PXs6FfCEjJ60zMPdcTuDSq4zomODiBEIXEHKClQUn56WbFJCh6K782hO
TgDWWDUR+C0TcAEPiQg0eSxlQI47Yhlok4g4wWbgOSNIjYnfoN1UQkj2KuyPv6BEgrS4Z93gbD+S
oGw8veSeqHNkvTwE8iYTw9Hl5l2mEFchnx0uhTdOz0B0tSJW121GsixC5g8GS2BTC8+P2FjAhB6O
o9OdoOQAm2OrFxPI5euQPEkNSVYaC5XvnpIcg9BaWngCv3xeCxlszrzPl+ATJr/EpiE5Dy9bt0hN
TycpPYRcqVkoq2LQvLl0T8p3XGstz/GnscoTQR31hF4nUjAUE6rHFyjwms5I8TzkUENr9co1mApP
VyhnKIHG9Vys78P1SdCj/PKXIASvWgLId5mMQAEcHszYdtFY6p8jDTDmUugYYcIbzY0PugweIf/K
V6QTzc7pZdvPYnqXN6qTNzQzF2cYqTbrVMxP3Q43PUoirjGn6+gChbE+IDdt7/aDwS7idhUsdM5E
/8F8PHMRcXk2ssLl5pSmTBv66XOo/R4VGR9SsuqN6bj47mqHi7DF/eTtpH8iTz0IIw9Q6QHSjNZL
gcy1+RHco6q0cNIfFPln6Z+Y4HbXuDpJqDFLZr07QMqMN9Eb5qpTVZps5ho3Fsu02nvchmJRGjom
LykMJB8ZVDzUI53+/ogO+VXqIYtiPZ2MBK/Tz/++CT34+i7djz9YTn7epwFn5c3smljQ94dC5SM2
oOv7tCw1I6FkjMSbYsQuObxsrrMsajago77xzWivvgSvsxbPjeLk4xofi/kYR7333eqrL8O7yG8t
cAYXCMazLC7wgvOwQ+Ru0ccghgPkaoC1hT44Te65ikR21BZK4LCKv/cC6uH7UzVa7ChaqB+xRvGN
ce/h84tNuEPmps6mspkaIOjEFdXdxtu/4aXW1qCGpMzLbnzYcGkJDofQgoer2vF+wkE4hzHyPzei
vy5Lk1GVgvsZ6yc2MKoUcs3EM8xVgziPHG6YUJ9UdqdKOFp1+z6C42o0NG+WNtvxJJd236cz9Hzh
GDSSQu6ffg7YdpGuAxisehnAlBOYcyUtmCOOV08PFfl2vLjevyRTsCvrEORcVwjKz9EuT/bMNScm
ITcqlnIUZLqsqttd2ZfW3BHdbaGgo/uabo/qodF+CyMhr04OuzwVL41+ICTkxX4Yx+7oAIPDn9fU
tB7jVejGgZmykve/kTACM7pZLI0E3nX3Oe/R0prxiYU14IAplysbq1wIn2kRne2MxdfUXzCPcezV
zq2qiHBOnFLF3DHQOQx1b3WkQtD4bEBO/0iK3mA2LvFdS/d+OrvYlRe4+j/ZTHHylsfRCs0FD3Ku
2qgqmIlkw9T8p2MFlV9ptqIM2HNZQFIUqpypMYB921ycf4U2wIDvSvbAsctWrjH0erk0Day2EXcJ
GIWevKHOG9vg7VPTMOt6DcLLs0Z+TTHfcp75UROor6kY4R9iwguBfsENxLiG0NfqVj0klEUs6ttQ
yTRygoIcEluGNTvaKxH3ocYpfZLrXOhNeDeD9o3at+bStuKGQ5qK0LqiDvSaBfA8JRNoezpSjA90
Qhdj+N913k76mbG2y0V06O0RfAnJH7K0ZJiKXs9rqc+DwBxRn6y39SX+dWfzZGUP2wevgs9PchnO
dWvrWfCa6uZIwNdFKAPVH7UsqCiQneWKO2PuEYtgYm5OdNcuJapjzHLjqXlY87QSbYOWrBRm5qKI
pmLVhs/Ndy8tmG8lNt2tiC3vt6mGGJRzhOUFVpaFcVU+REq9JCOlpl5uIoe765q0dZ4HSburC0EV
cigBhlTAfVLCCfirvTaWIOka3CXuEWf5JYXpvNhMxuVR7RB1jP0tMMtA1P6NJI7yala06oCO7fB9
RtFx/s8gsOBugogAbi4byndPaRf8uuQNJwdJrGIImBfntUniR5Iz2Cl3zATdMs9Ube49Z8o5FSXy
eg0gAqQM4fMNcb3+8D976KNYQLZE71QkIme8Lqqdz+yuNQzWQxSXQwncBB0DM7+Pcsd/S3iE6dEk
o5rQjppgCjJnRodhFb3AdHrcNMfynOuiq2WlFIFHp2tpO6rYRMNYifIBD42zTCysQ9AwMz1najgq
KKhCTbK2BC7VTqVq+QDOGFqGLw11C41TwdF1wsEe8GNuEjSC8MVyy5B+XZX7qRUKIyhnZD6UiVuR
3FL8W//t7es9w59BIFJmI6NhFxfB6nI7P0sKsyc1LONTgiZp57eWDxzfOkTfroSuQ+9EbFLCcE6U
nJJ1rHIa0hi2OmQYf8htEpXeL2m9mROL35/5DS2TSFMua+0fGBH6CCKppWQ/FzC4/B3F41tX1ywc
ABg0HLalzWM2az9rtP0fBaS9Ap4rCetNc5en/mFXObdK9ogqd4I77dfapPXyaCnTOwaWEI/M+jY2
BIKv84DtR5QNGVYExM5MDx287jaKZQuQ8RWuLvsyx1fZPl2hcB0CM7OnRouIZNoboaKlvhxvXqvS
lbbisPmEZpPJD3wGnBs6PefmnfJxiIBPc/0LXbkDyvw1tU3ZkpbHz8/armZYIYXgZDDxSlH+yikm
+tEYp9znR+GlfasFPrc3EXU34HZ7Q18FAXIjkir2DSIm7hsCxDAbkuf3k4AdxlYJwiGHc7c5AEbM
hriFBt/8h8LeIzmIsNeRtQs1woT62XMeqUUeIuAHciPJkylAK2skijALXAk/VIwejjxVmVwEClvt
JG/9+u0+ETQh9jz2w2NZv1XIJ8w16F1j6osI2Hf+90soQD0w+TZjPVrh3q6IeZghzX9f4AlSl39s
/lWIRYLdS27/+8pH83Ol/7eXZgc/i85yN1wck/ZseWAfKlz+p2CuAqGpqeIXJkFMrEH54dyeMshU
DOxHrgUCqKAyfcaihR466IUjk1Wf+6Zmr6CI4fDB/0gPhfFBxs3qtZujXTAo5iwKhT/BK/zpTIFP
hyqoBL+wLc0Ker3vYhUl/l2Z5c8NIzp9TcKJREKuLyQRGQSiDETugncdilM7mDpeUeQT8v3u3M5s
VBR5WFeZ/IW9YD2cY9xI76XkppuTrjdQpz04/mAZqhdIXDo+WEA8nkhVQnQMGkAEtfH8IB5rzFQb
VUjIEhpuz8v8oIOCJUA/aRVA+50YjyUYaYDOPN5rpOCr6bCz8vkdATglOhw7Yn7tVfWY3JRIgM5k
LR6UEesur1HuIL4AdpA86dWmwUDaoFg/bvA4St7BX0jNPORnUjetTblPbDIYaypDoBTbc4cyfRP9
cZp44Pm/luV8/iUkySUvDj4g6EyRfpAxbgZJEUABoKj5ObOXwkCX2uOxzm46liipPFqUNuTXG4Wn
WBnePBRl+wc/+wjO7U7CwgWJ0Jb6EXIeRoP2PVOjoEiKxt3jI4zAR+sLuGu3dZnhaHOY5pmJsJiP
qs5/XfhGUwQOn9XRGYXwHhgE+9EECvXmbp+/xDNEP1Oys28kOmiN2dLtqpe2yL492CYVnhoTdi4d
YHNs3PdlRaenfgZWIDjSH+bKsF1nJOV+L7kyuactHikL9WmUcgB8TTyWCRvsgz+hWciZCGnYJq3z
X+n/1HzLrNYYGx2KDmHP4xAjybyo6b/G3PouED5OWqUpnVUFz9owFZEOvPY3qTlVpSiNhm749fH8
yBXEowzP6WjbOG8HBIQK+tm0NTTJ89qwaEvzXd6B0h7u94m+9Km17+KrEdfnPSYgmpppPL0/4HKW
MBx9AynRN9GGHbVE1uDyZamdqzC34veexW9F3WXeZy//8N2hYS0kQkIp0XTEyjANMtQjMjN7pV0m
qLqveNy+R+pJlHEb6SyIzXK9iiXZIkHahPk3GNngARjdTMyqOzTIYyiFPr2trWrz13fi/xCXhRLb
+tkARy0bgi5NkRx3+tE/sKMj7ms9AxoTPX9Ylc66W3dk7oSX2WRUx66wvkVx1IWV8B/G9Uyi8sXo
j9CQaK8t4lYHovNXHjOzWjL92iRsfs95kPwj6sIbPSX094tTCBwl0W+48I2jHb7OKoOTToaVGcgW
aykPlx+l46yFt6qXEEwCjLuB/T3GpJuecbQGEGOTn9XYcP0LtwrFLRdoecOJ8ptX9lf94nvCSUHL
1UTW0q1XhRmyaukz8xX9CfDkcdUQy3XVxDiYdXPWRN24cg5CXLc8WSCFGrigvyEPl7DNZGJZnJdJ
/u3A3d1m0ZhRGZ884u+BTR7hLj9l59fWF1HZrG+aBWyL5r5J0OOQuHctPbuS6TwYhod0KfV+55fX
L7Bt5E8Gt3+XflPoz42FipBp2lW/RHkCiEzKyZ0rztDZ2YNVfjWToKtf4Sv1zD4q4i9104Lpht03
1OuSeyp2CFLnc9/zO0pYboEXb7Og0suaMRq+fRexvEggIEZ//02jxPppQvTctP6vuRVgkC1O72v6
33cUsMFDg1Y6ObVljqOgzP6tm3B96MS1OtlylzANo0L2LLb04W4OJSbp8oh4tUKp70hhDPlHd99Q
yguP6047hYmBBxU9kwyN6zX0gWPJ75Ea0fk7KnXlslP9p2Q+riviWHpGNQCKX9Ca5tiX5Zcvr5YU
ToSmI7hT6tWD5Aqy8DXAJFGi/Eh5wuG5hdbu8Jivq79yoYye0rKairaFikmOxd9ExoY+0eIbWJBA
AdF3u03HVGGEv6/4RhzwLFi8NCAaQKgxMZd8chx+zfg7DGw8YCX9rFl5bP20Kk6FAdtWTONeyYYh
lcdS9lCXRlT4nTdOLxj+7osBnUe3xliVkIIHwU6WQPFuvjwMh39/tSdcgkEKhfDYa6TnDCwVEG0e
0cSG0jDtY/W+Vt63zkzXTpEinN+hLu0LkFZBXGOxRfvPm8AxEqjyvUQK0hQPWubHOxwQTNOvk7u5
lBu9sW3W2Gch28KGQWDbtfoh6G+v2ty0j6xJs6SOf0a09qDp9rS0LJuTu6RwjvT9EyOnSGsJ4/vW
RoVr8JuqxurNyis6ckPhm75TwLJNYsNR90VfaLEhHxoqwv8YrAtebTnMzlDUc31YWrsixntph7Tn
XRcUfVAHQK+vd4CFrLGfqsmVPK1TPKtnlg+T+lpBm+IYDPBmfjwF0LPiNMfZvHZ0dLSYlmmo0FLP
TFTb+gvQ/89H2JlQMrE/MgkbuSQab5cH1VNMZhUZRaASmwY6f2YaDJ52hDkNa3z6iFCBWksSXRU+
FAhmN70Z3lxIbqsTe9NLHg/smy023j0CFsQnBbWl2wqivaYx5xM4qZJ0jZgXhb8vZ5JCAJQZyEN2
+nTAUbqIxPWeiAhVu5lJhd/Pxo13AEwHliYexTU7JKdcIOp1OE7wg26PyanyNa2q+iDdKOwLi8xq
5etNM5qnq4g8ymepwMOztxvPrCObwhA9dnIhE5SpvAzAnrj0HUop1QqweghK9aGQEZ1ymprfPpH9
yF61n9Emg6odTFTnOmD8pM2AKextFXk+g+YgF3ocn7aCwnZrjYYLWJDD38TIyli22ExnMT9Cygex
+pQp+IQZHT+VzLpmPXKSaGrKAU65j0kx0WK6rVnbJ3hUmu9CyKuA7weC9T1F1nM/HVOIayZ80qIa
LwhpVtUpObi/w6B5PKDWTeQZEPie08c/k9x5LNb3LTjzGrPHN8F6PVpfi3Nw9wOmDxRBTuTrC+s0
grMiW2gn3ZErdfVYr2S24JXzSRRVP3AZbBVEnSl52r36CSwahB062Ny76MhxTkp+ocJQUNc9u9/e
I0GJFZ8ysANBPUH9U4KTDv0S+WJHFVsqTmz19Vc3xwzrXl+StEm5gScMyrefDnL9XDIFrX42QwAZ
Hr2T7a1oNkj0awI/i01oA2rfnecI92da4+1/gsZf9nnpUvnCe1KiJYsDJB+Ui2wcUgg9zJbysIOK
W6OD23XZcBoNwQANF11M6R5+kLsYX38ky9beY20OIwEg6G3KuVW1q/4XDkIqb7IjwYKRRI+nJHpF
mieWh439aF10HEHRwhi0Qd9nTBsbI7HLjMnFsMSy+hIuoDKFVpKrsvTUOa4FMEeCKwpi3KITnMID
0UvC57otLNKq2T87z53gXSHCUhF1CLNT30rtBfcDBXvBMf/eRWCrHrpksFJLjzQtikr695ULP9Iv
n9rUeg9S1XJ1o78ozfD1o8j4b5W+U+94PCadGoErMxdAdUuJipjX7pYDwvhJPBWJfIOvX2pICtUV
j05EjjoYM50IipzoRtII0JwcpsrMC5B+Axexp2J4oUUvDmKWAJw6im1+fLcwglukrjEoNXdleUNz
gIgCvXOPPsDV7SFhw1R5L6dyfu2IU0W0xM/mxqUoJpCj5xa7R6ihEhB5VjvTEGXxDHLNbI6NWO+v
z5qR3UubjnDB128f3y9aRvj5+WBlxGiykZGNwysFBd+kyPG1U8EHUxIC/We9TVultZXjcB6MGWQd
IusTWEcF9kEOaSlO6Nu9HHRhIIWulEhMI1xbRs9NGkWBGkWuddEyKXUc6GX9ACnngHk47BL/WuWG
5/htBwUISCTlnK9MpqcdULM+9CTej/jC54/mc8Sxpe8jPwak0m9MkjLwA3ojweXQiR7qzeNjaCuL
kj4zH1aTtPuIHgvTkg45J8bS9FWN3WfhmXQmx/AnxUhzdY6V9M3NOT/9yY/5MTKv64WUTCwr6gzF
ElgzcfyZEqLvhFTJWs4HlB9+5RsfDwfXXLbecIQabvLUm22kY6bI3AvVRDJkfUHLDl+d8UGELn9f
loE/p28uz8x/TckVVI3rA8HydvYISh3VzCQOaHngddggl/GDcx/cs7jmTmlyddd/JIEphxbnsLf7
DkB8TzytLQBjih3d5O8XcD/u4xXp5+iU2jQpq2Nbmsfm1KwhPR9ozvuuGikV4vhTxqfgfo2mVwsA
yqyjve45YSnVv8X/OB6UI7HyUt1yQwLAGchkUcPy09lHmgbkP/UE4p9K+p3KAsistHtGpba16TTn
Xp5muZ5xjGd0upElhZXXqB0KjQ8wK6j00rXuLd2ufgx1HkB5wCeo7chcUyeaOvTK9rzsuM3JzmuF
yRXMTKkRjSUT6LrDHzfUGWafMKZlczzN4E0wzxvYTX/pSRMmT/4KR8tqA+BzJzVBSvvbjRgPYe4V
la6Q72hh//bBOCKw6GS8BNEx+yJDvYeiMGMwwtUPowM/cuf8grTpdKf7MC2Mn5LrCF30iamAwaf0
EjK8aeShFTCDUynKYslfbHWbAUuqf52ypQi/Ao7lWatGT6y8FseR72gynEPQma/FfC+Ft9jd6/Aj
DFF37+ndWhwwpJtA5Gm6h4I+wqVNq1nXr5m8YeAKPpbVpa+r7kaB/0C+bFzKF8Zrf2dxh4SUVfha
trUtyTwcs/9yq5O//0v7IBKbOVySceUq0N1R7Kn7XBJGiueH/8V53Ttcv8g+Flz3xJlnMA0bK9dv
Y+TrBJ2prwCAdrg3Dm9Svxxd967t7X0Hz3mklSSFw2BkRAc4Fk/xuuWPPjhS1o4pVA/0lyExNmsb
7/ait9yr01zTMdVxVxMUb9OROyZOPBQonqPhwiEJyXjqkm3isc2zhjNKVO5F80Ooye05xJ9tnR85
TxZuA/S09aTGnrOB/4kcDf4MOZ4NUH3Q1+D5ZQK5t1T2L1wmTnqZnaA3f6WpOJFfMGvFZEcdUgK/
dolv3QzeHa3JCzGN/XxVWeFJyk19KDj5KhxyuvizzMtwjIdpNnMIYBrIk4/+L1TItGp0MCO1fGyI
wXpiiwHLUjv90tEtsoJF1UMw8n8zqbbniruDEpprVVmWOCNY6fw5LXU2B2jwPrmViCSuzuDx9kgr
Fqgc2qjSPlMw8cQ3S64XMInSQwnAyT6ZqENSY8UDbpnHHD3i9qn2sVnQSkRTYBlobcMNF4X10OYn
HVlN2LMb/gzD3qappaTsGWVU+kIfq9gL7Mr6uza/r2ut988WakYEPlB4z5T9xFEmuR9GhBw2VdUp
B4vWhpYLWnos+ns/MLRmAn5KN8WTuXebG0ypLy5LYUafbg+c0v21G6FTC6QnMySgmuMC1V7KfRKl
jkj/vbmV5e3mbPymfEvFmhL+hEwjHEgkl8bupOYXjaXdWFXrsdYM9+qVR+VoOTH4Sfh8yh6uqrJW
VqlNOYDF8y9b+288jykFzUr2HsjBBIbBGgJH80yCf044qIuXG5evd8soSfxR0dYVogwljI3W+wX1
WSkqQc6DFtbe5m/qriJKCs1amS+Y9WZgXQbushax7gWuLWM+D4dj1erTSnLhOjKoBw9XbACDlph8
NBnRI4AW2m0Dfp+f/qNVuz4rd5rxcdZyDNLlOcqDvFN8F0yPn4mGiP06MGM3CVm/FWRSz7sZTYuX
7wmqtHuvx+xPq0xVAwOEv/j9yGfOwh8ngHvQLTVbBmPllIxizG0DFDMGz6GPk4E0LnC2mIypU4mY
0LsJ9aT3+8+jUoiv71YV/ywmlIt/2x6dJUC+v4Zz3g6uMwqDnjxVP1oK6+M/AkLdfw7wWsnPV0HI
0U4fvLz8RCwgtSXlebynqaKu/Z6/AM2IM3D0Up34Up0HIDxDnqamK1qGYNCbhDmRKsZ7SvUtyvoo
VMT+Nij3j+qFuqHUWuOzQJN9BJDJzyxDe1TULMlUQH1bZ+dQqi+ibd8gajtIw9nIg1/2E6MjUbc1
6mNL5C8HQD0K4+MMEgZp654iNVxVZqbVJTNZMmMrUZodS6sd96iFhTiACDR8kCER8F6DBZ/7mqe2
URLqtUti5dJ7eQgZSqjiSKeSm8Us3EBuQVECMwVu36YFFPDtLBsKP1Qv7krvsCNkiCls4IKlpbUS
6aw4QRS9X7Fo+x6NORHFJNywVJmJ7/1czJ/aue379TTOsidBNgkBT358jD2vRfvMAwxSQmFm0+tw
Dxh0Dga8CfLrUg15X1i79u2p2C1SQkBeh07tUQroOteknBwlOJnEFD2MEmeO+vdePQIQRhZjDTOS
eEbtDE8LvM2v/H9a6JBn0G0cYhACcD+a5FfAEnQs1iPCgAJaAZKxhNPs+bVL//Q1xX2XhtVqmE2e
J3OpQKhvCekb41e3MOpzo9LRSURkwugUDrY+4ZAax4vE5sf+PXfBKGjGKst2bqeT+2PS5P7mil4h
OI21fRuiLdcfO/Rc/p7ydSXdK8kBKKNR4vq8lhT2QrRxFExVHN+1kIq0ZebG+me5NHQsIGv/kJq/
+LD8ya2Htl3Mzhx8xoIlek6HoTmJb4JCUqlswi0frsO+7NfBthzR5Qiv4PppL1jgvYm3EjRN/Gfj
fdxRLmtw/MRdbQDU3D68F5PKHOlzj4UxygkqBbCxIu2d4gsMI3h3hfCy33cosapZZ6Alw8VXRV4O
mvWfpJngYVOgzlvwEFE12d/l3HZBm4ypuwh3CT0Ex4P1fRVfw8/8UNp4H+Iu0GkBeLYZnWGuAbOo
0Kywl2dvpZKJb2pcFOLC61JqB8fHN6DGvklrxqYWKJ5tE6e/w2bpSI/HLC1XevXW4vlU1z7XNWa4
90vu6NUi1abjPOAnID570K9T9EtRPewtumMjEztddevLstJJJcTv+T3ab1+0hNxSli4rTMdCW+vD
Pto3hPuZp/q5E+iFvp7vdzmT2DQ+K4rkwumlTMfCj+c77tzCHU+M0GJ7kqnJhCgYwThBdIQuNHlk
+MKDBb23r7zC3IUCZUnqoXdDyhpDKW/LoEBikVnbzuTaQnYkW+swOmWv+7u/Ol7lnyTIyKkvSfAW
Zj0f8QHdURl7fC2rjQbGOtV4DgSrkJb5BU71QRlnn47iwzFMA7AhAk50zBq94vNhBv8cSVDHAKBE
VZfnesS44SMf4ocUghef8qanc6q6pITS7EZo20V6NRRhWHmC+Gs/8V8MVbKKYQOSUZ7v/H5xruvy
Jq4XqXvF7n4ewpUO6HfOKkMvHy3p27cPDKTMNFDGEDr4Te5mDYpE6sVp7rmpXmLkI4XJ0Z/Blxhr
TSOLSw6AkW5XkktVLy+MyhFaJYaqKtqbEtsqwygpL5p4BfXI6MYf+s4QVHuxO90tg34EzkRadZ+p
DkDRdrHtekzmNJhXPf1wmuU/ic74bzeWY1NNSN4gxXFS5icGgG87GHJDlybDv3FysJOUdctV2Zjt
JiWQ9PC+NKqQilF7CuFEdGGD2IZC6J3hZJ3bydTGxDQJrltWq30ENVrBXN1jmqSddbRhBlbZp0L4
YihLvVn4GICeUMMEXT4qEMJpOSqP485uMt7lMf1hbTMLWM6kRhcZwlF2rkINtTEI9NVbrD8xRJ/l
EfjEwblxmphK57slUdIFfqpmRxc3fyWxGos0REdIEzgoho1DH9yoWo1YXEATH3PjZA8N/laUHBfY
DpyAa7Gf0n+tbiCRz//6uuA6xJgtVbNmsw1TfLa1kTJYtT9M8vHaT2W5wofan5oA/UlQVjDvMHCv
DNfwznbOP0OkxbrRxq1ZINqdQnNOy7QzZNWOCEzhg3b5NjSIjxIXPGY9DhMVou4YS5G5yKf0co11
vtBWJI/xMjiL7TmRzjjZ+5cyjONk5oixH2XpECmwf0rteieCYXmRXwhpwoBNIua8prW0vlYhMXTU
She2nob+jhoTt2X+j0t8eLr6X7J98iQDT5nUfO39QSusYtfC+F4CkxtXZ/1QQz2oN+8zoUXRFR8T
8KdkRQqfFkwwkG2xPZcr1xXkcJLfspZ31FJeNF9umsss/MCafqCOG4+uLxz1qEJj+oHPB+o7J7wU
VtoMJDBT4dZXqz4GiypvYqSs3Yn83nQq5qlZkTYNEPyR1zwQ6h9riHIOAzrd16bF861zMjmDUKe6
Yq4KJzZqp9ufq7RiaCiIXXeU70JkusI7I1Dv497dnWmdqvaDZdp3Xe0FkMgvZF1yLsJiz1lKjm2a
CrBzHQ5hY6bOvD/Et0F1JcMsouJpqEhXNhtETuW2Zb+pbfMu6/f0MWhlWh5FIx0zSMnO03tZtrDp
3L+KOCNcmz1a23R/0wSSgDVW9Yl/2VvZ5V1YBxQSKB34nJI+c/TU45WkkC+TTN/SNCNwnSaBt8bN
NlMJx5H89Vhq7M9+pAlX1OaC/7MdPviei/vQ/TcN+xnyKM77BjpzqodvnimUVL4Atb7mCU6qPm9X
F+cY5MwqeBYbZxfzaTly7MLIJ6J1LymoOI7RjFtEEWNjFZkXKiGr8HLgI4oC/7wr+5TBSgUlBY/Q
3A8Js8EBavrBNl2TaceGuAtepuRyNutQAGuV6WdNlABRI/MnLu7e28UTG2s+uvGeqGLBi/SNv93H
66Z51VMH5PXUOFWKtolIIgmNpd3PR+aNA3uIwC+wuqxIwVL+/7TRtn3NhipPtnPnViMZRLRoiJEx
ZxZvHxkfmkFs1NDOsOWgLZ7EezlBsaqkNMR7/rZnOZhXP4Ufsn+SsrPTH+CXnRi89p5GcGto4vx9
f/obnUAlq6UKewnp6RZlAPOelaNIqBmiDg8m/sJpq+PNHxCJKgk0DCeIRc+W9Tlih2dZ5T1Q9/wB
yqNrBrllldxlL1dtCWsYKmejnqobEkuBVzbYBnMbnTm5Gz8fz3iYw42zjwo1zyZduyXUCfFwo0oQ
zxTXsy6mavV7B8zCj2kPTX1mI2mzhYmjYMUp6DJwzJVU90Rzt0RzvohmbEYsJwHhoMjmz0X3rZEh
8VNaRdl9Qr+KGjZS2YwG9ukYRMWQQZLN93XDg3e6f4j291FopqmbgmwuZmqVj210ipjLdcjvnkOH
EcMgHrP0KElhEE/bSbNGjxqejKPII2oMt6OKm8JysQifKGlKax8lRf/dlRNRMtjrSUYA8tvjEWs+
cDlfMAvY7GSYJCLgx/CrC7M1AI+7nmSRoFRz4/d4z1Wf+OYNwB3U9EsnMEdmxOvfMBGRltAtm5kt
OPrsNXKOLMoh1JQMHwlL3gr4GJ6TulRUb2ITFyahi7DnM5KoeWbZYZ8cFbA+bPaAKzH3DOd8OTjb
5Sb3505nRyYWD4YedJBU1I2uC+sQgQjZ0tQ3pdt804YPNrqN30DpUL6Sk6TMpoTc7jRoYVu6d1xv
SaXdS6BgS41dEveSDHwLN+ufjut5R6r0iRA+Q0XLBoXDBQASo9izGVg+atVPL7xRSUtS+jrff1eB
AAmGjRdCPL3LLqlHeWlzJMsfj0daYkHajbSSJLyQyCfW3RyPLw3uRCSb9qhUN0zN6PJxyEIkQfvy
ZmA6+5XZsdwiokakkZHHZMMauCFc+qzdcebEOMHnp/Bx4r0AwD5XkR7f16xWrPd8n4YBtPEa7CA9
zs8sq/aaz1tHhbbNhoOfAFUuk1vHpqHo8EM3JVWpwZkB7BMor8YsLACnIrx7JKvq1upN22oxkUvN
J/+T3SiwU8Y4HgkKZZaDr9tZseR75s+XsQP3BaR+6Frg+smUhlBp2jg0o+/EAoy1qcdeuEI8i9/Y
fQPu9XtQ7V7EdJrvhFeo5ztQA1XgHdQI2NB5a4GNi0kAUYNPOYfTW7aU1i8+VCNRpQdSaa+pjqBs
0mErN37jX1hnmCI9VQQYGdjZ1tS/AGwjx8i/10EssRJ5ba9QoNVXDazrC1n1RLVIuY0AifhoaaEM
pcsaTs8FGBur1G450LfrIUBULt5mluEfkiFMzzFrGgP1fkc/ql3gA2Tpjeo3uAkfXWMWGUKd1aw6
NKYP+Gonm94buVDjezrNcL9MIEpf3vZ40E6RgJwHdo2902vy3F5pTUOHkH/SlOpje+5Dr0csu1fV
hSMOjSxQk3Yp7ZsW8c+zFhjJcGDhc4KT1diADo/W0T4aoG4JSuoc+Rln8eEmbFsc7gZeDhwCn+/M
+nrM0vP/WbztUmN9+KRe8dX6alCOm3CURudH8/iFVJRKqRCbzETZ6zCvpbMMogY7xdtmn/+VXlXM
vFxk5WiVbCwnDVpsM2tDfwHjJ5uiGNaqAXAHTWEY5aOSk2WHqK0p95U6KPM/BnjetQI9jjzw/Rz6
mdkz8gITePYnYWWH2ATpGcGS+N/mYRI5/bGe4sHhtqUXn6SZkb85pDpjECxIA2uWjsjRlS4IhrCI
DZvbO71yZt/ixlJB65S8N315fH3RBkv0Uj0M5EhXJJSBQH5fUxMEDG/9mrZqv40Clz5W7mjU2XRZ
IAtt4IcjE1EQM8oGpX68XlOjTaOAqePFcBUuzVlLuuMAtsf0I4XPRoS79uFLqblV6co6WQw7BcJt
k2Ff7ie+r1ynS7sVL8cgoWrxHzgEkgzHPl6dZ01pBbbHrWwMrYnXvy3OfTbcdHFhg6J1s8t+Mlwr
xyvpIAMUqgDFswhPtkXlaA+MY3L3uOKmU+hAQ0z4Z2DNC2rEt+1RvBh2bAn0WMPz2sjXhrE5OJfD
XFFYm++g4U3qa+ywaH7+SjE7EuFoBJtQhyXn6HChVvxKDHyrU6NQq2niWG5y/bFaNQWoVnBihunN
FfNoXXntoZw6ivnafFUIhPIwfIFD33V0JWIGW3J9/vHokhEU+ad+W9uJLtvrZrmWb/FYmCWsTJMt
64Qsd/7y1sgVsOii0qgya88j47bWiZTNvJFN4evAyhpOwOQc+Ydgzk07S1/YIdensIY3iSrVxj6+
IQK7Lhwn4T4tQ7nCcC6t6B/Jj1lVfnxwlX/5QbIYzrV5ZfAMoUcz2IrKwzv3LCg8fX5wG1A71ypf
6OmvR5tPWeoGgtk+y19nsqudq/FHHPHVAgAXfg5byJKLXNJsVrE+ggYB/Er/qzF5qGx4plgaGdU9
zYdb/35o/AyrSYpQT+tLD6G2An03YImkobwaSHP9qIMlK3tI3SkMZqsKcXi9PPqtVk2zhIO5x7Zm
UEOFW64W9K0GGeAoHcH0c5vVuGwAal2DejD78T66oOp7jBFGHxL6cU0i++acMPCZgYHCHnQ7fCHf
qS2jxZzHjeBsb7zZ7N62P9YMZZjsn7uU9Q85a5xq90ZNdMi6qBf9vITQBfwuKBRXxXeVRckisd1M
pwN6M7l8XvEZV+iNBrqWqVB4I1OXLznieVw6kU57FHtSP5w8VBEgR+KYPT0pmjKM0ZonUmlR1t4d
gPTC9E9vMLB1NuI4zy37URpPZownMCaI9Vkoxgm6Ntq8X4UB4QwLi1xKTb+ayE3nHKIY6UIpopu2
h6ee8N+UDC37sOvg5btY1Rzr2GKAUx9Pl5BxsbWd3PS3JJuA9AzCvjQn7eWGjsYJOw82ZL+fm/Gf
TDuDNVNEPitgmXYH3WkQjqs2imiVJj0iYyZW36fQ/Uukj2FznW+cyCsdeSctUvmUjhKhPum+oFdI
mB+03ozBimk8pbDty4wN8vm6vBtEqlgO8hZxCrfo6xBXykN5Z7pvQmwFwK4hWl6787FOuaQw3cME
g1/9gqKbRiI9wJxe4mcvYZW2vpgp4Rn1r+QfCHOxJBf0XML93YjHS46yJVy8VeSvrtWVK1Sp2Qqm
RZgrqKb4Am2T+nwQDTo2uLmVyuANUlBrOoUefB8qVq8Qc/h8x7wkKxMb14QLinp/8bXURn4AZoVx
thdHHxvvBprGnwBlS0OwIQ2nhkUSt1eLRZZxCk8RuoYQonXC3DzQWYPvFtJ2/1NCqhr2b6Yxs2DD
8yVNg8jFCHTh6ZhRiuBZ8jXbADVofpiycpjr6DNouAj26jrhMDk2w7Djfp1pQCKRwb85jks0KpUV
DCr/CYA3AzjIeE5MILB/LGCRgricLw5KDKY9uaQG9oig8sLPQclJFDQK7kSV3eaaw2Y6hQV7W2S/
ok/Gm1JTXOYGvIMWWgdpHpTdU1FmrKk1zLyz1bfjHDXqaE6dtj38s+lqNto3AMDKYdBW64/llyPh
R5vE811aur13au+kd2TQurW8HG4rWF1UhJt+07Es3fkxoxaOmZg9wcTx8aG2Ww0BvyoUqXa+hOSL
c16vWxFUGvwIc3/LAPSdn0QzyzIHSdiaxGN8CKqfDndF7LpmAhPv4WCXQpA/1V5UArDgrdrsiVDS
t5tRZvlUXg5IH8nvNApHcCL6E5IkoPixEYvwvf8ulCrAdTZNg0B8Wsfo1Tu/ekad75musRswicdm
M920avF3JE9AfCC2Gh6EyNkbytPR4/yYGwurCGzQVs1gq0Oi/f5mtsemlWU0BKH7KBVOWn1Ndlei
gfIU2/NlzggHTgqmMBp53W7QWmYzmg/xKiYcr+bj7FU6GIr+4dB6Uz3g9FWoqGlCAQVIlcXG6nQP
0HpdotrhvJEBe2UOaFJdsTgoUwtCcxSYR283gEKzmjO2Ns6WAmlzVMe/wtPEESjjHcsVEGxAI30P
omztLCvn33F20WBawobhRqr+9hic3yJMmFUugQD8cTWFEgpSaURAa+iyvP4/Bl2Pr0Z7Vy4f9dPf
OqopGQhghNHCtgLIhuT2EFOqVJmZqmd84gKTV8gDige6nlzujVTCu25+vO3oh3fHLwPun3QK8VI3
+eGL8iME6H1hvZrZO76tM8sbGAvVCHSuEPK1LkrNNs39l6n2Oj3T60K8/uUFiUYNOPSL/JtDA46l
MidhKXCbcCpLPGvyjHpUOMqKB07buwHX/IczBrp791p2A8cSFsZUJdGyVbklaoLV/gwaAzEifP+4
5HbhnWZXdTTWyVUwuqeoCvG01S8iHSRHO5RrqiPiG5v2baEG/y7D6Q3yPnaFikmDcB7JP+Q6g+54
ICQr0PSi9eLfMu4yg/D+jdzvePbcIA4aob9c087xLyHtEWRb5ww2qXnprzygFKaV2y9z1fIx4XQS
UQmNEPsWjYMN/VjG10Jyv8aSihMlysrJQ1jKpXcj4xQXroMXa0cnvP9b2AoqHL70YvdtdN33/FL8
/wrXSpTv+jAfMKFP5qByxXEOtdaZ25+NEw7TAeJGzV1oPUZ6yUJ33pTokZdLLv0IrFq8i8ReQcEj
bwD/Rj1s6PSQodCAEVidSAQM1aWClPFU45BgN4/v/YRlU+YQfoCKUhYnr2Oxt4HpG7o141x2cRKS
Ri6gY3xk/hTGmC+EJuCEO15pi/GWkZIqm58AnrDs475Fhf8k2syI6V2AHxYhZHgJKDBLj4ta8WbI
dQ28zcsdtZQWMppNuwGj0DuRiLZbv0cAN+3YybtLGwTGUwTG/A+SRQSkkf4z2Tx/0Pux0IThPYoO
0B99It7fT5cxEHu0GhkxezTOvChz8aJpaAJIYCVas6TRSPBru64TytA1xrIyk4UdrjQ37huJmN4+
6v1Bd1wKF7f23IIaBDsYZZxfwdEuoXh5TbmB2C2LSQaiQMSkUzvreCQBjhAI4elYFTcArVMu5rfz
k+TXkL0nJ/uItBhLup/qBTf1HENX2BYgoJWl25r6BQKcfxcLs2Owwozi1uIfutpTykiIDB5GUhW4
eH/nbWFu3inXZdZ5DmfBmcBMcI6sRaKIDxtlFRy7rh9bELnDaQFoKfGgogWbvzcq3jKV6iKQtXAg
nJFhxhP9tRXF0D8xaxfieVyMC4vfwqbMl6YwsxEGBiJPLwQ6TFwLxXNMq1KJ2TZ0OlzsotAhAEUM
rX8RV+UYcCrM79Xbv7b+JoWLPO5cMWChmaJhePBfyfE4DICZWZRYbIjU8mMGl6Dhlc7eqktzBpR+
+ihb8mKv2RP+106i5pufZSjFBQVw7Hw5OZJ98GnmnzQaHM74gfF2VwBL36dJqrSIEbCTWMcUL6Xf
wvKnXfUDn8RvKjkQ+HKkg5ImdJG7J4gUHXYw27MlwhXzuCSz5EMAtM2oJnWEB0WsYBAuA6r1LNoW
TLvnUljG7o9HV8dTDXDR0GTr2GhGf7et9PdkClfoEeJ+oygAbgiAjvsc7QxnFKKh5+k2+U9Nihqf
zYanh30JMPsfI15m+aAxWXSp37lUVFK1rahXMR5V7UWkzIv7uYa+gBm7LSwrpsWRToiJL5++OIdR
Cdt2wNdnd6ef8uiqAZebRq5UK+A5fnY5LPmiurbArUJcVhwZUS3jTQ8Ie3cr0insUtnpqJwZsBmX
tjzVx9r+9svrKNh5eBTU1yO/gOUCxQsMVAYsQ5V2eZmudj06Yo87Zp25/YQWbleENWbNb3qHJKZC
pymH0v6Y9jh2/zn7V2iSk9YQmAcMYFUoOozjvwJaDszX9KNmnghSUSi4wk22kjXo8AKXqYqbLiuw
IfSLzl2KJlJH34DZPBNFi5mIaS5UxWxyxt30yN72pfv76H9dPIOMMXoDwtB4QzakzDLDefgK2CES
8dNYVZYPVH5eZtDe8znv1ooKepYwkd9qrjTzOBqQwI+muWzOyzHXNJuJ0AUVitMKu2iB52Sodm30
JzH0fyAbnK27ab60JH6+Z0O2d4RcTKB/8bsxSZqIWyuyla+r9jOzYU8TIIbzZrDU8JVlYObZD9po
EbzNW77g9UAOZ3adCbhGinGrpbY37MOMvWKWRGqn2Sa0HYyvjt7xjRPChxuzgxoYWHDxpdVXnUFb
wHlV8obaKMyU47Gmo65+QA8EJyJH5jPuvpWssybbib1gcRj3sc1UKfOYkn5sEH+nwvA/TjSmENfY
1iHOnRgw5JObRCgXHmyNi+DbuCN8xE70Y2xLSmTqQ0hOL/gxaBBWwXnMQKZk7dEcCGfqesCnuzXy
Ubtgcb2LxVsn60urmkt5BwHlFoq1MjnUXliP9zmfZtLdY9Tk8dQobiekenPoRVo2HS3JoJKaVkrY
4hBNrGMclQju58Gwa4UV0EMFTqe0jUuzzvfBGa4HzqvSTRySh3WAbCtxABOL9Inj82Mi9Ekm0WYB
H2LZmpgVtTgxGRPz5QWFHWKo2aTC3aaIMTMr6v8tEKKbp3KyRUcUBy20YizyTPs11FX8VjPV26qj
zCZjbeE27JWWcUiUeiovxfVwXRQhXUtADnmVUrbEDxs6c4njiM9vC9czB36lzieIudAQuUMMXLCw
fpByHufy4ksZnTIccTdC1YEX97go+2CvNjXPX8VrxF6Tee9l0BS36HLiyHxn22FSRVdJfkIxojyO
q8Yqv9hfaC0rqzPNgTBMqH3HQ613QmNfFbuaNpjzVcBHZTPgDlJTEdZllGDseGOCnYxsDc4ISaN/
lBte7rKOx16efd5UUGn76vY2DLrq8fLvCnr2szCjGE7o2VQck92+nfS+id7/N/e7CoXXr093u7pD
GpxPZbOgmRXN8uK+ybI0eE+FD7O1iBcT81Fa/lShWXcYln4pudyCY4G7o55sbVFxozyFcawrjd0l
d3WuT6eoqjAYGsEd/4IACzPxaZWkriuTHmR3d3uE+HvFQZOovDqsnvo569oVjBwj9IepFPG/UuDI
XgDfpwSpbDHp7KzkL2GZ9aVNmxPsZxKh1dX80jV6Kqg9bHkEjTDhSSrKwNj20Dtc4E7LL+3s92y6
K/z2RGP/VHYvr9WQGblmczvwBQc9vJ5gzwjkUqTrjpXKWurzKx65nv1ZRoslswV/OrKQHwwKvkn2
0wsi9fz4sxo8h3ctHlmQT4kvGVljvIXS5BlEiwrch9iFcmej8ttp/k4605tPjhdBgDjCuvEvP0hY
/iZtKUYrkwGcKhxw1iTW07kzqdG1LvC5DFv8HBwCpM0xCS4Dzjed8f8Qp487F6XTGeKXScIgtOx7
yL/QiGG63rgdfSFqNpwvYuuic/ZNMxOfVMkpN0j8qwJgUhrdTYzKVTg1NxCZto8PkZ2y7vtg84xo
FBguSN7yubWdycqHh43djiC55dB9k2kSxiJW/LFhtb/RyoMXv3mgB+gFeJiwYaUcpcMawGmjyoQl
I0220qkRETnnM+qH9QxHilf0zuq+NTyLU1by/dAY1rLa+HNPPItQRLRZyFA0Nuz5do3LVtBVXKa0
Me26MY+iCFkW6h1qflj4etqYp8BUHHmUHe+WTHrzcMFakNFZRfCAHxCVRXl9q2j+Rhv2b/29hqrP
r70JaYAMmI20HH0GtXFjL/RCdVqgiV+kTeynljzuHaL5vGJxPFZr6HoS16JTAxoOCtFVo3QwqIED
DMgtSUC1rgtVafmHOc1MJ9BWHP33GqeS2jTEnX7kX9JjkyfpGoYitQ0ol8dnTpmnz0q0MpINR2bZ
b2/H4CpskIxaFq8V5OdeC4PcQpesP9q8wow0syFSh5xciqZT4YiKmfWF5wW26SNfg0NafQT6zC/l
wvTGNU9DU6RCc7wvMTogrwsKieIlRn/wUSqdo+UOyv1BYi8aLB90r4uUsxAIpdU7ecp+mOHoe44n
HlxxvczUHDcm1YjIt98KyzXtXATSE5c6bn2XW+AraKvI9N3M7wvHX8W4sMjdH5YvQq2eks+pqAwv
zEBjo5TfZACnIM+qevG7eDxnzM8eP1GW+i4hb4ZcyylNKx+StSThEE4cCAktVLb4e/dOviffdrTY
HqIX9am36oMmE5HmqYEsgjNTm3ZyVQyN8PQdT7UYWI+6RPxajut6TcHAANwoNgkSeorv3TEq44E+
lRYSSpxAsikFecK8EdGQf9/C9Vo9W9Bj16vKFKGuUoXscIOiBKAPzshaCWZ7322/MfVrAl5foKF0
RiA9OO75v0GybLShQgt1koV6KyNkg4M+CaGdkq0Ybq/yDReOebkOztOY0AIzzMIVd2/rpYdBByUG
r54x27cFSz/U6xrctvbVbxRRVSG25CDLjW4lvLeqxanxbt6CGLL/23xplDK+ktKVqWPjSKyuXyHr
gsFZbPBnwr1WJB5ntkt4lqzz+9dsdRyC++IAhw7r+PpuhE2kWw+rB/yNIe27NPOSHpKnO+ay210L
2OE6DoTn8Tikru8PZg0aSVtMSSdOX5fDCQJjhcSMv+/MkIfdcVtxVZa2zo5VIhX273qMQj65izOc
bnd6pGR/WAWUoOBAiG7xpRtmqTs5qx5E09pT7pwCBacv0surReSRGgLbYtLLr+SDZt+QfspXaoO6
Cye67ZsLK0cileLVG40Z4i5eugnHxGYRBedlvgljLO/cldb5P5cMgQyYJh7+9A0SMdCVOgzdoR0F
perRnbStQy4vindnu9QV1eMExi2tVAoWjnrNATjjJsBsA/7SfGcxVblYZtYNq32ItX54VNZl2UJz
BEBBN595RZ/lRkyJ+vMYP/lJ3/UWMTsTWfkRj4v7LI0PegoDxOKFhNcNaf8GvtfYpNiXM5MqaNUh
w96aoPfwuLruIZtZ+ISSmcagFgkTP0pA+h39G2u6zP+5U4bVCXzMRYF8IdyNosuZya+bsw5DE7RK
+4orFXa9N13p7vO1+R/X6ao6P1il4/+vrw/RYYdBh5K9zPo5ryf2VGTX+C5AEZ8oDhALmkSVaKWi
OGGNnCTrMXWJ74MnR+cTQ49dYGm0Jf2XN4IZcWSLDysDffB8jT8SUclK+Qm2aifMEYWZ+Lcg6pFy
Ui0KTZ/gDzcr8BSnBact/7sebKg3OAfakKnR1Uq7aWp/igHFU9KDZrIO06FRuvmCUzR+dK9wXS1t
tmsvPmVA5P2dxornXP/VivyApk0bFYKtyFi2GuYRS/Hg+EtYNUXdB/S+LFuc6O5KXUt1IR9ZIz6p
iTSq8QcMtv2/y3VamkO0gxmJ1ZNmBLjiiE2msT5hWqmTu1QxOk6RyBrHCxLeKqgB5MdLsGFd5CEm
PiauRJDabkC5lJ0AJATYmbBOypCDhrNDKK1EugXjV1e0HCAgDSiDRr23EIC+YNWHzJslc95aUcHY
IrEdG8daO75ORdL/D6Mry+tzXCv07XFJdgQA1FdMoEg668NXuoLZeivQpuwl80QoR+atD4yeuoqY
g66Nr8GzX1fwLuROr3wJ0HgbBZO0cmoT2tdaAJ90CqndY7dLVZ0FDMN5E7umASEd8mpLjaGLGOp0
iybj0T5CYMJW9v9kFR8B5fZx8M4gCjJe3q84gHmnZ+M+hOyekFyjKRfS8P1/tq2ryCfKX8b5Qh14
HvIEh1k7DKxgoDX7abX5x2cVJ5Vhh4VAQV0xZIxHvq6QFt0RKM3LaXups4hYEsATGJW/mjsmLXyG
hRYo8MKLpD2IyTyylcqDeqCTBgaPFN3I9H5GKxEYYkMdO+02heJunWhKvY7t5ZZQ+rp5tP6RiQbi
cp4aVUI0nvUlAVRoxZxuctOp7eO9ZvTZFt3Ws17WJifvTBTfLD2y0xhM53hwVc1parNKKhvQ/SiP
tfJy9Wz06bdLvBCQB0++ybgMlKB1+NaWaM/OGW+u+3L0J6XSqZt9LI9NOVLobTQmJjfLuKPBsaO0
wciqCVesdB3TfpU6Wq+bhAzO4SLVlahxTKr097/m1E/Jo6wRmO8zsCAn5LPzhg8cmWpLuUDhmPCL
1tX2S78ImTt9WQFLbaj9mQeFBWjMyOS+l84PwCusFnjbUx0HYbGiX3ySPlDvIx7AfmzAkVhOpnfN
N8/G1LJgf1166fzSDJ7mYUBfBTgwO3BG2HoijngiLaIcn/W5oqdJuzZm4tCkUzcovBQf+JxaurQ+
6qKu4uv3oNmPOuPQCvBaQ3EelhNmFywIXtlofMHcbLvwwGObp302PUEKfp/nCxyr0VOaNbn7DojT
pBpY+uSmmMrgtrIhHDwPhK+Rf5KJ0yrR1s79G9n9ITt4ouCvzR8+8Br6eTpaWw7ozPjKsIyfPhab
40zWPHizMomMD2OLZB/oLUQ/pI2Y7OMeKt2Pr0kC57gwv+uC1/Lw4s6cHrqh+Yb0FGAzA5IHUKCt
rZ98ip1MDX5cG9gvnhgw2mBBsybZeuxoyp6jwQoXSUCtPLoeYyt4/EhWhXp0iSuIuU6j5fSk0nDS
FNL1P4Z5w6f91Eftyqb9aGCustHEBs3rNKzIWLa+vllfWi3K9SNzOueMcyRoalXpsXRbxWVdHJhQ
cHBsA+xCWpqcOYVKvY5ILzNtNiWjUVo0Ytj8avHOeKPAP1VqBEiyhAw8Hd1qYdtXfMrOhATN91Ne
zFwkPISSdoYObYOSTuD71MnA8qYX0unE+XoZOS7X4ptpitomIhpfnHwDJ7HiA7LqppctDHchK8FQ
71Qhk3+tiSev34AylbI3qaLlBZsUQFDXGnr5isJKQK6j2jk5gJqFgC8r6KrEJWkoNdaL5B/I9EBd
o7szwf+Aeeb6RPbFsImRf8RZl+WNIRFxO03E4krmvA9iRP6kjM/V0TKpHTGnRFf17LeDutcX3/2D
fqqT+ZUPYLc4gJ5DjV4dGB5P++NYS2/tA756JfOjJUKntkwUsTF5Cp7W7DPhwJXfYlaEbVZ1ESMI
LYci9ZUYtCQXxhaWAIhXWMIiLe9bLcz8bKsa+DjX9XQPE81IeltPYrcyE4RipvryKvsNZolDNdwn
lzWGNBZrS62FvuMLCnnUBJLLxWwP6UlPqGrW5PSive4CrcQQ6OKI3i9qju/txk30u7yLcpi6wGSA
PFNqZ6mgYS4dT0a7LwRfhKKQ5b8AQfrTpC3Pof7F4wUHlsXd0abZKvp/gj04KSL7NJM3JxHB7/nv
zTnqjY1ufYaDBVrbDbdWZOCzbca58gtmkGf+F1xtCGAmbJwWG8ZaTElo5mwNFyIKypajb9MPybcz
TS0s3h71qkb5TRewXlkKCcNF5V1Qkb3TWUewwdmRx9jKADHOfCLndyHeYoh9v0mk1Iyp9V5zaiuU
JUwcxJE/nfxdtgVFsXKgar347sOOZzesL+Lub/JvlOn6vOE/e7FFGhxxxLias74uLTxtz1hYjnwb
JyLQi+HxLL50REucqUnYJ0YAfa/u4XrlezdaFUStL5+RO/GyfdnQYINIcIuaALrHXCqf8d4zNHSz
AO6rbZzjrBU1JA+zYSUqiHhi7TnwfD//T3HVDKqLigJRak2yBxc2Do83EhBlmDqbJwyDqMXZ6RfE
oBPX3EdX8Kn/XH7kffQXkguAKNNCveVYixkpFqGjhokQkcG9bjm4fOj4fYDZ2w/Xl9mfFzadna7p
RtmIXo7Mjg8FM2FNfwFcYQvNl9kBJ63VnxiZ+AnTmgtnMxJUOF2FYIuQpRM8LyHSdI/YhzOACgeM
h4mNCBIHIH6VPolzBm0aPsclQa+BblGBe+gAgHMn4125TPwdeSfwfJoxqJ0XUhwVodid21dmkssm
prltdc67i2ZHVpMoz31zyFALeNBsbIeD9+5DuvySUhk8mjaPcVvvwsswLpTmzaHxo2k17x6R/mM/
+33/b59qAnILODmoSBOCljmFEzKp7kiqdYzHWH0z5wVbr6hKtUz/PDyHPTiXlMYksngLMA4gQN4n
Qic01D7v3s3+/P66t5VEGsxQTe53YbWBAUOj52+xg4NP/tt+Yc3LWzHPbgvzCZm7hQdADqyzEpSE
4o39xz+0+zrdis9W7qiRg0LlPuksoMdwS+Ifj0CmjMcuwwEgQz6EYl5axvV09jZj5zFXjmW0KlDM
Fr49kTs3N07XqIN5NUJdrdJr7LezTNT+PcpHhjajvrDu2ZWUrgqAuEhR+sKabl5C7CoHf/TxNgio
3LfG2SCM38SG79lvVlt5l9+cd6UQF248BvEtXnPHujIF7P2gs7rrXlAD8omUdBqNBvlnRWTasVOw
uZONfZ2xGeSbCyQTzNngn9NocOnqa+9ca6Uy4bbXaprzuBeoy1mcu4hNIc2gU19ZRqk0uUU3efS2
kCqLQ2MexflL67p3tDlSFJZD4n40yg7l30Zq8+WKJ2Mzu+ov+R4Alr99gQ//64P8kl9OZF15BtkI
ApLjguHebCcBPM0VIoZtZnKGAgCoRJhZ2Kt+hRLsBcrHfzOEx5iNuYc4rRApvZ0V9VN3/EcrZ4/j
VdZ8IbRkhxrDgsyKJFQ6IohxwJNbow7bu1XOFzpMVKFSFkePWDWQ58RU9sg+8rzcuRC17kAbcx6Q
CD9Fh5oZSIh8daH+xqMOWoCATwABuF5Yy+0PK/YqF4a77HfPcQcWjgN/wdclsEOQreguE7HxJHJ6
IVK2ao+EHzVafe78I9rrwW1drOV0mkmL2qV6Cj+Qmh8iMP3gYvPobvuwftY58cfkU3ZbYs+TCEhh
/bqaO9f+Fkdi8eADum7Y3c/OyXXquj7Zmem/MXVmG6gMjCLYGWiK1hfLKeizQ2UjtiapuPtXwl1g
AUzkR3SULQm0V2RFqXJXDOOjP7ckhUiantq2bdQTu10rHTC0KPpcCERpe/JZlNkQjPcdXQGhkYoJ
W/XeRXrsd6oPmEoE0Sp1yMzWf+ng9HdpZC86J1qCLag1mKHbulgxw0qdoqQ6MXgsQZcub0R4j8cS
U7Nu7nRDzZwrg51Y5bLMaY18oBYJEuKlFIt04P9j8d9GPw16DxIg1s0H0DvTqC84U3242l5wd4pb
/RwgT3DeYP+kVVtb/n/w+UT20DCITWXpbbQU+2zC9gf10xrnH39DywbYTVwHEFHJReSA60MdhfHD
ih28fJUO6oaqlTe22jvDEX0LSGX5RSLhok1D4HVyxKJOwaY+33Zfz75lxdoT4uZDTefJl5a7fiOK
AvicaP0vAbS/Tnv7gfk1ahvx3aPQdhpTuNncKnW6UEmCrL+ub0zjYB/1txdW2Z+NLc6coPYaj9Zo
pMRCXltX9c6NiICwNh8c/8zXOIBoTQzKxAyXf72dGy2kCjGzfYpWRQ+XmfeOeTFSsH4C5AlFURzj
4yvnl3178GLSgnPp+ZetOALsfQ71CJdFKtwjdvsQErFWQ6X/hYXLdBXQdhJ4+NHiomYa7WaF1VDD
m+3WcXLB74Pz2GQzVwRdHfHqQnxaRQRi8po6+T9JF+xighl9+qCZXrXBBhEUxItzGZGIMSHV0FYB
L4HzdscxpC83E7CPah13n6QAS4qjoWx+pImXzL6QzL/JyEnYCHYErNMJOffGGYnNrRsQZjcExNWc
oXnlAPC7P/byFWA1zZ71Q1MWJ8tSFoX997/vKsPaPHli4botxYbKcDXM9Q4RhYyUSA6UAm4Np2fA
IfiX5fFnbHTHRL8CR5Yy1OAS1vf0+dQgDE4aQ8YWlZneIq5F6wldxYLwLYRG8Un8yuLLWZgZcbsG
K18V6zyKLo8/BYljdO7Le00HrVplqjkzcli87RHX8auKKwWPfTPxyyP3vLrlNUnK2P08HoFQOTB6
J2Gf7A/kpKB+XfG7nUXvwel07/tgeao0DEjg2NzrcVOqnbA1eEPgvUFLmvsBKTF2WitW2YBG3nm1
cEnWwkKbfskcayNgK/MBxdJr8UDTgen/rk6ExuBQGVQSDf9KhRTBmcAVQUiNgp+FPFSDT7EPshlU
SV/0O1N1SjtNGCDtC8OpNe3sfuYaHoKkI8ymg4sw8V5ld61f0FpvTXjn6SFniyOScP8N1N5bULor
ayH+xL2lwOtmr30+vcYWzXQX38ybJgV1K5te7tl4ulYKnahQhOnCmswQaXPlqufiFMZ0ikm03qVw
pZVkioBXapRDdBqxgq8aO5ru7wfIszCuuXZw0QFTr2UoAmm2jv6J0Ii1OoVx6Yy+8A/2a8qc8Cpr
2lSCTio/PyRhsaZUTVmlirPYpCPkyXHn3I8YNhwUkgHLh1RlQnmG+v7Lle+II22Ofzc225K5C30a
HaNwO83rdkGv1T6/H6004l1s4//KAf2cc3ByOVOQ1MmnVJ2aZR+HarivEvqvxymkCdTqC6fKXeue
rKEKK0rjczF9w1IE09WjmTPGLEQesafSluv8IKR9NAdXmqXWoJV/HIRTasgmuvVuEsrC0/Dpi3vw
i8Nioof1yNPVdnITS6VFMwVxWQFR7CQLHwUnT7v0Vyni8J4uFZkl02rdn/LE7uCyIeBxV4b2TQZx
97BXhPXKD/ByXhZn745r7VqogdQXtVGQaG1ARubqQ0zAYCcLfcDjTt0qFGPMifzY5NsjtVNn6/h4
IKCv4TbJgyQijSqm6Nlz0bf0n3lnShv2k+zyxqZyLwZ4L764Jqo0Fgu6mojKf8KUaoFf+zJeIKsn
ohJeogWQw9Fml+voKFsdVB51eInSsCCPOSSa8IcJOdGXNUgzFaipdBKEgZmvCHlGJa+rkxWZJriO
BZYPdTabaH8Th6kxESB+7VRg+/YUZ1qNJ7EXnxGUro+31MH9aQZUhG4mlCOHrAFXO6NNuLCfzO30
OAr+bgO9EflaHZNuwpoOpJgH2lPyqafLLqyv55eqw2FJz6Pdv6RYauCeJTmiRuwL2fl72588UM9s
UU/KFWFtvR4pBEGiR4JZsJdeIojz/y4ZA8nt4Jmas9jGvvLJdtGVSeaRGUsN+uqphoZm15l/Z33I
twVHMj54cu8oAVC6mad5ryPa1+KkS2kreVnFvPL+CHJFDOSNZRE5da0gPToxu+Pv53w9B7o+nBmc
k2dHnozHCsxlLNHlJKvYHRzDL6Ba/02SmZd6zirYE6Aq1ABJ0z4rHejw3oLiL4CXg1DhgZZaXvJz
DhSo0U9EOs3O7iFKND5qrKd6CTpo4Zh7QVofi7mShX7Mpr8PbiqrWUixmpWE9B7d8p7KkXMxv8RB
At7DaNwtYqlDW/7qcIWuY0nUXGLtcphTaRNDfxe5Z878E4vyUeXc4uE7VvhXj1Iy8cmMjNs6MFLk
pmad/t3O43GCDLnifSOy6bikqGTh3KT3hrgRoDkoUpwi843z1eVY9EFvm8m2/Ci3GxLhBbh3MUOj
GjMNuIZ2EuA6+e+0r7C3HWepz0iLWonccw5JFgnOF2uj5mVBBcn53y0wp4p/BcBsvN0XuNX5hugD
xN5HuJzuVrtEg1UvDgMRSJuse1XD5BYFSlV2RxD9UEouAYqntniPQb/cPRbK+ldRy1g2P3rvz+La
/r3rV/2RuVtKW0i0oTQ5gXZV5/GYSVMq2KsNuYwGW7lA9FLxdI8KyvqgRbxcbV6jepKggwKQC9Jj
gijexUFjR8Kj4Y5MXuO87FmhAsWES7KuEsn8VvLzXEu052oUPbSbO58Zq8rVA1qOnl/KUnU1M7W5
J2VUFFrUqucv+ofugXeJ1EJFJgM5z7Lm4i+tr6ujNcYHY1xbTXOFjGGZyg6I7GHfVlxQmeWGXO4C
Mcmvr7oL5bJkWDWPzxC/k/xZXVZoCUsumFRS43P8ibE4RQ0Y8krPgXRvJHF/zRbixDCnCl+i0VEo
TTV5vHqFW2+642qg9Ck1Ju41lFX84TcZ6JVAhHyuoiTzw3QwkyxBB+OXfeIH1fztWzGedGm/lcyM
MJu9gcTVnmnSbIqsd21KgX458Hb22kka3FrfOkNKO6VbSgumdVUVhG+SiM+VwtEhGWRPgnK4imMu
csS0aKm/BJYgkDzOGE6DYLcCxZllLy3X4DMMAjczBpr8rQNyK+wbWeZKB1w9eQ9mGt2Pxy3EKW8Z
kGEarTMmkd+4aFaCVYUkqd455WjHQ6VzvGLaUPMwDnA68SoYCejSrRgZA8KfF7/OWz+N2qoFFd08
g9wafTeDzDOG3d8BvA/CgG/vBitUUS13bNUtTjAS3qJOmzRyTlIaWBFoatJM/iDeC7kcBF0YX6CM
0YW0NFp1kBkUNN5bEUuekx/qsJENr/kyxGsVVNgo/bi+UF0xE3DrjXFhbglpxDGxQmVWFssQH8zX
XeSL7oiPdI5eKKk6D9rGJe7MyE5cgAFtAa7kQVzV81F/V6KxUxTVKcBoWWynEx5iU6BtJ1obMMO4
RsPMBw+zEEDGY8xw525LQe+/GrlgNvqhWz0LagwyBllRJxPH94tS4afKz9mlys8cnqrxdFt6t8ww
NPKOd0sU0vocqAZcq89qzd7q59XV+B3U8TBAz7tp1ncNgsPzOEPhxaFcFb8kotP0z0I6N8yCq+8e
9wAudZw5H5a7SEK8EYJpvSItUOcCWiAqGwx3Oi5zjLN3iP08a0pjWNcUjnBJ0JB9SKfaq7M5/gK4
EfLErPO8cyWxhgO78BA6Zry0ZjQsxJupRfBPNwMvFHERlLRxoUqcdVGkub/v/XqcJa1oW++XPRsq
piOtaUaPTUSoXspLE9/qnOjLp9pFXEE55fV7gS1vmQm5/cdPqQvr028eNQYJRe1DmvwC5W4Rxmh3
Ev6xeGtqn8ZbjuIIf11uCLFgMY3Ad9QJDUFr4S2ABEKEa3E0DjQ5zHpRjQGGFLjkjGTIxEzu9UuI
yQtRsypyygZSid/Gf66wPcI2SFkLbzYuxObBd4Pruot2KdZg9v9LomFLS+5lvgUsBe7PJPN0W/zM
T6aUsG6O93B0R5vXp54H+gJN4uamAapVkqPV3zL8W+nskZmmJ6CkJJPQtzwCZHZPiOOZMl/kLYZ+
o2WvRyQodkk0SeS1QhhxAvPz5aSv9lgcxp7FLcxsZYFKuS8dlTBxw0Phh/FjFia1HT4ZvJXUUgm2
7jfC6RE/oYYSVSEIAG7voJ8y1BMZONV7gTFlWkZmHui3T4bFD2AT+wtAEaJTzqtvypGocwvAcWWq
j21piv6bkU3C8qBk9aFhIHWAe4cm/QDCEYJWzwb9HAELoVdXW7BatzF4TjyKgD/0J91m+uP5v8Ar
DAsVKZitGiYxVVfR15+7YZvquXM8x+2j+Ei1SuDWTOnpEv+FG6Go+Un7XID1SEw9wEHjAYNca1vS
Ld5jX3Zc1/Ug6olJuI430roeyHp/WJvZK87EkxZOa/ZzRfqiYpz100wUKKWNXbGASk7HWc9SQaCr
3fyLbiLcnn7OTmzCcLrXfrYubThtEmV64vnu+pKYWGB1XcNRyEXih4wWhPL6xN+oif14ahLfM4xv
ZaOGRUM9PH/fZ1RUv7pQjF7wzGaC1ZiX/SZm+I2Ul+skHLjfH+qaj3hyjUHq/5bf4fgdhtmNVLHd
oPOqlN1aeAvlZgwE0fOvu+0EOXPOEiPTAu35+sTNOwoyyYBYps4hiYA1zswKOc/sXCiEjRJch+6h
VdEYmK/A98UvjZwVsz9AycQBcJaHHlhQM8Ex2f6/dAfeksuWb+F+1X3n8ixYzKxcXcWY3uOfyYbz
G/FbcaK3IL1b3Y4Q/XlOEJDYe/Z7F/IkjASTn5bzInGVtGJlXEFtp0oYg5rVbdSBWBiRga1sNTSI
TL96/6qUdvyCnU+wl2bnxlZwXiYhIEtTTMPkbh0TZ7R+sfwgVDZsJZrH36HfLWSMo7Kh620/rJI4
wz9b0qsKKxbQORoykKF5SSg2F+dmC9V1JPDvECUgVcCdOmkkbLciJZL50+f8ZuD5EB46ZxQEFb5Z
YUn+lT+SiTKKzV7O0vWEVrQuUy2QUwp7IJ+27vunGhTUOWtLifIrXgFiwNxz0X6FRj4vZajw3FMw
Tn/ydZ3MN9M+HJN9tL7/dFVVwOxMb01NaUuJZE+Mr5oNW0IFK1NynQvTslGJJvELZ5oa8THMuBQq
j+QwCtDBdnQ34CGxtWZ2UcuXYBtPSUaKlc73CrQEgsgYPUqgHtM7tkbGiPKYuM0nd29F4QhyC1+N
CaL825Av4UUuBf5hXlWAz1qxRh4T/UsUR4IuwTBLVmQiU5qXJlKcT+snjyIsxsaQiEzuUDE1rwlR
LwFEFUVX4FPw5hdyDs+AVa+VhRS2I0junqx6nw9iHiC+1L7gACherK+2OE2yLZ5nuQXeWaZeknnt
t4qjp5YnV5FMR7I+3+vnxKO00C/Y5YHy8W9Nis7YXEP6geFhN3q8bxot8NmLZ8sSSlzr50EHQ+lf
13VfRlzwg+OvduhkOqQxsmWVFin7OnNtYBHcYsCLRmms1olYo+BYdD5ij+TAfEJeT69fOTkR7hx0
dDfkgaazBEcJQE4Zh+wXLx4IbjerQcFlKwjrXwON0lvzCmiJ41sBXS8Mkq2/WmD9Hc5ZRezJm6ft
FDvdGLKqhN8LANF2petiGjIDXsZ6yAFIQ+y2oQWGPP8hxogLKV2I3yNBGhhppLKdD11eYC2JArQG
Yd8qgnV2r8Ph0W+A6N1mEmVk/TTUQOovjMAieObey5fe9Gv9j22U5/xveqbHCx80cdcvZfaZMyyz
r7ydGRL2/ZpOPw1kz5WLAra/iARgOSsHlWzovVvgT8eFJ9Q8fxnWdivZk20VYfKyGNqjuWd1Amfl
KJnbTnMUMHYjOKOmCrgmJ9JFiSVTAw+3fDd4jznKVQ2uidDfcyqu9jYYPReo7rrA1H4FAhKcdhYO
oj7afpOOE2WVu/3tB5jKUV+L36PsmhuuiJDGlA3IGG1gqRhdas4nJHzmRfXrkzCcPzJejvl4OYar
YVpxbTBrVS9LeWY74UVN2EQHPsXz8/V4cuqmJsiPWGPIZWGNA+eQIlrR9r0JCgBEVehD4vulkWA7
T+dkgKPyFNUANlJL1iVAu23QqGiVDpRUXS0YLhMyHFfRLlr18YkQYWeuTrF41l7UcKgau3seDzVn
zuk4+jsh77IkaVHjiwlTdDCSRjXHDjf/dQ/JwV2uHxQEkRLftrsLlAYeADQhZrV4AexglVhb1TCv
BcNG8m/vRxlBQBq7JYVAoMMUcASEjRfMyyZw6wms2Y2ua+WmYaWYmVdVbMoe5MQ4kiezCr9WfMop
TMlggFlPJrYdksNNnicD3oYobiy/MfVsuyPbmxvxXj25oucJcbHvl6UPncGhavcxq8uYD/UBUQoY
GRRQq786eDHtOS70v7leu1NSAGofd4WxGe9nGPXVLffeuU0zqdUEaMP++BVwu6M0e6Dv9BNGUVCt
uy3sLuHi53H+Ip/H401JTMsY7SkPX6VFIwUoOo93Na38CaC52IwDCnepe6EDOx2c14hHt9RHJXh8
TUxbrFzI3dfZkmf8eJRzC1ieL8ctXLU+h89FN0h9K7ogpzxVh7Rk/JS0jPkdmkyoKCv+Lb1webmw
a//8llkz3ltbWonAegDKfFOOnymFEyr/uQ2hln4B/qNh9/69wCBniiQoJPSSa8MYXfRd4rwOeo77
Ki74mM1F5sPwR6Di3S9n0pU2kEdEnVwoW1GnCQDj6nUHFR216CbYMAwqE7irqA+6/vpWjv4LXvVt
u+rD0yrLinq/IdvQY4V4L+Xtdrmb53/8z5seGqbHXvT+HcJlK15UxDLXoFE0wz97m0UzW0IDw2Dt
KpzsXDA4EcSb18HWiQeEaHmSmhV9ygjN6s/JxmTWP8VsEr9j55yZgD4arARXeNarcPWtj/Ka0ei2
xBXqi6DpAsTt4QXpwbYtgPUUvDxwafP2hq2HWkDEW3UUoQQxFzirtQJBMXs2bsZpT5Jt12mZY7Ki
fEM44hrQpcLE1BrUj5ZkHZZ05GplO5SR0mA/1LtZ2XWa+50g3ddhQb2ftpWaTDcxzGX7GZa1ixMN
2n36XpT/Z43RQicKxrlaEfWOnBAVzFHOlJhugpvDYG1Rh4aJIefqUt8kAY/r4gKi2XXBP7ySNb9V
bbp95l+CsD92E4vpUZsSldD9ri+rui4FLhkzCy9IAlPAVYGe5mcaTH05znY+Qa/ETq4A9w9cyhQ5
EU/PMuOjE+TcVnT3S/90fdxbKE+4tfhmG8iu0saen8iOPyZAKPgcS+esSU1LN9ex6IbLvJD4gU7m
V09IZbIcAu556Racl4HAdqOcKflcaxntqudQnnXy+K02ym5RpJ+eUkA6Ut7cWJNm4asonsn+2Sv7
y/KbzkGMigG9gOpApLhA3c9Ugx0FZSmZGe8hy9LSiOMZVscsulG5lfl4GniTPFEU8biBJetRNOgB
KOoPSCOA0vCsSqll29tLc0RgHYo3MN+3jnivRhTZ0+bJU4vzELhpzLfYf3J8JwTSBpFwSlbxDYOn
i8e+SkXeqe2U5ugefMWS/xEN9hXf88HBDnJ5jOXYoIZaphG6J+umwKFhm6lsTE6IR10WiM0D37XY
k+aMgne5/AFVtAAx4XWyJtsLqffFvWv0atV5tpyzqEnuFkAgIW54EmvAC5dYiJS8ThexjvQPwwL1
7BNQVAHkORuMJxFRF+sVfgtOy+30Bt3b1IXC1CBT3gw6qzMDWiEpdMkl8SP8U9qyCQPVLZARYfJg
5WzC5jPdOF1awOj3jiJGbB55y1pZGJmzuuaqXml9kdQZv9wg+moFcC4J4Uk2wUgqEd02uMXQLqxX
i7/Hhu1zDpKOLH2BPHINv0qfI2+v6eNrtdT9sAtAP89EOjkfPFlvBhh23lD4jrHHEYmUkzp0ccq3
ZGk2dKluckc0rRIS4QhJhSZKWmgpl1sFWJCnlNT/9+lSKAYnmWanKmuIm0M5fiWUMsYCSTuyLq3G
6ucIibp82dSllHFMUcsEsVDwjSIqW56Yvqc5ulci0eLW16T5mPRoUgNYa0n0c7n49MBfzo/fzBNM
Kfnyv3oN3dLtebDLa/OJne/ApFR1r/ppUIFVFFwCyJlTUNW89s4LcTvgDZXKvkSxWQm4cgmkwwYN
HMTOQXoHCznQJDXEdVKuTuYpX1ZxyUt/dfzcoo6lHGNINjQ/xyQAHBEZM+DBS3zqmT9Tsogw45sy
omf3w1gkNmxMnW4NAx+rK6Khf6K+kanIhGlLb7du2z6vOsAK4yRGpqdErbsMObe5Xl2L3/HtHTm9
8doTkFX8Il3pQPgd2hwxA2BuHfDch0DizlNW7qSadbrWS5UCiVYQ5SbtE2kOg5T1vw+zwJUL/i+r
vajIO44PMOq2c4fAjUQJ0R3EFrgaJ1qSHZwPuXNrVudG02NHoJQN3UQqOXaHIvejw7X1el63BsC1
RzXu3F5wqrCVoPcIXRkRNd+orKxd0czo+y/6i1i5HdMjU9y+32JMfD2PfgJBsbdOCqYCzwN0L5N0
16mfBNlzAn5LOEbtMAWnhjZm2RF6dDDzUpQ6i7uwz2ycksIWCobFlRp+KeGOj4AtFO3gFeHsvrbe
iAHkMX0IdMqpakGf+Cp4p2VZQs+J9R2nKZz/0FIuP0jVB4nYzZa+2wMCGjpo23tmXfUkrG78px0C
Ashb8+fA8OUxZHZeoi9V6Ak/OSesRuJhD/7CqTIfm0EmjfyoOXU9II6NEZCQoULpxYNE5rKh238h
vE6HahmO7Oiorm7ASfEPflpqAeS6aUWxrQEPfR+10qeNTS2VSU6rrrozFJAIbJiMem+Zmj5DXx8S
NEPjINB7o1X6C7S0zjUucIiX0kv1gIM9+dwnDRFhsMkKrOJEEXDVT1oQKg6vrir1aI0kErl8HGqv
0zgevmc0O8qgp6BnOsF4tcdtfNzWMfk9I+G/Rg/r8egA3Q3/OzEaQvZGFtWR56cHatzORj+XJQ3u
j47m+kKOWsNtkOsh78sB/J6je0/TDuFc7xLXI4GWAQhDa0V/gQVUP4FPvgwJCAsEt6R8ca02Vkgy
fCNuWE4EPwv+ZpVMCDDB8C6gJAhxu+2tR2yTIQr6nfOxXAI4GvU735LuaeEo6syjPha1GRc2ahVH
MDbRjlNmNbmohVluk3piep4Y24edhdB7tv4qgA81eCEVA0tU1A5GSzScQKsMwwktOVzUHgMiOQyy
U7JFrCmNjiKMx4LKAbvycl2RZsgj4c8EE9VEAWzI4vSQrp5+kJ2wpmbExxsElvIbPi9zTnu4hQAU
OqS+ZrnNJW65Qb/AJ/0XLE47192QLyQET2t7yZ39AHVmCzxAXMRF9j3W+E0ZcbunKO+HxQZuxd6S
Q+ihBlbb/kHEvvxk+iQ90eR2uDlNJ2TpHp0gXrg7DptN6VwwMjjdxhuAHRZcxMb9SaTkyDqRDW5s
VVHrmOvLBFabHZDqPrGT08KKI4+rzV6hn2O2LPRn+c5EiRSNdsQ99FX26B+v+8Hftuqusqkny2/T
Fm7R3h/yFEKjz0++m6d5i1PxfiHbnrhIP23x6fX1vlpWuEgx2/EJwF5O71HO769wXKTsoxSf6pcX
1QOXV3wthmVyIKJlctWg/n13bE04FgzXxanX4KmXaOjnKdy/uo+vCeQ/QBqqzYAPNDoPA+04PyEL
7tvIWUa40mNgmVo89JFxAWQyPRxQEVHtCJjSNLAwrTuvyM8ipu7agCdoNxRHy59FpGXudwz+GfL2
wwOrE/322ChNZTknrPUrFaH7nDPFDWgKjkIxBE7cLR8QG2VnG+Ax1PB6KeVUWe6BurXPLTT3lBYr
iEwcIh668MBvcJF8k9jjLX6YmUMgIDB5wsOr1Ed1f2cbNDZG8uzPbMGEOPlxoSV8yO3Ba/iZeGaG
TmCS3jUfkTkX4s2YjPuICkAjeIncd9aEoMn+GnII3Fabx/Cuip2WqmJCT7LRmob9JxX4YaEl6A8m
cVTY3ELlgr7ilwWknuzPX5LHtaVOax53O48BJ2GfHjbKqImNZ2CI0Xrqezim6awKphNVffrBBWw3
hT+dWiQ349OijqRuJ3rjTHR78rK1LtjYBhcdqgrRBycS5wp/TLmVTVVWGPta0U18HN7w4PRF7PDc
uGFkenxxzPoUF+iVv+24wCmfGUHXXPuP5eY3nL/aRi8Fns4kiEFm5vBZSsPlia5xTHD4k3BHfeRP
OyrabN/5kLsMLomtw02OSJRm8mSCFgYSbh9Mzoxn8JHg/20p4Ia5bYfmmpjjFs+JpomD5333PfIl
d2OsqLR6Llxv13NvG28kZoiUcO2YZy53K6nRggsHJM92MwklL7xFrWz1UpnDRbGFrRDUjOHpymlN
ceZtSXDSvp18Tx/91S5lDpv62Q/KLujx3Ga8BQAPcoQlwFUzeDSQ8QrS4eiHGG5doFfutpCKMN4s
0yqLfxMHfoAOi2lsJJ88khqIXdQt/+reiy8eM5DCQzaq3NO/nJr6jKRIn1reowp5SHq3VD6viubw
cYvo+QIV2HzywLZG8kH7581zrRg80QngODTcRZ0rUsR8cfSioxyTjdGSeB9z2HXyXvNtFNOEtNyS
abR+sLmS1WPPh74cOrKfjuyDv0h9+1n0S+ePQQiMXWlcPyzmzYZ72Rn5MSi6T50D8w4/ZiBMUTo3
PxL4Dvj2ghCVqEc8hmZz24sW7dOrm2lE/qE/oinX2v6We9UeToRaEoZO6MiVPr84itQDJo+85Ugm
SBcnrCE7jRUI+UnX38uO3lQvtDBQNw0v+lO1a61emxbwrlxN2f2UiAI+erpb9MU1FPJrlHSKHUzj
2S3JsOzOLBVcByJoRjT6hPJICd+3JdLDorT4a4oJeSlCL7j2s8z0EUQIuBCBBC/fwOgU8Wo/+EE8
JdRF/AMVhIbqyHQdpk1lvPk8bu7sdRbqzhJV+85+KL91BcYyHz3WOwT3MvhQsvhHeOn0niR/oJBx
zGuODtLfVZelPfZM7w6zHtJ1hOainjKyfuG1PRPlf/wDRYzwkh/n/+j5qobaAHkkq//97fHTm47N
NhQzyk/OtXItZDZbA0OYGNvPM8A1zUqF+hPO2C+fR3Et+GENKyYT7I+hQHzNxi8ARqZuvnh5G4Un
zKJarNILI8mEGO6aG6rUc9lWlBnHZZuRonpNgzZyOozqAj1/2UZWUSdke/z1XFfUjKpQxVcoqEEE
840Q5uUldf0ZSEDPVhefUk6RHW2qpSqZeRHrBQsta8XRSNac4XNsf5GdRMy0ZkAiUqGywK2eVpOl
IlzzKNFXC/1SipzGdL0vnAfa19PUjiCCYv5E0uUcB6y2wUpiqvu4vaGaO2FqJhlZULe7eVIFsXeR
1rmNs8pv/Bgy/cC/9B+YrmFng4XTfFnQyX7YBQ1KClKPbvqlh8DLBAMKnNMixo0+tsiiVbous7Ek
EoXDNKH7ZjwkyiIpFMdrUB19eOrQgVTZF8f2WifuNir57U0wInhT/Ye5E2tBp+oyPyG5u+1Ql1ce
hWfFt4DaXyP7xTGsnfk5j05Yd4NNFy4irMj4ZNqHe5cv1XFa9ZZbPvomt+B+TXjsqEM9wi0OwDUH
zB9Y5PbkVNJYzlS6qlE59NNpZEu3lGrox3+wkFFuk8WhnQnktZqoC91Yyx5EKN12jsZGEwjc6I0o
TeKzIy2Mo6TCXH6RPWYqiygH439v9qQyRSphV8GugStMcAx4YWIy77TPwLrHBwgpvS9JNeGJ343D
xZtwLoMY9rxWQqcmgL0PK2GA5LmCgDphCpt3J6jp3xG85SEKa/MSZjxolmPcQCQrGq7kzgv6xdE7
d1u3FGHLkXULWnVMiFEyQSKS97aE7FPp6rIq6TGD2hYj0q8WsKGFNuvu18c0xJ2bVHMHwZ17nOyl
NZndMo2PHSp0f3gXYExwOyaF4Am1EW9eTN+Sbtc4vB/zxVdsywXNRpcTYm8EwVx7TbpB2+k35fpq
xWY5kFgjlWTBNfVByV3lJ0EBXUOSJAxT46NOPSxMjaMyYo+S2qOKwWxFiHuJtYyv+uGrzgFd7NFO
xJ12sND/kB6msn8NefA8rSrMCfGbwG4Ut9jngGVzhm30r1maW/Pyfk4Qrty/IR2roOw4N67O/byL
C9CdN7VU5o3VPdb3UipXqTfMLaT+QRI3h/QEJ8HvoTuuirScjP5iU1DuJ+4wW5XvsuNZp+812URR
M9PieWmtRju8JRFHpPoYNesoaluwd5+6DQ+E6itamwWSTefo0QrGtZQEZcZaV6XzXx5mH1MuUnpU
nKks0NyyzKyMIYHJnsmi/b4WOvj1QO8vErXblp821ZdEF3ZSbQu3wYEY4SPKugklQgRsdwI8je5H
HK3Ll3hhbln5vswyTrbem5BO1u6qE2f38ZAWPTRTsv6BA6ucmZ/H6UTsBpt3pnGWTriygWxtZGo+
XsU1BVaVK5SvSZbLm0UY+tTWB3vc5C+e54ETbgArqvu7fmZ6hNU23XE9tzTPSpWeXh4qv5ikCgo+
yWailVA+JsRtTyh/NsacnpAUM8l7ve83j7dRMmJwdW7I82AskZG6wm0CycF5zGbZ2SerMRCu/nW2
t3WKpoBNCVT2FIYNLv6MzBJ1k1VB98caGR0R6EoXd3CxpvQhFjwJHZXedpVoPPnaoMkyNnW3i2LP
N/szFKO+c5+wBFuzQ1oRm7ynU3Pme0Pcf6UuQ25xtrl41HT7blAeB8UY9YS1AW5Vw760o5Cgf6CY
c5/gMi7muvRssJGtoBO6ylNsJtDbGUh09hlQPypQz2IzT7A1TJECzSsRFU3DtMpbwrAZs8DQ29vx
MdakOK8Efm1pgJUkLpdre7mED6h6UadtmbNddilK72WR3EutUMFk+TxWDHznbyoEULcqsrpHTRtQ
8/qef6jocdn3MIaJtJHBS54eLqOaeOfYL3O7g+H7emCZozmYAT03w4fFSUeSSwWxlbz8HXHlj5yP
9+6bDFaZ0y3iffoPDOvolTXAIohBFXlTaZYkpWwzu/b97YB+yOE3d9bvPiVQPvBExpKV1646F+fr
crSLfEkBHD6qs9QLsUttJl+lMWcpwZme684JBHcuwYkK+D3myDqCEUcOm4oN/GWS875fMba9EwCT
lLgI0mJ9TCWyJah/Bgp7TsRiCG8FLjBMY6LE18PjjeVxKEsHtoNKuNnik/Bamzy7G6o9a/4QRHw0
svDrBcQvCgkOjhWXX4ZjAqxSxSlPnhoGzk+Kt4rv+l8bnuQSx1qGet3BcNuwTRxsLZ719lMnnLON
tmoQ7ADyNNZwn8Y5I/YvkMywAQnkCJNwQgtwGqI5kjJMLDxiu5LHuvrrI4W+hMTR3Zq2jArmM37Y
oo717TKaGr2dxhrCvWAjoe0QMRm6hMqqp089eyTno9/Yc2zqndeP9VAAN5YbFP18DVcQ0ogFKB2s
ciQB9qbinvdndnaHe9W+GfJHUgXa3fYXtNqBtI8N63i+oMm8mYG5CMZuRqDQJxDz5emJAOvG6NYK
H8prm3Nhe507wc7Wxf39wJE3GpnCB3I3JARq3moAS5d9Qot3hB5WqFvIBJKP3A+B8rydcc1bV69q
inA2wV7E0RsvpBGUSYLTjnw3ud0d4UZAUztKVhhWvZ0OfN3UXFedbDL6HpeSAJ/LxE/XKD2hM9d8
oCuN3+pG+GE2EYZspvoCpOBPF25OHISkWPHuM8L+gwTxx8pRYv69PPdgCz9+4dcAZpurgg0b4qiW
zaTJpZkMueUZ6MfrzdrQzeaAyqYNQxdvWWCuLcCRN6+IM+6OY91ZOdAZkvspRK/a118nnuYNqLgM
0ozyuJH3TWe43WrniZ2+MT6dhjXP0VF9Wb+yGscZQJPsymQn6FpTYbaJvFQ1yEF63XOgH02FRYE8
R+KbVsfFerLPwVfZDOgOIR+7VhbeOv6XE7d+sjBW/lJEo9ddcqmTBF4CPzGIJu8BklL3dzEV1vCc
zSk1ovijXAjNaVxOV4TtpJ2o1O7yckdp4zBxTFMPoXsAppFXTlgETmyhu5YkmQxuu0DI8zDHoeLU
7EDjXB4iEdvy7e8qbMadVDYJZh84XZo54m+j6B8wQ91cRTMm/AFGxCy+42tQFKj6+LKV83G4Uuag
zPu//cHu5UjgTD6IyhLUD75Ni/QTotiP9NNPQ4ScTwppk0dfXIVFPj4GSuPBPVACU0Enu9eiyafA
R4tM2YwOeKMc9RgR0NXNuGC5wqilEzFOqo1VuyRMZa4h0v8/KfRta4gY+m088awlIXN2t0OjQtLj
+Jmix0GoXtYsnlHz6st8vgawNKbLanf9I8jC/2vIFzLigDhv5ctm1WzXZpdU8qy1UITNSLxz4142
PP/rxuBPADItCxyxNpj9gw3I4mXgqfFGilRBILIrXOcbr/enIiFJ6Q0/IbfKTEHJBTnQTTK1duvo
5v69diaF16Os3zHHvejMQqcXP3vRtPlAN/0JmiQNJIl2Z2zDxLEIBByD0MVIVQSrMhkH/49ow1yP
ax1pP2Ums/4KKldNVGF6su0QGeJGScD+qJY3cOH6GlW1iJa/CnSQ/p8Ic47/uauMo2EXkD5zW+Ut
z9Mqe0rVGzcP+w61EVg5q0mrklWg6RM7aFnws8fRrBGnM6PRD9WnbUIo8j8z35+m5jltjRvvgHbt
OgeC3DTcSVFekqcyWB/PsG0uIwXk9R1wUaK5WAOihiYJCROBqXMFudj8D5A2I4rtlYcITGrZHKE5
OCHv5z4YSckYnLBwY1W+h7Put45Ma7qHxmft059Fqc0IJg0xMJOR5eslzcWg0nePe7xZ2kt6Gzo9
J4GGlTqhNWUOW41RiL5/nHD0ud4LhfFVyolrjvIpIC0zscyrt1YCmdOFznpU1LanmC+uicyJn0ER
enkws8Be1855mWvwVg+4S1ZcVL36/5wkhH5ImG0Zf9+q83TLsloaXNkPQeT0hqYMvoa+YGefWzM1
bP4d+nHibV90Do0cT6Y5pglfVm5sFAMw3tVLSSN+DZKFqRGSxZ/1HXbA2bCvptiTI0pS1/ET7bp+
tOH8Dx+ONkBt18AU8CzC96wMi4Yq+dnEHM5p3BdB84wRaP9UiDDCcW/VLs3djkXkNCGubdhKUVbf
KC5D2v+qPZ6ME+e9BBtS2wuwXm07cw8cHkbn37PBCQnu5GD81WUpIAhbzQbK7cTqHFoehFbwRaGV
ercEZANeKb2dNAH1BaJdAbpMCooXq5hea608/ROxs99CNuWCeZJbXhsl9MTVBrmMTPTWm5GP34dx
cYwtmYVkc497RVLQ06Cirq8ML4vE5u2nbmjHEz8yN/7f0TjlI2EKzhFvczkoorYuk+SbUqIWKz6c
BfaAl3ltO8hVqsVQAgaAVv0UuZwHbMsUWuvuEVSo69upjeqpwWEwnsnYqQES6fR9BADJpuJ8sZtK
PyFGoFrFRWAW/19/zOAacpfbJHXIOmKCBLptTUlePdrTpUth8DtsMaA+IWIHOYypV/ak9gVl21CX
wHRgL98G5tHOZyTetqb5J7mttnqdsS3w10YtLWkhhIJHgGdr7/8q40OdUibEyuxsgdlKCkOk7x+S
2mix/l2lcU2mjYqrqW3JOzsaQHK3M/r0btiGaE9qXZtqXJ6CeBb+vEiT+1quzOZOgAgyHJ3rvfXt
kyea9NdRo38PPfXsyhaFGxFZxzP1wBLECKWwyEhJo3KrQjnCndexDTGvj/8i6L0jO8chC2/ajQ9v
qqTanF6vPOVe2UJV7lXWA2UFloLECgPAavKqHMa9fVqZOxxPiL33H9Fz00ZiaDgk9r1bYc2HlDy1
fCkYYH0hOVoWr0kNER37uKKQZ70VvneJ9waM4UDAxAa109AHJeHXST3BVojIekWHMLsNZmvF6mT6
PvNJdVQfdifIAo5HFikVjJghQcTwqXXo4oOkGACHW+vekOedDK2WDyiMHF7IZE0Im9nCiAdzZ8SP
lMvybxNeoL69MohhqPCsJ0MVZrG9pkUxcIiZmPRM1EzSB9U6pVeYh6zX4ikHcl62VF0Lt/hcLmDJ
cV1i08nJwoxn0X5AbMxRa+UbnypnhaUev5mUKA8vN4nkLi1KDfaAsRo/dVX6/VMCCN15k7WcnkCl
++vRP44ELne5VAjZj9yqKUBj3qbDX89+bSVaD6UNtZi0J5QtaYXYgW4W0rywEgJpN2TNCYX3EfAG
fs6AA8/ao4IHqvhuvAakKYuz890n8bWILoEZJNYptENDs8fqT3PCsFFsUhdXJOlFfwZ6qcj+yoUL
Zkmgc+kcBsrFPl2+alhsPwMC7K6P4LNh/EsTuo4uVYYqS/Y+9AVxX0W71bk7mkAj8HIJ6pUAou1g
hgRgoweveMAVoyXxW2ZTbSu5vszQN4sZD78xz0gWSYoMhTxqoALn3csHGpfDhnYKDPDGBdk/eVjW
ou7Q1ycUsS0v5RPB6goMh0AzSnaeTWafU/cY2odtvLiZafrZE8UdvCJorE38Q1BVR+HkR5Q+9a7c
foTJIEh7YEHFS95c2P4OEowhH8Th2xkwtUEBT5whk8eS8CTTBv6KkzueLo8veoOtG9nx0EtGd0eh
ijla3QCdtIjCXt+NKHjYqpRZ4MKyrfhqgi4NPpiE4oOOEger9b2NqrBTyLWOGAWlReq4oqS5swjc
aGuPe/tbwUteB2YGeQ0ZYnKcP6lwoRZMyartL0IaDFNmfEjE3Lrg+gSF9suRU5zJnapnCB/qKT3P
Mov3IzL9NfZp6Dvslhekpa0OyBd+sWyuN4V+aVZFixEO+YORvfBYl8WjsY4v0mPZ9sTyjm3GBYNl
0s9XlIpMWo3U9LZKAtLJYmj+Nt6TcpQbmSJtankQ/bEHavgzIjQkF2yKpKQSIPtC5qnXMGybZ09O
7PgYyh4AcWNnIKiozduN23p+15jvVxTGKZ48HVtKEelMPIeo2PMQ8oxujYyCwgKBW67Ww6zfrc3d
Vtd1tjOIv2AFA1s+IKKCHiFCMXDMOyaehOjAVUQdpOFj72YGn1XxMmBHJBzXfhJTKynjjSqaUKF5
N2sIo2K39CIfs/VpkZFIqBFlI4JUk4Ccs3OAAzxMWeCYgxlwYN2Y9rKBer1r9KFWiWEExrD5Nh+k
Cx7ulkvPq2GjWIRrrJa3sPsrghW3Ywz8puZcagRxtCDFuh9NJ1QuMJXD+2EmU6eP/FCr+vfJUOj5
rwSkk/RO3Lh+w65PMPvTickmysGIndHhHeox/bawXQc667Q5nFyeqtDfsJ/R+IsfPEIKRFjP9zpc
IDMSfoIG77zGSmiRkYEGUhWj8R0IeeBt0hOpWBct9/8PrBEUucLEpAR4UCBsZfN304tV/+oU9lrb
csPCfIyTzhGJsvdtYmA7hA5qEsZULLiq1RSrjfLSDB5L3MS4BnQU9b0ehbduqfUdQgdKDlLhj+EY
zz2cRPt2PgDvv3EcPPRuivzMlfYwmZU5F5ttWGhPPSwhbp+4BcRNXcE8QXWN/VKvRSZ8K33vLLFb
N4HNSjxOwHN0yRPiG3/8JUOkpKY06vIssi5UzrFi/dATSH3WzrU7zE+ZjFP92u2NWPXQOQWH0HYt
AnO3jPbUE1axzrxDqFJQ32C3YjOeq8shRQevTLwuADfvYcrCH8YMs6XpQRxbIet/NRAk0aXdRQih
H/vivJdxmfeHLCSq0cBiy3dIIF/rqfK26ydllI1mN1vqA4R4DwEybsrij0Qd7Vhn51Ntv/TZxD0x
lwV9QlmbWJ8jvneSo0lWfoFCqwQiVpxFBICOAPtk88X3UbrubMx5JK/jVhuMQ0B+cHJUe4uIcYkc
LwYS8OM1lc2oG6SiD5AYvJqCAGDsrLAoAoAzZlT++NHdX898SV4fnz2NYRaVO+BR6KEYVGpxGWVp
fHh6xiC+nCp5aqqvE9/D43+zInJJhxlTN6AhegVIbJlSma/fLU3SqnLsoAhAiuC2XXdW0Mg5LQWU
NqVmUdi+fcXQnqdLqib3lIrMXolLL+YRv+YToXIv0MZp7zhNHTmfMgoIwhXuiLiwNVswpO4bMxxf
42dDNPPbzrwqb3BdgAunwEdyCV1i0m3MI+l8jI0EGJk2YnKT1xGQ1Z4NY1dSeNUOnV2hk1IDUQyF
QPBBnIE9QE33PaareJfL+vQeN1HQEVLxGrH4srbhK42qII6N1cSm6F8w6fp5MGaKWgql4sDhgPJu
1rL0YsZKOe9Scvr5R59e8i8m+KJOh6GgUyYSKJ0s/OkKAy18bnGI1WozqajavzXTLUJhiPLXcQiy
j4mMKGQVAK/DeV2FvZIXLPcFhTASa6Z3j8Bl4O3RId+987DMRi8NpahJp+MRI88e9ycdMbVRD7hR
kQfYceaSTxWnCv9gvsLsevLXN5lHhezpcbInMOAGT3bTUaoyHgbUL2LcVTHyiD77KCP6kBkaL3nf
B6e4PPZoMJCZQC6bR6J5TyboXDnb5hALvJC2wuMfj1NTsgVQUoY7mY0IaKzm4vEEAo4IWGXUiMUl
NzZbaz69ahgX2GRmw/FuZC26ZWQEtyc/4kAe7A9q1EgiITZKAc/wy/n+l3l9zL25lFbFO2CYdaxN
HbfmOWUpq4OZ+l2SLlASZtd0bTrvhFkK5/BGvhc4gm3gAQzMG2FIHaAqyTZhwgFSYlZFRV9qVSDb
LzD5+Aa3dxQe9gChhmcBU8jX+zsR4ke5AEi25ODm4P9CA4EuDwAZUdYfb3pd2Zyyi8IzfkfyNFYa
1scsy72kS1RM4jSjcbSBYUHV0GyQXAP+yaxzqBDAH/d8NizS6iKRaL75XjrSCMtitWRkfq7sm4P9
+s8Yy3apOO0ec8c31yKV5uDhcl9HYxGZRDhB8LDogUvVdcSputvgY051g+LUYpHNgy3PpR/2jzcV
WuE9l1/o7PG6w5r8Qt2teDg8JvbsnWqA8/vG8kxxo2S/bJ2OzvSlPB0D4lRgB+1wSh6X3XUlCkZi
o6oOoq2L5p7I2HUpxTBvHv2tQYik6WhSNLhispIE2AK6jH2e0cun65gjZHVHwNnihzX5pMfH/6LV
zWNAja/mox3PvJ+Ohx/v1COOqdNypfBzHlgBDpUt7Kaq9SGfkEHLqTqpJI5CS1pIKDWCxUBtP4x2
ZL3MFM/6KO2p5DFK4RZcq6UkqafA3KUYNrLeFDm9VzwEReqHDt6wSSVVQW7GmfYCwmwWuV1IawB2
9LfhUqKE3gNAuvZ4P5Be3awRU8HxwuOPHgGYquYhpWS0+b80kfxRa1RdZfxQDNqClhDm9wP3I4ut
BOW9gBvwRv/VDTuDt1vQNlS5w2mVB8yuF3Da5Np5AYminI+WbgGe+NABGf7ZsUOngO665RuKDjbf
ZShqqHjXHDYMpbtswBxDnxeIhxRswcb+ul+GcjvRVIWnZnR7UrDbkhlH1zG/h+yq3TO4L0R8wG6Y
a6Dx8iAAmUnduAq+wJec2JDhYKZcqdgImfh3Xz3RKnYFrBIz7tP+/ZrZmptiMpnwt/esufeTYdeu
P4/BJtWWQnC8RPAVKcdR5YYW9XCwJT5mK6yeYWVKCRuW9faF1SPjvXRnOLvTBcZ/zljMNNkTW/iM
++5mBjoC21O2qF1HL9/er0sAYNE1RQ5HMod9qythrG7+j6EAgfVcUzQHjL6xIZ+RXnf+r9zwI2ta
tfQaJEPO5jIYTOn9pTLU50Jy39yReHhstDUJQ07JHijfEiE7VkCvGRPszjQqwO+oMV1bT0eweVJX
4hHnWpWDYvPSwcTAMFsOPWQ3aGtkzmeANb5lOxMCUfTw/rulAnE9XhTgpmK6mTNCixrgUTJPriD8
nN6qoe5qcMJWiTGgtClwcue1xcuxzjGX2nr5HUHNMN6CyrSHYCmN026EImy5oncYTPCIpwoBSzM2
o7zKOORPufiwn+5SSEyf8eLPEXM4YbPYdLlKJKwvZMNEtwxpNmEj3B07RZx9F6MEa5Du99Xzoylr
0qeZNYL96RqZst1kBLLM28lUajc7o8/Nz8EDHJrcy1bxPNk5FFod3gwtLJMxijOxrzc+id44dii4
JbjYoWXWh5bepJqVi1n1UMZqAQJzggtDib+sFMuVU7FNwxR7HLzQT6FXIuppR8Prn0T5XOSH3WGa
n+qDoTAIn0xs1MBtCw16SDuqVdoOC5AqhNZWhdl8JifzgSbDB1RVTKhZ9L42k44S20XrhYrOVuC1
t+9ZWBy/IKDXH/H7u9yJ7GhQL9BNr+xUD1Wyf4pAckQblYK/zDZ/0gOsJo1+JFjvAIyHMRBdyF5C
j5iZN+1hR82/HQWD9V7U5tqV4yvRE74VYeQiusVTSXAcMHqtsJc9TwUdkdUBbvFDaPHd+Mhftzcc
PjRd6tLo/RZhD9bab4pfXtbCgd046YxN+O4QeOcBcx/9EapCdFz3Qy/pXjuG1Foj1NELwafpbck6
WPm/tVdv7Yd+nG7alU5SgFEAm+s2m3R1znTHIB/si/hTK3jZN9CYyNeSoz5nV6IaN/zpAxynCNuE
Q/LMo44QwidO2LNBCIIF8tJQoYR1tKGLSfCi7WohNeAj946rKCoVTD5PKfwrC+rrA7DIrpEB8R+V
HFinDHElP6ydDHpMJ+B04j23LzwYR9O72i6vtt0SqCrxTkwaIIs1jOO9aLoyE+kbCaE9A2rs/6nR
DrwE/usVRg0HRlz6bE6uC8ah8VqsM16iYi2JweFylrANvKZpGUJQ+woxc3ZWeGeEDJK539zIh+pI
gXOvo1B9k1t5FCO91BsCD5u6ZM0Kr9+8RQzs8kBtWur/pM3mwiuCj9aIrFRMp4sX2EEluSLzDqFq
GJipr5ydPJY4/QGePd5wzypzYLzEIzAr9zJySUEQheRKs4KLtWZKvKx3KWUcGIgxfYKGul5Fj4yk
20U+8sqSsy3FNlO81Ueoe+LlnMe/WnKSNVW7XbH0h9TvuTT/vzgbTkd8ILvNEDxTX5/n3PphAH5w
IeMTjK+9kITyf3sKE9iImgJF2nrLKRvZInJRvjxkh1pJnlNga5yiS4rW+SBkUI1v+0uypmymtFpa
4xcmdldrVIshEiHHaD4uJcgwFgrixJUvvRzw153qPftbz9pKdg5u4fscN6O3px3l5Ifxc83LNGva
0fe3PGA4twFFfrB88Taq7SJXF9dH0dc3aHQGtVNSD4qS3ncNNYym5rTw64p3QwEVM+E4oCD3BSKX
H46FrdoylO2l/aLbQ2xi3/xH/ASV45CzrmFIoAnoJQr7WrB0mvW+wcaigr88CUDcCQ/eUYdFHM/M
mZrWUGUL+qrEZXQscFUgRCHqG7giA5QqXjJa//kAP7RiQE/ILfKXMZRioSvvY//p0F7B0mayHitc
vXkNTE85s9oOKercoyxGD9excPRO+lBP3u7Kj98t5UrQti+zbp/kBAI/eLrwnMv8W2NRb6YH0XQd
+qqfQiEDaIjkRy5NGMUtjO53AaCOY52rPN8zMPyz1xeTTw3YV/1V/Mxb8f4t65qeOiJ8bSxtfbsb
hcQT8l6C6OHdbE6OtOd6mAG99diT7A2bA8lShtz1B9xCfY+STXL8JsJ/E1+eFbDtAPNsjHgLcFRG
K368XD3k2EPSXmt6nvCWlM63ggP6cTNJWwfDKF460SiuWGHE2xELzrqjzvyyviEupdwfoWNh/WnH
TeElDLB/mBND8H9h5YVLCtien3pdiK28bUVIRj8G3I8i1lAoW5k1W+0/3qjPzPwQNhs5SKmgGf4R
unLCPzDjYGLrLKtAJi2pXUzdX1KtMZ4FrZhQ/9kXpyenFhWkqmJDqG3qtPZZut90vA3UQtlA97bO
YKhFj6wGz05nSgX2yd+sYmCG3bu+umtFhOcdfOCVFuA/sMJf8MBJis9PiUKlSDVlEL0kJiihB3OP
KMr4RMfrFpBDCL2aRG1H1zq7WkHntobfnjMoNyb5CQFIodwptMdntAk3eZGFIKzU7sJJXWlTDSC0
ZK2PwCNqOPjNFuG7q+M3xLPuvcKcOWUG6xdG3oYVL7l1Hu7rmLBknyyvtnR7XYdzzT7Zprk9C6e/
FUOtPNiM4fKZIylEQd2pJfOzB8ieh2mLCUISLq6wZikJ+r/PIchWU36DQnHbhdUu3zl84cscyKp3
iUAmhzoo4gxScisrFLiciG9TA79WPB3gkpN5GpZwnTFD8d7xybRrjrHS7z7GlRVzlfCTX2UxnKy8
Pv5wbyHuAKnL+7hFPvdWFfLW5MKrlOV3uWMN/aA7SMFKAUPsOyn4D7LfZKwKonS7ngRXjsgyUxKg
WW/d4aYOqOhtq0PxO/3q8rXcOfaQfZmUUUZEPQCow9FGkINl2i4+IciFOpu3ZNa8qghd3kF1/aAF
016yZkdXUQayLuFkJBz9bLmTLMIyUuWkTxZX0IwPD1RQvrPe0AR6pC0jG0JA2D8AyHVP9Ttb+qVj
y5c+JeeQUQCKdCvvtqadFVJgTBGdgjoX16vB04+AkDSZlqQa2fKaLMFkHhuIW4Fb/w0m1jwgMf+C
+EN2/ldOMy/uFvFXW9ipJJEcOZwhdmHMnIJoNTtxlcQTtcJz2cwb6rHyW2/fNtk3R31qNQaImTxG
pH3DlPhQcC7RCwU9eWCiU1G3DZy2LU/ghdvqxgXQ7cVKVDX0uKOcSwWnzq8sVeR25q+JVN4+ygU1
eVTi/jDlgMmP5PLUKMSn72cCj74+HPZyzOf6uP1pNJgYU9e5aiEgC+1dXDWqD5QwpCWLCY9L6cx1
6/jTI8U4T7XRgBza6BHbL/K3+gITiXDiXqyncnN53WqKML67Q5DxHqXyBv8MlQtfuAAFljGHAatt
foz/GHTGC/dWl4COwnH9O2S2pX9QK792Gga5FJ1OMPnMUn+/tg/IFX3BjIVDxmN+azWl9mImJEp9
3fIrdHBBlPaorb7JMU04LAl0HrhWMjihL89g4uApPJFb+6+vJDF9cw20ojcxXl5LoRYcO1gLUCee
LW6vZUSJyntYWZdgJyrrLefwKjEBpXFusvvQ/agp/tGsAbbB7ABgKSYQa4aQMqehlto3G5bYZksN
vN4XvQTHzUi0noAd/Ip6FCV2giCsuqO7NwN7IwKJuSrU4ExpHl8Z9FJp6fL64wUXHuxhKT9I5Ekk
Ty2JtlyLJmtEtKvFV00p2taA8vO9OIBOpQCmX6GYGLY5RuAlP/3lg7m2BHUh0a8q+iuHP6DD7WAA
xs5zrJw2x+FvErqBaWInLoCzN8CnzJashxKyq0KPCONjp9MebCUSDrPATO6/h+pWPajFGhZRj/FI
YCUL5gBk1dgC2PGlPgewOGdhLs5E+GBGgYogliC1ZZb2QUi6/kz/AAu5hTr37VIE+lPIyCXCyPC5
na+yLDWzqu7s2wC4hYSfsIR0tls+9qV3g29bTkSHPdNubPLblWVEw64A3ir8DWG+PsIxKJUugHHS
Ao6xVYlzAAHtUuxPOyWctfVG5sOJo6IELPSkcBQsfqPlb3krpfBeY4PsJLdRmaeQzncut716cDdK
VoEXqqCbycY4X9iHtpoyIiCtYEVWPO77Bw0y8DmgBi2oEm/t4Lgap9aFJC+pL6DqYRbiw9FILmjh
kXGtkQVfb8+QBSf6NNLROap4r+9CFqOe41PcU4qIgHU7LbX61r46xtLR8EKNsbCOXrOCk2NoMufY
9Ti1x8viG8VTI52dLKDQWWPjKBOa8NTUeZ2m5wVORGWAugpZd1SxCIWbXZIOVXcKBZq2YzJKMVsb
vF0OgzEiTAR3RDvriQ0CY3YhAan8xVZiAZk3mzrIugvbvqAYmEveLJX5HbBQu24T4EkQrNcuEXZM
N8cv6zvG1LGCta4CWUpGDu7sg0hb+KDMSNIXLudHGA42Ld1SWPDSR1Nubwdy4QrStfB11xuZ3muo
MjeMT+IBevr9QDPpEy6AaOK9uMHM8GACX8EVVFP/TIrRV6Bjyz279iZAYXTwk9VAwqadlsDz/lq2
8cFWLn7Yb2IxMGsfEjDKs4G3rotjhK3eCngONbRSJrf+IwPSoKDSEJi9JAQg2g7gSocTW7lvuCF6
nNauOnh2zQouHiXKYqzUBtapPBr/0kHDzvZ2CKGQPUYD11o9QiCIqIhvUtKxiO8DBWDvdTzPkTvW
pcqAgEDpkTLhOtooBrRgN7B3lmlhZdXXxySyKTTSLI3dnqXe8/pLLQKHGCHt05fas7knLtb0AqtD
SSvGitDsVJfUcUTbR1yAzhZAfgo3EUdEKOBOEqHoiVhoUuTG3sv28o6+4EyQXRT8skwyM9sgebbq
5PkwbZe+oSgr4zg8Pe5r9HOdqhE2P8ngw+xXWpyTUmCkvxE1wp7wW+gnHGRnUtc4H4YA8Z3qUTiC
DwzklQcwdlYkgEYSg8npxeuq9nQioSLT4q8z7GA8vkmgjHkskCX26mEDxlHwfzohUXEVPQksIAMp
HErgqf010ZxV0myZfQfJAPyG4a5Nz7R1lMacu7ezomx1ZlY2rL8m4+0wv4x1jJKL+cLSTd5VKn72
KZ8WsRCKkk3F8BhCp78doasqQ5nCRpJ7NXbi2jKVbA1qkbRQNfdyWTkrhWN1PlpYj9mwHqTLBHqE
FkunQk1G+0JSVEWQHEe4OtecOrAwB1RyD12Hiadd+AYB5fgek15bHM7EvgO7z8/7K7OixuFhSSt+
zaQXk2ksJYfk0W1N3J/bOevD2BeSPpnaADiCKtX4B4uyfLfELGYJsNsPuKWScTIsBDInljRIoBfW
MWHwmcvHRF4lU/9xfhh11muJa+6YNRl1GDmUIlHEnGegATlUHxgsn8t6tC5bwu1Tl1rITLexhDdk
YBUNq7Jd8soa3rKl6rae4JkDDJpHdsxFV9r9sB6MuKWgRMyA511R+0n8MPk/ByjFlfShYjNJZYFG
HmcfTKEn9irJ6uWg0A8lPX/VBV26+hc2x+ig08sGYgkDOb2ISpnjd12xnvoXVCCYfviUOpH3E5H9
t39hU4YpldGgMda1lzKXkm0RsVOsrw6oDSZ7StQaNOEozduQaYBPgmh+PW4um55LEeILcV0xFJEN
I+/JQFmLZST7INhYj3cKMXL9O/AckuxxLYNmbMzur0w8a4SSudcXVBtGGR6Pg5NHUPMPvxWff1Cm
nn/1UhO4rsdM6zDQbss2kq90Ro8XGg58kiX5gqSqCEiLdq+rLs1pdj39lnhAtOTOGz/jBiaIK0+R
e5oLxbnVADA9kPsYOQqVhy38J0SUc0imNCQDw7NXuDE87F7920OsuJnUvUt1T758FVgHjiOj1ABr
vNwm5DvUwA+SzIJ+CUngXaoZiE9e8jCHILatqNCVggtSXgG2Tbv7r7U94jGJqPnr7ZiO6wroQTY8
nnD5SZ98EBcDtS5i0zyXJG9iY9K0Xg4DpLBuq4227IzYrLWuDvhzf7L7010zwPDJHoZsYg0mp7Gu
HfEMHbOERNAjrttq/6jGJkDUPIDT/lP2IRxYq9EGLob8a+gJ7MtuchQrKk4QkS33AA8D8ew66su7
6GLcfrNHNUMVpwI54P2sB1eyINETNlambnztUJhwBw8UL6jueAdLIpxlF+1qlDpaoV8gAyvl1zn+
Pn/exWoQuIIxM6sPwcUXDiLCKTzZAUe087w4wwGD2WWi8bM4/TbfmzJfCmJbyAS2Nh+G+ekrbCwc
6tljNT1SJy9jHU6HGOwVA9YqRbfITJSENfeGrHgsaikfvBVZssOgiLY6KbThBJBkC4SG/4iT2zE8
HvUxZJR5Her/K3Rlco2zG4Mg9ok10MyWoCDUQI1daa52cwoEqGW9PRqBAz5CSCmp5aJ0Cqe31luf
982X41+YrT2vlO7WkV3PhMl07nOpV68dhRC1iiyALnFFVFBHasQtG3vGqq/MSPXLuDc/zzX4DzOY
puY4eis7o8WUs0SArDkrHSVl2GNmiSQkI6CGlulNKgoBgFM8hG8O9slE/5KhlQqCnycfKAvbeVHr
yleXlWBZV0QnPKW/iqHN5lKcH0RKQH2fOFE/aCGgvMaKE5rgRRM1wp+MQ+frawsLFIXKUbYNjYQM
PjqrN4aQAeQZZSjzEYD+g0qrFcfnROxAHN/92JFHW7wD6egAUbDNhcaRTroe+yEjeyNnDU/PuAX5
lfgkwokOpLE0TGvQYy0Oypr++UIqNlnk839AvkHLj83Em+jyB5bpW4Cog7swubGkkvzqqqmx1eri
HXhr2EUUbkAhLIQyUTiSgLf0qcLk9k2Cfr8BlEw6JG2/GGoVKY2EqJomOzx3ZzTmekt2bytkMhic
M3bsNjfWsu9HXUae4gM1bxjnkOOpR9vg4517T5ivd6X6Wp65ExVaotqB3fIbONx/aBHfX+iQF3sm
gzBdEz9FseRNz0QmrYqq9RgtgpRx/1NjEf9udGIgbxzBD+4Cgrf3+R0N+cB0o3snSsNCwJKGa/Xw
+TEVX6MQjrQ/uWF5pZMwbWWnwrursherZH39yvGyhicAZh/OvnScgYBJiSsNJ3OtD93f209P2bTf
OiIt+JDBJ8Mrl/dBHtpguZZm2Ccvg2rBKVCFwipT2dgyvxyHEEmJLxCuWg7olwHsnAAK8rmgMdoa
a+lv7k1UqTVuMVcYqjDmpzMQKzz2u23Y39CNNnwxCtWN9S4UZqgHH05IQZpPyi/XtTWmOh5rvD/s
lNpMMzpIhv8Vf+rLChOP3LIDCzdZ6TniATA9W+TsThYy5g9EQOaglXeuny/Hl2gr5tBebgBx4+6v
yaiQrUSvKTOaxEK8TI5mPP7KKep53MhtVhoSu4QnR/5pIVGnqu6vL1lhQ2xAbDDRiT4VXzOwe7tM
2PBZln1ETXmSdwlqpOVx9Kn9yMX0WRZFNomQJ0kZwihkvBCekN9sjzLTBAEzibLLazvgVDnro2sK
DOMnahwBgcneEyxO0rNPStwcyCgaevppsmE77DereeOOQKhAsNiS8P7C5aib7+W8GVwkdUQush91
aym8YUMGeHnPJRWRXBs8XcVKS6CDdMTle8UPHFqiNw+WD30Mkvhib7T5SAkj4GxbpQbGDM38nTIK
dqcTlgXfNUFu3p+aAFf/8gocza5V7tr8LxVRxFVolNlA3KRJ6A6kRZe+hg/FhhtCCxyi3UIKYpa7
X0vlRYt/lJ943TStwlZ7r2Br8W6FQtbV2/lhsMv3vse7U1m+lnKojIgC6aNlfat5Q0Fu/jG5BK6w
a3547TaPez88j4vrLOz0FP+/8FlHaxo2lHqE9uSRmr32WZ0OxfDty9MQsvC4D6paADc0GkCG+7kY
OqbsuVe9TNhwCxtNEOrBzxoWXjUFc9VckHbf2agfYlSjwySRd1TotAk+Cg7JDz96FTi0z7F/b12I
JaKRN0aM6XVpUBUKa15GGVe04yjgpKMiEudx2BcBmS+ZSACSTWTDEbaw3yvHFt/V0W7K+iMS5WUg
YejMbxADqhF9ZAKFB2A2kHWYKzlhJwWp+vxK7FM3+DjH1Oc0zgoCByIBRWRLEIWPCGzbaxAmvx/p
oowb0xjUszJ4NhnU2bLmhrajIZ8w8RULQJRLDIyEoHCZRw8DmS+CJTiQw6V9IQQd9DJXw5XrryWY
wYqiADr5bYRihr/t/nXGGrQYRSgAcD/QCOg2raGsDRPgrconxIPag8AONNMERvR2RUU6MUOxF/gU
9LrrneyvyQYxL6fjUE1/2AUDlyXe6bAr0om7d8JfLIQ/tXALfXcRhvXBADrmIbTwOPa+ydLkwanY
Kt5TQlAH90Cvl5DrgWm1fSTKrWNL3jemCzi4/Vxz1To7n7lsZjo49OMGw9QlvC1OV3LzE+JoqPlQ
82Ld3+mjG9qwa3e5Xm/DgvCKuMAuIdVuDAyNjj0NshG3Pebpyssx/JaMzw1onjXdkKXSjB4gLQ84
6G0wdT+ny3gcYw/3Uhhm0/JxSa5t2UgQf8uHOaVE/7e4Ss/UY02ThtYbNiTAmejWhyUbKhHNP/p7
ziXJOjvj3T1W/PqfYYE3MsJKdb2KBBprl6fcXaAzxNlWMqbc9UC5MQknfJN57x0onCWcrJ5xdjgi
TisCfv9ey6M6jTrAuml9LthFZ72Vm6FwSeFBXeOl7ORDfrxuiC/EapZJ22kGpp2UD0dXaBds6D7q
5eHqzQgFiv06BcDeZ50zQ/NShCYrchZOv1IJJBbuXQZMso58/isTBxb2x2R+QD3hymSKnTDK7wvP
lyR7thpnig/bhB0MjBYYWsIcqrufunNotMPJUMljeNgcEo7R2s8RmUHUwz15r566j0F2cMM63TfB
ISxBH5cERmaLqu2zw+SeR18ltg/5U9DzFknAebrK1+Hcg/U0O2Qw1UaY7UUgU7FJw5/oZNS7VJpH
Lf/uli3cV2D7Nf/LLGDNG10Ybwfyt9QuxJRdXDblIzQQOWCqoIF7ChdimpHYfB7a0fx8OHmKi5zF
s6EFHXZRWnGCYxnBF4jraCdF+fdSWDIarovbFAPuZ9512sVqjLYtDBRUHkoHr1MDCrJZGxufqUeI
n0A0EqCL49CDzDrGH209ZOY97RCZdbf4Y44CCwZIsD/8guUGLSyoztICyxvqrpfW6bP6O62YbGC3
amR2hNvg1JlPATA5bR3AlucJniY21O5r+kMeNcaelnCbALrq+eLrk3HLEtkyMgywpLY84Fk6XK7V
3hZxXoRqBFCZ90gB46janKlrg03fkpyYjslY4jTOojE+jx28JMun4d+rHp4/9EHa/4aT+QK4BkUe
2Strbd0tg3ostGR0VPX4gJgFliwuVokPocnb65IHfqGoU6MZvKRibX4ZR0QEmvPt53XfB2Q5+Noe
yaERZslOyETjqRACuLjWAhC7kfgGuUqU2ae9uHe1Go7OLhT/MgyKVE8Yroi2gOipXIuFyQ1ndQQ7
KrHOkUqWq2P+YKQtR7Oj23NGhQ3PtSZM/Kuh1aGcRr60RL/GgQbMjf0uPCpsHO3E9w2y5qwRpb5L
gUIouzOu/ASTgu8UFsuQd6YPGx2Dk3xsEcPr/oJiUoX6KXzB+wbAzH4+7wqj3XcIoXml6DIAeyeb
Q6NPS9JXv2yT9IMo6mmmTWuucxfFnOEXnGYaArZKCm59BoaV6tXtLgJa7B8wSv8GCTSF5dBJ7xfT
svFlMaP9uMO5IEZAnrJWvg/hB2x6Apt0JFj+RXBk+tL2E3qF6PTHWpw+TEXoZySq0XuMUBGHRfzH
B5TKCs3W8QKwbGIuoMQOgyb/bYhnoQjcFFeCu72+tobfxtAoefYiyNrJp4m4k3o5enULiRmbRrI4
mVYlbQNNlBjicvoUeMcJLOfwbdI6/HWkJVEWLcTGo7OEAc/RF16BX3KCqmAOhdGtJgbOugAbvAvc
eMGAJ6F/Gh5/p9iQA+CiQ2s9D5lTwXjeVuQ5VKSJHjziuE9Nc4tf7v10nZwRHYeNpiv/gsGxL2io
8Otj7Qn6KtSAqxGU/NSU6JId0WJH/QYaVM+ohz72IkQllHWP3zbTDmdxAKKuxjPuhL+TyK3gQWGd
VRFc2ohrA3cUl5qlXa3v/2WTY/nXe0HBVVa5t+B5A8eU97kj8pckSXvyWqfDV5Hlo9T8wSY7IXHE
rM/5/zyqFrF4ktu2mRR7p5rFhMwb0gswN8xOQLS9bSdcQFAQ5l5lUpk5gi+bCy9mHok6uyFUedf0
4DNnDmFWLAx0M6zdoWoNtEqM4+xw0D45KOVP0RIAzJf1lP9oVpJjZRIkHIeKXckBHyzJxVEe7jV/
Aj9k6KKJyCc+nDGTkBvOgp78PTFOa9KcMtf0jVXfaBzv4nQU/f/emiPWEU7LXk0QP85vm4HEtePo
ikLhcMOwNLIj1ExY2FFUw4fKieE7Sb1yvrvFqlq+AZV4r1dl51Prc00BYN0SOJx+NVMsXWcKAJgs
lvyoqUXTWSk0yaGus4lSm7kqiAjFFhLN7qXRhwcr8wYJi8DTKHC1SQ8xsU0t9jEVHzV7m8q3yq17
n+W68PFB5qL4OFd9+d06Djejt9HGnPbr4e9Ni+PloVxx2cjYNK3pPXMzhg5dLPiXXk42n2wjoHln
oYr0VUtkZ8nqjv9AJpjTguQZDVR2oOv7G9Oh48Lj1vGbVbRiT7uLYoUR2ZuFlNVQg19YNo3J/yg8
9kOKXvuCtp5OAEe4jBxt/9v4CBq3kVIgVALs/7N1+J6SItkuzPNkTEjEu431eDKkQ3xsjSSjkKdI
4MA3fPGbaz4s7zYPvclEQH9yzn3DkwS2pvYlJrtXlLB5W7gguKR8BQSTwc525xqNmLE2r5Eky02N
bzmh9uVme29LBz3vbkQ2M6Zpu3dHpMFr18X0Co6r0tuH/zcKKlmiXVmLrPMewW9oH/Q+6Tp2Rnzc
Q+Icc5YarPhRt39fuzWjPhCDKCuklY62HWVgAPpdfB1XHZ1WHguwVHBBY/GmhOY+m0z+ussjMVYF
0ltZIlG7vgjCla713FLqkJlDrVktlDfv3aZ2CPcRq9224xhnhLmdpt7doil2TqrC+TF9V3OU3T8G
yzubWCb+wb8Gug6pBv2qezH6NwT/yJ3R4BuQx+ySK7sWG5tCtDeTUfYHLvlLwOH7uNUTKpjL4pwK
ck/RfvIU/cy/gywzVdJtVsIW6Dz/VMa9Rj/GEeDc/uczupZAf+BYMrGGNkPcEWjbudXipAQpAgwm
InZ8EMHXpz03uM9tJp/sM7ngz3Zpi/7ZGgardUoUOnKJDVdPBYuYBwtV2MGIIBc1iGqA6YkvlM84
MjSUZNN48gfTNn6BYYStQ6hookzfgK4pTIg9k4URbGzg/jT6yMIwcIPECg2mFVt3rrdQRYvzEOs4
MaQc4Wvb7HlYFGI9A2Z3VN0eOauAjDbZP91bjdMi/LVrrzDlNQNyq/uY0674Cz+K++UZ/QROXhPu
IojWOI0aPDXVrgAN3f8LbpxhS8uXdoVirnojp2fiVFT8vT1ybD61Ey3XcErS852+glaDbeFNVCI1
5jApuwlODpndJ3ncQOPe4JMrwaEpsp/J86AeXGJWZWjh7iaqhDSorb1OZk4yKnklTJjX5RUPi6vM
35lyPBuc7Rb1oj+lef+4xvtz71+bSEaX1F5d1E9T9Hva1DTdY91jB3fZyIGmSZfHGcHP5kFzxhjB
FmVp10mSswi0HuE8oQUEWoGNU8JIwUFbMjkhzjMeuwOVmyRPfNKhB6LktVZBRty866FRuX5ocWTG
wpITp1uT1UdqbVhqaErGNOdpc29vjzzyS0EQxGz29rrGPCGLnzWqrpKL2ZEzv+5qPDbxWgsYaGQ4
NHqwGmhpGTUJ+b4/fD2N5YN/S6UzRfBkgrqUovt02YnURiNRHwD8+067ksS6i64a3EQkbgT5/J/x
KVtAckUdqZxpxPB2Fkw0vTaN5mArjAe1+MFdo069TQ9/g1jW6OTBe7TIkFnuFZS9BLOEQh4SBXFx
DPezmBblTK+zgWoxpDcnlT2eHftlWsO7DzTXhiFkAlLcEuk6HmvNFUSbZ+nLWW2RbkVQXymsKSrM
p5SDIU3f2gH+bxEri0HEl2xZpcVqCfopfJnlHJHsiGmfIxR+aLiISN6ASidwK1cAjJUAvlf/IL4N
GSvwitRwkY1l2NsPW76cVR4l5jaGVwCtg02jtFNPNxqf9rY0Qky2K6O2LIYlUNAfEhj80CKasFKs
v32pf0dHf9uyXL6Mv/nRVWSBrxYqfYb3op+BTT2c9AiOsS4XQ67djwlUFD23A8gGxXtL69bh7GQP
4tS5or/9Oe5MK7xT8XThzYfdfV3qtUdpqlfSSSJx3T7AtQMg8tamapR1MUsDBbFZ+KEN+8TPpBBq
CyePoaokgl5t0Xy3T2xbNvymemZ4D288GDb1FqG3B933lqCT8Jfw/zzBmQ+yVVNDVKmZ62sWARnK
SLfGB3UozlDsk/CPexMyZYV3EPjZnXUNW+gKxiZMcF80RndTOz/9ITGiEfn5pLS6EhcouLymfM1l
mpVJ33FxY1GGB8gs4UCod/9VSOMtVHxYqd30zMciOmyK7YA/7NPwlzBHjdek6yC1eZpJZLMZOZGO
feBv9pexzmgpjjhYpd3epXiCp6iimFp+FWD+wGe/YJSqi7jGyX8oyfu5TxDktIl545Hv8hr+TKUj
oJPwnIN2aLpyFfhcfSdHdv2FX/4DlftDo/akv5AftJEXp6RaEvAMnHfiqmGvkZTNMLEWB7nnjUkZ
vkdyEd4aUYE3x00DssoXR6CMort+NVY/ROoSaMAw9KrxDYn0iandXbKngonZQ9MzJSl9CKwuWEiY
NnHjr6+5jRs64b6gmSHFgMTJqqs6ePuTwxcpZ2mic47OVsmEt5dAD+9dqS9Bwp2dkPxumUDqHg3X
hxvoiEFfCgyDBO85xbTRUQ7N8hj3jW51YG/ha+dsbD4pi54hjPHCsnCt/BMQ72wzVKCTwKzYfj1K
tiLPWrHCqqJkQl78BYmMZp1yKXydR/9xL3TYatLp5AnbZe0AYOm874Go+LwnN+4lGJUDk6ZK5pN5
Vz+1buf6L0zeSACnlkZ1S47lqfHSncS717Wm+UkWX+OOIXGgXhsR07SIJVVlHT08O4V9E6ZxEXIY
WKPT1KmPiGZrYTz11I0WNkLK9IuHf8cmale5twbC+Hq/Yd9cHMQojS8+zn3JcXza/hVPa8X7OCTb
DC1CBK9UydQKV3oomgZ7G1Ooiog7n25mv9cIx1CZMOOeyyHm0AjSSvjl+yzl4W/q6FM+CsKqO0gz
w7pbvCUSFtC3wx5OXDndZ87JYMsA0NceKEawIAN003fW7vvI6IzSesh2bVSgT8ul3WPPi3BSbWoZ
vVHAoDyfoIsFVNRejPHPytW78Y1v3QAXRrjyA/bwB3ZAfkUzBe/3TRDlctsVINxzkWzzmpydI3F8
jiQfsLCJwIQyrKbgrDb27wy2y1yvAdhph491Zf639QKnIG9oYf/0kD3U4Wr6QAwoX2qXvUQxsOo6
OzlOUw6+HqTaiLN7xJUBIld7K57Is5y1sn6hsQH16gPjQ+WbpbqJoc589hajFJvUSQteIC5xMrDi
uviO6lS6HFPKamQOkcbXSsw7yioYDYTbjf0Ju207x9WCTpAwWFPcy+k1VfNDeQLiFYyZlSgwmW2K
fiqWgVZfQ1Jps+fYuNhSJenG2ySaX3yN8YTYjNdBF52SLWkMu4SJcJVi7tehnM79gml6cS3ZtJJ7
M2EWfqcNJHevL4+cPfUQn7GOaAlOmQL3zNQcAad7SlaR0QbG+P4XHiV3n7jlWMWKflZ8gPIBt4M7
HFMC+69lZSRXU5JlkFzL4+/ToIm3BCD/8t8Tbgai6BxXFGtjcqQp/rLj1L//1gZlUH8r1YWB+KpO
meHNCi7C/JEUU2d3lBds5riAZjaAJf1csplBCW5Q4ldxe20aUXNqjcjNqrddeaG1jhELV2PyldKP
d7EqNzd3SL9fpAjK5mfSFFTQSEtLLLFz3bbUGNSbPV1t9rL1VXd/9RkLrDSFBL8Od7C9o20oblQ4
OwOGx02HoPWL9e18PQPXyd9nwBaeGs5vQi0eVbe/R+Hd3ECs3bjZct1rsyBqs/oUt4UsKQtYcF45
LXEn+Th55DBN29sthGotb9M3MEwVd1fGMhYQUaH8Jjbt0hvCAsJomhi/rLt+txZTrsQIdAGe4HaT
CojcWCIXCdG/hqHeS9H7dlInm1TpNaA+jnM0peyAPx8hy4PEreEA6VAhdyp/5vQrpmof84utUQ9V
IsL6oixs1VPkDJn2me0LjmcPlk6JbuumhCC9A+v8ohohbsGcuf1P0bWFE3ltaD5+XJmGSubbxM6G
EpUV3sJI9gr2wlPriYBa7OHSOc2202wQMBFMNxbWlndZCaNQ7dgDEExZxqQe5y2hXnLFx0PnO6DG
2+CVRbCStGgz1zrLCMLyU++HHF2iXpUu1U+pdR6pJV/hek7PvArNP1DZF6/L9BCn5w9KNl9DzKxq
PzOHpoQ3SNaWvPltLDX9ZanW75MVEr1QgIqb34uny+NFERHQrHIZA+Bj1tf8kehQyd0m1aAxkQw7
0/2jL6Gt1QLKtUhSKn31N27RW2sv0Oy10cog06am/k41TYWMxmgNmQsNtmDNFpcZrmaSh6+2aVnT
LVSGfXHMLv6EnaiBLwojNid/9587reGk1veE4zZDxT8+39y6wON+8D85SpPjbxaMp4UTKTHsJIgB
7Y7a2EoPh56rH7yyQKtui7S+m5WAybueZ4EeEA6LuKm0+mX/Q76XIBYTHSBktD1rgSKr/bhXAmVn
qk5W8Tg3+XSYI9qSZFcbK6I9ujD0WLSdaoveryHT/mbgzrfzg/Dnij43SvTaFRN6p/kkTll+PsWA
qzRqVhj4uiGSN7tJX3yRiHD316l8KgzYFV9xWZFrFwr06Y/95xBI/bA5BE73247vDDEAtmlT2Owb
NqrfdRJZMgYCV2vFH4xizGmdxZKFFND+5N3Or3v0fQA2ldPe7Iosf7/ygZhSeYYB9aPvnjYyPp4d
fGBjDrAe1gjTtHLcePyPXk265v230Rjc6PtP36elCcHmTBhEIU+5ZsnWBhhW/WmBHqogGFDk+HDQ
r8HwlJ9FPfFcgYPoEg4tlcpf/Wsom77LwqpVbE4HIgfr4ewc/Na33Tn0gJH052GDa/bUKbqwU0kX
656oiCMrcaXGaMgs0Rj9MX6dGDlZYsipw8ZtHIIrNkNuqKTJc/myjWljNNJYt3zXYR3wbtheyJ69
6kdtfNo0sZ/2SbN+ufkmttCYxo29WMDlfMrpAls9PARzB04IKB+0AvV/zrs1rrAECMBEeVvl+U38
L7A59enfq4XgRAjcdnA1BYcAGBc7DL3+qcKlWLo3KzyZy4K8ZPoMp+CkAeBqsidNtLrlYTa1jFMH
1LP/ebh4AanQFaRKui+96bzfJ7QpbfobgofOM9j3a0xJgdwAPC6ql8VRcg3cEWYece6QBVqXf5rf
M571syC9uVvPa9zXeQtwyxVnvzGc1PpDj3ce51qZNNbJFepjOPCO2C0FeCptWhmCHNlpAx4zo8+x
hekVu1TfuFWxRn2mS/Woqy5wLwOtpk5f05nfejycT7jhzT7zGbYzqbkQJlkQrzmkSAtneAQmE5iL
ig5JG5fU+c3FaaBToS3rU1AMHuYi6xumpKX3nIw5iNiym/OBRANOnw4+j5vQmuVbWxXwrfjf8++8
JOUPN5Llq0iWcReTEjiFwBY9IuoNqeDjG8sq6wbJvv2z6c8sOjS+/Co+Z2qC/XNQ9idk62lHXHzy
cVoYZni8Mfh2M8NglKq0rn2JlTUCLhDJG40QVf3AImzWNHFdpsyWi8qYoXXIvDLlIjoeO1oGFb9N
mP6g7efVcv00t8CaizM2FEEZEpFmEgLoSEwCayr2YRfOYgjVfz4foM5zm/023s3lYnYDWL/EbCji
4y5mV/5vjQIlvjUEgc+HaIwciSnQ11egeAATcsSOhrTt1aAB0F0S6aDhx2Ec5PypGHhn71bhpuFz
fR1A7vVeS2Xd5pdIp8Hp580K6es5H0JBMExxehf/zLMwWXb2uxgiCFzaz+eyb9J3DrEu2CgB+NTy
5SbrVkt63uTpSmHnzquaE6UEZtbZGW59mD58mQSpXqUYwRWmmM2ZRchbssdpT0cH600Qj6OVmPq5
B9K5bawOkxE5sNmJTq3iiTEvv+g2HDJQdgZDhHeZous1jJbVPNvfyn6Y6KU8Emc5UFteenOuzF6s
8Xcr4wdMS4MGYnT4brFSIE6BS80rvnEo2r4HKwiDVT7kHE46hx4EsCYyvkbGR7ZY2OfNq/XKT75d
HLyrEOU+vKO0m9hGY3hy+Zt53/sYQ+3TMWPyeD2enXNFwddb/kXJPAqbryphhqt8+AIyMpeXH439
6wh00f4vfmk1xDm6gLt+bQ3v4vSo8udFO9b4fMuwFgDpvb0RUGF7H4Vi8owI3wgolEcob6yV/eQ4
UXZuPlH6khhyFiJv2MbuFCBP/mKbS0UwPlpTRhjn6FhKmZ8E8D+kqc8KZkEc2OhpA7g0XoQMlyOw
VD6JNu4zqzS8lSHLBw9CBS0YONgTMvgDpr+n0S1T/nHj0ya08fv2sLdBADF4D/0l9/yb2alLbGaB
NLTzRkgRuHJvJ5a/GRFy41PnZ9D6M/B4dyzOUnC9Nr4bihOFP1fJkNEGWx9IRmZluO1RciIdMegO
dL6RkDW7S/B+ZEVc8iHhBJCzEa6hRcEsT5oDKxFl6xR7mVMAE4Kaes9gJ+m0xHswM1UEvI7fLffb
QB4/H5PVUQyPsuZcUa5w1qC9K/dScF+Oh+CdT+cYn293fEwPPGlfiX4sI32Am2qzPhVEI9JGRTIT
8Lcx3IpErMoA9c6kw10dEqlxVeh3NLjKa13wed2hBiPgMzJPAk/u91Kyd1iDo2NPgpvuJ5yEQl2+
yiDZO5TPuM8lurkVmDDpe45NOKd60rLkD2l46qzqVKTxKINu0epr2XIyG6jrFkOc0Z+9DwoUA5na
vyHiIf7kUrz4zFak10dWZr1oPRe7pPl/HijWYQXYV213ANlM9iiCdWt5fH1i764MOeMcMIXHvMS8
5ULLAt8dOCy4zigKlx8KDqFAQxOBvzmUm1FxmobNHf88I6WHsqLbPuwOecnnpbCilT/BwyR+5wr0
yu8ZTR89XyXYlM9QW33BM7Z5vIzAIxSoLz0FM+yvj25UDnYIAUSoBk6zfEl+V464f0PCmkn11+8S
gPJ4PJp0kP1DTXPL4ysXEP2DMTMSE3Mp/o3WLDa212NqrO7kmsI3OT27SNGHmTmY0YVloYWVvikt
sIXtpfUxrV6Euwo3xhs5+IWZnjsjEPIm9cIya4EN5iIkMMNZps0bCvGiFTxfVvzcoo5k2UL3G5aJ
QkjaUU7SJWdkUsKYb4dkEbKhzLpaAhj2MWNBEL5nb/gRXgvqRfokYEBPrSQOLFKoKdD3wKSUVlp4
DvptLUz6OGu5ESOf/pXNuv4hcDO1/RbXn9Y7Yqa1N815DYeFaAaYor7AhXfqGGZrEx0icgV2VxL8
hfe6/fJQwRrOqCWpqQD3AQYU+DYWYeJqRPoEESLW7mQXgCObCtirMov21eJEe9NsgMoEKFgEwjSk
Q2hrNtuOLotiE33jKRP5UtAX7iagc57ik9o2tyDCz9v5F5L2MJGX2e4G7Ga3/ybE9KB8KqSIe9Mm
qilPJ/8JYjs+G+xqfKKwSNIHi0gmFZHL828n5Py77LkHcVzV6uacsn/QAKWGruzt4bajtDOdmStI
vsAdsvXBtKxiXRMOSXC96+k+TBOEAOqJGlH/WheJqAmTnHcGKXauRptx0eBGqXvA6E3YDcMgSoG8
Z+v8kVO+gNErZVXmFLLC87urpWH6WMLASr2ElA0uve3NoQEhyKPWr/fPYBLbGGLeFtScvL0azaIw
m5jIYVzahEtuCKZQbWo7aIuvXkb7k7dL7lt2uxvBXw0nbSL7iSwsSxtPv6gSWRpArB1Kna9eR7Uc
oWg20B0K+6yFhv1YQz6Oml/orLwSoQDckUN3rUo73gSjvd6IiLdW61aHkUdM4MwahPGYv0ICiKx2
ktWV+UGLfA2QK89VwUwL9gNR/5jY2a/vr1J1MSlFddGOGWXPJ6cwQ1opB9nZy8gZQcd3RaeuDCnm
4LMWMRPg2ivKI+yANOXki2S8HwS04Iy6So+B2XTMk82TM9TklSNWXX0sfiV7nVBp5vVMAX8sJvkT
Q/plVABJlVLQx+F3MEBd50DaldR/HL3qPGL4R48apveE6sJyxDsh7AfQvTNMlEzsN1gt4vYCKMiC
xarF2kxN0d831stom2vpQJ2i6d0NweycnNnrpz+4AJo0yODGWwSQv3r1cVNZS0FxaDQJr1I+pV5F
bKoh680P0kdVFtBhzP+9Fn2K7xH/JPK7zEJTsfPtjqdGUT1dV2saiD0c3jTxflONuTQKUeQG5f3O
Hyr73F+eq2FGSGf5Fvq6SQW02+zySol3Cj/70XZyh0lRpUIB3+Hs+2UgnqqaoWRCiRi/pg9p85fc
1CXo8j8zQ02c/9YYoeCiHSJyM7pn7L7Ud5ge1dRs/ZwNG8PFwFtR3wHwbizJloormJzfQvtsPdKH
C49BIXsZZWRZUc5LenVSA0uLyTL0xvmlGwbRL3mo5kE1V76vjQtaf/3fXBnnGQmggmaW0tt7TBye
a2HoUrI+hozjwq34Mdp6Oo0MPsE4AGy01lvkpjjWBIWMjhpEjU7CS2haqxBJ4Iyr9DJl+GCFPhNp
J21THA8DzePXKtODgz5ncjYgD0q9W2WF5gAiB+qfnfDOzTzfEl9jjN348XIc5bSB61fBaccbc3T1
UPtkok6GOxB4w4TQRFIb1WCKNYzWcqx2uExzdZ71zx/Y1j7xabrxV5tPQbBFR8127PozqRaETaQO
LjyouAT5eIZ59AbUQ2M13YJBUaMkr3Ct6ESFWXpG1ts3QVSvvKhVJVg8yu3N/cvafYGczeW7le/7
ryVu5EGiquEVfA7V2QjyCtdjq0JLad/GySH0DtZMqoCwvEX2JNB1iCFJG8jRK4egDY6olNxiS82/
qBGaJFGDLVtWfB9yqRyU3uG5eZXmkQm26JB2doQZ9ZsH2wuL9gk8YYyxKDhoh/CCGMUgb7OX0NMB
pwQfTfW1v4K43hfRoJSCBf/BN3YLDLJvckT/92O4rkKJI5TAcb3W6bT9XJ3/g+XCxG2l3/ttDS/D
NlcUH8riSnRNswloPpbo6HGH9Kw8ELBDNHkraMyMbLVVzFYtLmOG5KInPoKQS/+Gc+/2qmqte24G
L4ipYwlvcc/WxhXj34D51OfZn3fjYPCijCaGjLZeSA9ADEczuMaeYlBTbdrUyPNHwYlFBLyCZdlB
JzL1tDY4pTUrMSFy/gkvgAd1NF/BxrtNewVY2kKQ0b1jbRDtykpTV8wYd79MB/Uv2GwmsmQLMc55
aPUTJzCRa4741js3ThjMwE2QUpmLXmxUtOmAyVl7JZhvM1xt1LCnuTTckGlhsfWDoy077QSRkz2a
nqXlG4/OUqCtOKjMVqkDNtdtnDBUm2PhR2idvUv5/hnbueHuQrmIM72cLINjj/stxLw1IW7LJDYO
/jdrlJzogNFi4dsYsn7zX0TsWgmEpMoAoI3amqFShU+xbqEqpnmzNO5C8FORKcqZJiBuXMKFkf21
EOm9DM1dmI6JZbw69mdhq2kjaR8tiafz4ZFfX+6586E1XO/jizWUzuKrY4PtGcSf/p7zhDQJGta0
d4proFtUj2Pz1+kkZntiPVVRvG7u5kcEt1pBhRplT7CoMPb4OzsBN0BFzEOb9zkjdS6LumzJKiKM
uniEgEYuRVnFGz5M9ehrHitEWXnvMlQdyXRDX8mO2/h/SXWS4xVpSWqvURM7AU7/HhR1Yy52didg
nZfGAeuDoKtsQMi/oIua07IK9sP3aYjaXg27IiMzpGFzxacLAKq04ri3uJWGD9nGQUym5szV4u4O
wmfm1V3/BC2DaccVfsdxlCZzaWecXdvaS50ikcvOYAptWjvebivlNQOiBG2SSMrr7PzzwxNMfRZa
qQfgyFMxylAvnVxfO/MZE1yS2nAt+k+PUFKE534DpFpfJKZ6aFHRdeHTscblgjnXc+D2LnYbXGMs
qeHKrTnw8u3URSVtQ9mkrH7QP+7v1i8g5BNsMdoydCvFmRDoiCiG1/ngfh30IrCLmVa6ZpQC4h+P
tDeP3HpnT8ZTpD5zdKX8hiEkRhnvkrjs5UERKV8Qn8fadgdZ8bAAGRtCcWNtCHLXKQo57YXzJvv2
U95AO6S4nNq3Z8Et5Xs9SEgJJZmx0TRYltUd22E4vps1CZ2IxpO2F4f4UK11fUcL9BZrXhMLihJd
jxPuMCavWyqLdNAW//g4uXh/Sv6F7yfux746r1hA3tb/kzSZPgSYVt+Gj6v686MqdBCm/hpkLwGK
Wtc+pFVBdYwB4nuKNI3MrGkPR5MGCCh2PPWfDJuo9kNmb2+bzPu89mYG0oaV1tZndffIwQak0v6W
TeYGzE26W1u3UzSS9KsRA1ePWlTkbwJ5fysqTkca0mJcpp8v8vV1KWAHkiVTPq0itPixjWcYCWot
q8jjcKRAbtGG3/paJirzYVJ+kPrLeXIXmsBjrJb1e0Egbava009Gt2+1wcIQFjkP/EnG2SdNXCMT
vFR32FyqQ6bYoaonFA+pYKknb7ckPUgW+JnsUSmfl3ItPutXESjkfc+49U06FvGb7kGhh17NHk8v
WJ2U5zfSNdkKrTYaMTOTil4s8u9AEgpoUC6YlGV2PxANCnCx6fjgLfTzpdahUjeEaGdXtUVj2Ztr
8gy3YBZV/gPEOEa+Tyxohr2vD0OBEEG/oHx+bsAd2W68i73JzgGqGeuN97Apr+bWALoi/qmG2roG
Tnkl4jkvMxX7xFFgRCbNgL2BriXA5GX3M+pXq3lMf14B+FmaF/iarvnzl9dcqvhTXGAe0VF5eu41
801XI4EdjfIJPtRHq6LCAyF2sfQxuG4IEUM0xX4eEDk703ZGalys8a6/VihVUecKumbT5hPQuszN
1QFhMoUKNqaUUImzBgvoWWlAkE9BFspcwVIBHLErGRzsfcq8aUUXMWtTpCDD9S0+WINY08f9SuzQ
mTl4jQA32y0PuU+LUFwet7OekaL2OUB23cwMACFWypnfC1DBMnReqXRte3YA9qJ+gLOQrtkyfAJQ
n2xlKlOjuBxp6t4KYXhxxJZkCHu5CEbkEFtOLeVOgZINKu5xHWCLBiUzD+m/td1uxtaVBukwt+a9
MT1XT4/40TyiKCULKs59HrT1BWiy+GzB9w79cJT9ZVhaWAdeUgxxmsluz9YRpOJX5j2ACDB11nDg
HgRN1lHzS5biHm9WBHLkdwxghxAvCJ1XI4XVVwbXdeYiJ7qbUE4mlA/uI/3QpUsVJh/A7++J7Efr
8kgtqcCt1CKTw3hjt2cnTRzNsv53LCKGbVCKOhzVS//gmQPujX5vzuJz+qUh6NnqdTWMDCSsuDWK
kAV2Mqvo5sRjg0QRPalmlS3oMa1G3zmPn73xyPcpTiC1aT25PL2Da2NDmsS/jo7+/gMetsUBxteC
o4n54N16uMbw3PE2nWs7OFgq+F4sZEnMk/1uX1dqFFXQ6DyflGpqRX3oN0sw+81jzF8YSTDAMb4Z
JukqQWhJ5wmpJTyamainhAHIWMwjDEYrRTjOk8hnIzqOoe0HG4W3JoepOu7NFvGjFwN2AxzmrHag
JX1YwYV7Ux8WYJ7RKDKR3SKbet17B0T0JqE24qoPFqtXoOcEYHlqLSXKmMvDxMTVLsgwONM4hPs1
8fnFa86/hp9/9Tqo06HkCYKaqmza15+cZCsnhDoXnbq44O3AxGCvfw/LlNvYvZtMMGycBKIgQS1t
bvIwSqXX+tXLkQFxg7Z+1ijnTBLL4xg1wMJXLGXN6ZqJKKp1QTFqbxklTmcccBENk4SBRouSaDhb
wV3QLBfdxgpSZ0M+G1oNVlKRLNPRBWkviBQgn7bddNwyfOx7cWBgF/sFIFi0hGetjCYSLdgiOSSR
JUUdFINjeVVmH5pryHjdXXvYqRconzZ6Wa9PQmYe5xnuWqgvotjYnT/DhYeX6xyvG3qw/Q+NsaHO
lCFk+8OZa3Sj1++KizwS+amb3itCsQkPD4gDqC8UsRYd8lHpfpEiY3JUe3Fa6rEYPBMAUH3ivVnX
JICfbcGS82SQTdj+nJFjnq9JwwuHu1GYSWulWzc/MNucGmpTKglFpsoVVY9ru/2xhT7i6WpE0cR7
M0XxEjTCGks1FxMV8abykBv5l4iYXgu1ATRJP0bMpvMf/zV4CujmbSbQ60VhSqyK8nQ3QJV683tE
0OQ4rafFWb5yRIOP0r5gcI/B3kSYs/r9W8b8gD1/ClH4shprll9dnST3PCt3/4I1gDLLrXYPocph
MkscD8Vfo8/p/IJ+dmFEa3uM2W1u9r8e2+vp7bE1k4x+DSJTh0Lnv96ORGiCh5ErQ+2069tZq5u0
MAmWsNHihehcVHpb5SRZyxq2KrFctj+ZQ9DHLS73pRBhuz4fSTI07SZzh/0oLHNgyrlP7HHvfCmx
JCjqyqybWXMAoBaHb2aWnXoOOcZdws/8xcOwH0UUtfrq1IDixqHDZ0y+QUBfsWahlT8FjnDfk3Ao
pCJty1NpnBhQLKYWBbAX4c2dBule9/KPjRi9aa6iFw6HZMSx9nWotoKdVO089bahtJlFWYP7Sxnw
/ujTZgil7Ecw7O3IPMCK5JiOYk4h+H/zb94tJcbdk/REvadVeiU4iEbi+yjRGk4saGU8Rif/an8n
GbgoJ1cwFl6Fhpq8XZpyPQ00GbzkXabNYl4lEXiiMwlXQA06dOYUqR5oHQ2VSXG3+g7GDZjqEkur
Ecvu+++uv9ypFJ66R8sv6TgGaXKNJZ6JE+B/ix7bk4NpWLCttvJzR7padxTtfjSOwhhV+57FteHH
adDMRjJ2ZKJkUT8X8LpC0HL9tAaD5JIkkVduYM7A3v8x1whVPeDeMXAXoKFXaWn2KNpznD2Do3PL
Bo9psoUSskL6Z2qFqltry49FRyHtcJ9B4yfJr7BnYgUHOdoWIW3bmgJK+BhDu72EqrMkgQED2o9Y
fGANzbKnzbaGhtHccbkwL54/t3WJ+0uHPA/pfCxWy8XZ3Rqc/c8j0mWZz2cZ/7Rr25oNb+w7UEUu
AJaM1eQfwN+RyCTzOHAGbZpcYvAj1jUpA70uMPoRIbMW+HPux/3cNPhJIpW3XpdgM66ltK1n+2G+
uZId/v7kA7dYTWW9HRsoOAPa4FgU0LCcocXVpazmFOIiB+Y6M8jX+4i4XjDvjbbZjahpXv2noxtY
ehSTXaXgDTSeeoWEeu/exOxO8tTYslLZAa0lD26Cg0XHycwm76+HglWrdxT1Ry0XAvddc/+iq0ZZ
8LeT0yAvm9+Zm+DQ/C9QiiExDQiWCGdUXls54NWuvXyzn3YXrqPamaHDn73MEusp/TxGYqGBxHsa
fM+ZdhuLbrvaEuudIu4oX+4Cryn4cMSEssJkv/ohvFa6Pl1M7HBzuf0iLw+UqoQEAA3Hujrc6tPX
zr31sd1RwfpYBjRji0qHUrrrOQJpsPLcXOfubE33Rq1GCSVeWLr197vBqDW/QHlNieI+uZKPUB9S
2wDmG4eaJPYR/h7c87ek7dQPhvXrAgHKhCvErUdmmg5g19kFqhTxRK1kbjkKwyNXs+9903TB2w+/
HMUHKBxOb4yYW8OPGWCZ84f7oY6qvvdmZPoGiuXPHvd2fpEwTQ4C8em3wjxD6W/ifLrkCIp2wOb/
jszRvO1tAfytwZ+/4Xc4M3gJuHVW8CjnswrrW49BkxHweCDwRJbsS5gnAsdefV/XciUuxN3dJJXT
A38KBASqCFVl+9UfB9nBZIUMMspKOKTWMdHqMEeY3jv1CUkYrNo8MfH9kfcRXUSFf2B433gj0j63
zwXL7A5mLVK10nQRJEJm0y0hC0xIdW/DG3c70byv08BfLxViuRmVQbSUq2J5ZVQbblbAqU9FsNiv
8mR6nyUlexF0MjhaNCosWuGTxag6dhcf/GRoN3UA+Uzsqha/Bc7fO7V89EQ9uxmWV7edNXPC4kMd
zKo4ikLIVVgUabkyf5nrbYu7o+JwQWcVxQo2MjHXgPppVR+V7ZH/QAocQwJWS4pXKEQHy42hlrcl
LlFNgOOkJMdz8yuyGw4TbSePvGOe3pLmBd0oPzzkXpSnalpHDL4p5lyd0TTlyGen9DWGLLMTyXab
mO3FtGrSvWSWByxPvYKqM7tCLsVa7X2kMBqsLtX42Yjg3ZEm5xjtzQYoUEuWOB6Iowq31jl4Y30K
jjG+C2Ky3c2x6qAApoOLhXKSRRlqDNENhhQWoSWMyJBYz3PFx0gwVHhfNPfq3+pQWtIpuquq+s7e
yO3FEEvUm89jlqzDOzg0ZqpXWgSfhzMK8fd3io/OaYULcPTEs/B5XHA/xK0dZnQE3TeoQf8iJ4jR
VotiiKilu4WrzpkzvUAp6vWuhi0kCoAsS7JTztCbrmjbnS11N+SdRy0sWreWGNcRPTJ1zayk9O2J
TTEwF6vHGEnxY/BKzKZPiJAdnudUTCXwJ/T/g0zLafqhDjaUBkA8NNSiDfQP6xFkM8QxYWcepVcC
AEXB+u3x9Mk5w4ItYzt3ItepO/ffW0Lbft3W7EeGQ55mGM0I+OEl0L+U4w6Vww9y+/PJptO0x+I8
KLTpZ5Ak2loRzpiVg4cG/cpC2gAtIMng5yfXRx4MpxIR3UzlG6FOTHEFsKV30nJA2p1L7HfqRVAe
Ig5KSoKsbtXfaybwRI1Y2Pff+odLakvh44b0zqguqfvr8WIHutfFz2HoBPgDF2GqU0v0L99OaeNn
6TkPIilS0TEac7A02g2gIQgtEdIPYRa8ZPzn79Ed1O1xI1F0vn6Bof/+xW2IHKy05X4FcuSmc3xo
ORbPvxH/LTgrR4Auufrp/t+x4lsMyABPkwinVL2EudR9tkzf9D7Upazi6hklTwGKKAO5PV2pGdpI
UUsUMwdAkMKJbO+FRfdkiG5rFH1TQKtTHuzYC1UwaXO3lriF2TRFuvZ+vIAJPYowQSGuKr4b+erU
SxblfGSp+VpeiTbEwXAdR8jwepgyrNEkoLAYUXVzAlxGQzyGiX2idTGyy8zx9DFhmOiOfRG1nPe7
GdMUoh+ikHq0Wd47ukRColpEhlWKV3N4UkcUUolN9ROnUL5PX3JUUF1AF7B6JBGBt4jGPJMAgtjm
P9grwu8PgiW3K8vsgW/4zU/qrd4cJsuvEN+dhhBRkyMd3Lp5QWCcopP8Zxp0ab+EAVRBKcoeCrgU
IYoGphYwVzDb3JZ9xW62wB2lrMinZS8ETDUJv6NXXbKKn2H2x0GomN726DPIGaf/gy4LP8RWimiK
X38AeyFnMar4qLdneIMLAvboU+k0/LDAn+p3fEC9TkMvYO4XssG1IzX76v/FS3fFRTmsUmQQN85e
3BtqugBCv6XlqAaujJ0/PI3TscYeMrUzFGfoNjwoG8vifa9PKGUTt2g3Al6svx6DdmFQeBIk51c0
khL5ZUhRLWbZik7VdsUwAR8JWfCrnG6pVaghW18mgoBRT/78QQ/UUz/tuDHGNlPyGhz7tAhU/czs
eOgrYPomF34xF16zCyAyuHcyonun4BkjPO9J4nUq2qgtgcpaAi2KGlbVgkn8WiJ4gc6qzuwhyFbN
rTYsUKKuArwYz2H6E4lRUZyAhYV0T9s+7fVe8vsisWiO0ediFovMp2NrRHoQIF8gZpScxak2x7c7
Ij+PbL4Ok8erwCkWKxu+5UIGjCgvZ63IuV8lXOW//dNwTtM1o5ZQGGze7Edkhsg7IVYpXWoHWCwL
O0FmtNstcmEaPWjCJuUz5AiCXnM5qlSq3MFoyOmjryuai+SdM0YLHaWM+LB6ytarSkRG5JBHORJx
ejqONORCa33m+kjcmlE4YTeHOom17deO8D5+cdLbdZWWXmCtrlJVoegrByVj9yK9uK9xJQaErwIc
M8tyHsIdKDFCQTKMPy0bN6E6Upp2m5OvoY2wevvanqJ8m2M0EYmBq9rMyo+ZGI392iUeSBW1tzry
Q3/gsSv2xLCUgRQdEwXAoUy5jO4QS5ivjmGHsRPnpdHYnK39sqgmLWtvFx6EUXBcWIeF9QhseI57
0EpSIkAOzfX30nnUMt5CtFdLayD1ymV6AtC+LQXlWO5mSRtYxWPhzkhU/C5WRp8qofjDzZ/o0mtS
CyP9FOgPQsvXLbWg8KyP593pdsOHLFSV1h1o5ncsBN85baj0eK1kQe9saiIgIQaZhOceseW+iXLT
1ixOCTbhd6t4htTJiulIiOuzaLjlv22OnPg+hL+Og/0wtwtB7F7haZMlISJN93svfpvrAWm/Rg1R
dj9k6zg16+rPuyO3gV6/6PLMYdjbM12nZ+ZN/uT4uoU0Rp5T3s26H2oma1a7azUXctZmXG4e1NhL
mDEAM0FYqK1gfQ3U3muBGxihChBFzAe++bDzTx+WAZTHwgQzX0gk6UKDMa5bgfpI6X2o1Omnrhu3
jfqv/OPde4EW3wF/6lDyXEatzwDaGTTbIhIPuA/9Et7OwTre7HGzJwWMbOZ7jywE4lANvQEkg3mu
hTpVLhgfzqqDBXTI8i7j9vAirg81Z8AyCzbky86dG7nwcSN3+J1bNDvzL28m1uilre73LNe7Cm6+
/F0CJ89i7I+13H4lCWMrJejBgY2E/99kxp5LUOjDUYuIU/DRHj5En4a/a86gPIzut2Fz+qC1ovej
DaIYCQokeWbaSG9eVllV5AvE5ZBh/O6ww3xRCHIS7F6JGgT43SCMDX26FHeTDda7s78SoQ/2VGoI
X88SC89YeV922mZS2QFA5rTj6ONqnXCEB+FQuJbMQtNEPA4B5jkBJ1MZ/58MTRy9I4ieFwnp2hEP
H5WTrLB/PtqfZlP0Q1vuZNz3i1GhUA28nDd5xb0hinE7f3FWgjW/d88PLcMLuHjWc6uh4Xn68ipU
NXio/GItHdjOTurCUQXW/6OAzgCQefo+7O4yKBbTZC8L4nyIaUD+OU93pxt+I0Clobs2f9RCeoLq
inw66kUQJz+NUF6pVovd7uxhWUKI778ENLA8leAe/tSU0WdHxEJIS2gSWU4dkIx48bVirbK5TD+2
yK/gaFfZ9uA24FuPa7siZBbz3xX4yHWM+CqR6N/faaNCNSYBrvHjmjZWa/7LCAI9w6n0w64C7ASC
9eqghbGc0rwBwYgMovEE0V2DXbHKm3IkRoXYNATgz92NjfdOf4QXqRgbTLtSx4iccjvMhpy70t7y
b33a7ybmLtkE756Mb4QAKywkkq8e8v63TKog/z/FJt+r4RI8IKszAPId3zXMfaYT9l+M4DcFntA3
LCm6vHXQC0ZNPEVzZkNeN6ITH8hzNcOzv8As1cigOQWDAxsCcHufcTEiGPBhiX/nE0sD/lhqowzO
zG0HK/dfJAumDhbZUwmr2qV6V5gfTDALhBsLwMnDBDfZ/Fdlcs1/7WURxia3QNA6d0GVyAJbJlGJ
o0zrqg05PqDb4Uk1AFpo9dZb+KgaIBjJdB4/NA/JVZJA0Ch2iWe1eRQ1HDWFeODAntsDB0qRnHgw
7nbB6YHv1bQmEBTetIn3qe8+MhAeag78tRjjZYKsYCDvlqVb1F+/iSWWA+fi87iEq6oXoBw/XX23
GccVHNrD7BmUY7LRFFrCnJtsyN9ONmsEJqByUW4OJlMhEiSeNCo+WibdvsbhwJOdriWn3WoQilS7
iDlMY1ICzzYQ8Aaa+22PLb3mPVCaberPV97vPA4/w6dIPl03ZNInZrNGqeIYBvGHo+Im9zA/Okjs
wj8kBR0Z9fUlUf2E4XakcRTW0TvC9LaJOJUaQ1vsP8KQbXUbzfKbTx3+t5pBrB/wA0zxZbRc2f3b
4vN5TcZrFTYlLp6kQ44TfUsBm6yXfclqodWwd6XARLMAa8/3joIJPkgTCXAldsVQkeYpv5y5y0Dz
RwhI+zAZ4yiMlKit6dHMNpGZon0FAn2CKA0DoYQ4jCJC3dqEJz89XfiUI8o65iXrID5Q9dGQfGx5
QuRB9XDHBFInE+25XGN7NWJwyLvu8PuJHTSwqIyEXraMmZ8BBiY/tbN/vCVtzUET8S4xIUMPxt3z
e65uaU6oVmYsiSgKnPvXxgVno/b1mKMqc0udHQ1dOZvp38C32XRp+80YKmPT9+h7D6+SLhFqw5ap
CCv/EIcu6zLNNYGDxCD6PyIFPC6+Ss1PMKb6KuYtnOp6fO9nS9hMM0hl3b3B83K4ZHmMhqa0j8Ck
480uu3gaSQeZLThMOB9gjjofUKqWEtqguunppnyOAghYEC9OoBrn/NGCwO8lVbmV1BmcdNI2Cu8j
1LtxJDFpJ6G7exfTpDO2YocgdfGpkuSV+GptuqFApPEpStgxyV+msGrxJb6OYvLRNfS9WMe+KN3P
0hhnS69YGSCAPHSZYV/XpiAmptAUHQONqfYCk7NzpVDs+qOw4c2GH4r/gHStF++zmU+vpA0NMT/Z
C/iV/yPmLxsuR/SaSjowMpBqOQO9Qt2e1G2kLNYn6Mk7dt5ORGr9zMecTyDbjQ4UmVYKloziEDYz
Phrvp5CxlymmbLkP6e89d+ofeDY+sOaw/gy+iMF7bn0hk1AmYiuMi9GnZ7C2+D47mjJSc/YoP+9Z
Ye/XRuRlQEwhbtDTxG24kDk59fEB3PaYgSnMh6/U8eEG6OqQk+VcyBf9paTan+Wjwd70kDCCf7Ea
+9IqOr81nckHgX8FpHWOzLg8eL10SV33VQ+c/q0rE+zgx+in0MTEiR7gDbw/d/8xc9RVgfVAh4/I
P3eAjpvKAmZ4vCCERQr6E78OgptSN74PZaPcSxHeGJCHu5RRVyQMISivsPRGRxkfLtM55Epfp2X3
jRymYnd/LPbxhe8cFy0XMkpzX81hfWjDGjHBIZzQMG8BQLCPzGAKElTd5WyepDAlLJsTbHDpDVg7
WuZeoFPVnW/Gr8Q0nAH/WWjPvej8lyB5HbVxS86vzwYwtvP5gZkWwU0vcj4eL7cEApYEpRCFkja9
gnPBOnj9Fj6V0gOHlav/Gb9KpxBA7v5Lyr10dSfQRi1XlpRvPyaZZHXtYD3EPh3JOedtcW1DaAuA
dqLJgoFU76Edq0rdKmAZh8nTPBbqwpqC02YGR8MjYSOtr3n5xOFFQCoHp3l3NavbJfhUzuf+zNyL
Bv2O1UR6IYIs/zKwVC9ad1u3voaV+iA5f0/RXo1rYiPoblCsCk1UlfvXsDtnrUtPyOH2m1XIBkrA
0LtemFmJD+sKIdSz4yX7lB14ynNgLY+wwOA+IMKhvuv17ZolnWs5LOSPbTTbPmtFDm5se/2FAi1a
KZ7NH91pb/CYWJWSBYPShbZY6PE0KewHNa6Mvm1TX8JsHi5YB/KT+Ymho4NO6ilDuJEXfAOeXVDU
HiqqepwMFxBsIpUR+4fndqYhJTBazYQjCQBI08CR/yW7CDsn9Dg0EtDXQVU4QW1RMR1eD/TKaGId
fL1Y2rpiZ36aC2wtO8OMaswfdy5WdasLnD3B8TPc6JjjIZJ3JLUVAIhXJV5GZ7r34D+CsiZEiz5L
5wUy4AGN7KRT+zf0lb5DgsF5mRKuIPTngUrJlA5x2O8c0tbTU9rGPqjv5qtq+INxDB+izRTAVZDH
2VcMQHb9vd7RZGgmtVysgz9TSSr1DaYyJboCQTfkypNq3g8InsZ0sjxOv2JPm7jXZ12tpoYLx8bB
6+Wyz4iuKDfCnZLlPkH3qkFoYpqcl4cerwJzrMYJCXUWAU+Xxcej/H4FY4/tb8QOUoZlPkJS1qNo
5N+NrSnEBTuqYVV9ReLQpAUK
`protect end_protected
