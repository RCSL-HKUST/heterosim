`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FHBj3Tv3BQCGb6cGB/O10CHZuyDxkgOYlE1RDKE52patO+SRwJE6sMr3Gpdc3WYaKBTCc5YzK0u2NVcY8QVcGQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OSgJqEVRt3g7ypst+jHjkMM7t3DG12/ZAqhGgo2b4WG/WquSQbm7YOW0T8GDuZg13UTWmzv5HoZcNvwIHcX1g+RAx2C9BEjoYAcDyY/RrqRQMB0JUL6pG939mwdp7BrgkDXhHWhGaj7/caHll9qhAWYT6En2qKoBB2+iEEP2i74=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FqogG00UODkRAUso87bZdymqz2eHJhXUROJCAzpfec6V4HKtkoyKJ6kgwaz/zGb9FLLVG20ifAusF6fDfy8yp51JQL4cHDj/RaR0ua/tRRme6NzIDmYMtQQCyuQgnxBP4JRmtwbhPTlg6noySuBAZk93PQvRvv92Kj1kysc0TFL2aahsiezQCFqTE+xwFTgYkZTnzHFOT/wDEaWOCBevM3N5NKSQX9p0KP+fbPU3jvfQ1NThOPIzLd1buCm8lIAjZcNQDbPy8EXIrKS7FvskAHTlUMJmtq2S0Ut2n6DUPiMO76uZrgSqxJBFPm2PzZRyGy6euH2R71lJLxGyAoXfBw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iPcYDll9d4ZdxkfPrOl5arRz93xn/AzL807ZQQtP9stEdSu+d62pJ3qexLoBNwl/ISa+87bAZsWgrWvlapR93EMSOfDE+kSl6XHHDYyAmQfYvq8zCL7LkCb6l9rghMsUhS2ttC1y3VmPwbgViHUUlWW6DlVQYqH4Cd8qerc9zNs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BwTYwARsoQ7OOqx4+kPptzGDZmssk0DoDbTZbVY/TWP9k4DhIXS0nxvMWx75bk6t1o7230ohTD9i2ZodaPFMrwc6OHE/39CUvuIHnWk2hxeBu/PuYaDI48sq2elzrRC+TPQw249eHKokNkP+IdvgDyLhhPR6zfqYsqQPYXlj7L25yk8L1upfhDn3zjoXdJHt9mxqjN+8mUkiG/idI9dAy6ex7nqgmpzG913YASdskMssfjULrTKCBn4Or0L1h/NiKXTxfNvEhxOeepqhJlIbT1UOvtS5WUqb3K4LFQPn/qStuQQvZB96cHO4D9sm+4pLMjj0BjcNBnxQj+eiRsjOVA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 27292)
`protect data_block
zMXvui3Iaunhqx7wGjMSiiWu/PzOyyNpvtYtE1xp7PhA5VTd8Jcvo/VQLBP/HhKe9BEEiYjKrW2z
J4Oez6QGGgN1gC7n9qAeYZ8p90Mn3pnANDwoMejGzATMrGlH6rqjgO0XA04GFSLtw6+Dvle4PsXN
XN2PlrFM134MBEiDn9/ilai7ivA+HnXtt093W5MpLOY+BHoCKyDy6MyBkSPbqZw6cxTPob8lXmHO
qhoPFtXLguM4VqbAEm5jkpNccR680K6rdBMk+QmGzu//PRuFLAMwQ/taBi8G4EgPEhmR/3Bl8SH8
AvIwhQEUvsMd+UZetYMy6EIUYgdku9Ji7sxnUhNSMS7w3vWWTaXWGeDBQl/p/ZnrqO0mhPBafM/G
k7QmFBi78gACOWNfyk1jUAOnTAa9OLzJb8AwAmt4+xpSSHh4gV9bsX/lv+03bmsch4sFCHH0o0tq
EsiZddzY1s1fMQZQtqR+fAq17oJmhm5W/w24NjVfjWBiw2KEB/QI/5QG7AamBGRP5G7h0dCYiTkE
ebi1lq39R6Gzsj69ZFco0qtKhMJ/3ShaEd39Mzl0MMkrd3/P0CBkIa96J1vge9J/Fg3SPzHDdGd5
qNITEPNEALDyJBguZYxmi0ixC1K0awAXCFit6qE265K1WxkmFxrBsWquRJl82TY5X7ZC8qeWXFun
FB8jkwtqzIS3+8d6Ei6slxiWBFA+vrmoOTwdGm129E5DZiVyQWWcC0cXSqVVd+X8WBgX2TKbd1W+
46PTK2keajJIlN2sMC/XwaS1rim8uK876HPX2TvebGlcYDCTiGcGV9TLH7hmCZhXvCZGt2O/Rtra
4qlwKrKfdl8i1m/KTmWs2P/QDdsR3KQHLv+kQm1CFczMhyxmzxNU5gyE50TS2GlSjTRgSdwdqJKw
Hlw5Ao3D28ki06ZOTBrtdQi0yUSUG32c9xp6HNDKXEdggCjCGM9OIYs7QiExIr7iO/F/xh9KrLTB
enKMQ/itGjCSHe8turoknrRMxPiNgTUThAafpvHJSDhndhlqwxl1zg2SXwcfeKLKKu2rA1e1r285
XhqbCgOfZIDc1YTw+jeBTxrxMbnf0pcMPkPei3KoREhHucFrj56USQ3mjAXe2rDR4AYx7OnDckXu
eyZwBumJGT8ueU0bPdHpgNH6VNLsb9lCbd96SuCHSvLLnSwKfY+ElBEtGfUJ2GdezgP6vKXs7ZcC
Yc7F1uU96p59Z21yD5fNw+izJEQWxZ6yEji6RFLJcsknRLwkD5C0YvuGHkky3nX/cb9PqPzv3wk8
My0pjXt5Go8BNdcJbtwFIEneG2oJAVelXwBFDbwdPUg0uKRQpeVWE97KWqOLJJ8afFsKeInFd7WX
KyMnJ70+Wy273OW3hBY5DOHOmsrqaBvDFwS3d6cv0uJ8hwGTWC+PKGkI4vSHtapM8cRO5xlpDWDl
wb3ekbQICCCDPgOegFNkOCj6rzc4jipkdJrY9q3JnN4jv/lkQsZg35nMukbL3mzHZ+f4XQuBZuEi
Ds5TDzGAEkQqQDvA/G9aJbAWUbJvAiTmhr2k9xEejXFJdyiwfvo9IlVRwJzgwTipi7mvjiN+0crf
9CPPNJ7j2XAEZ3PV1gsxNBj5xXul+Jpi/qZf74QLy7G26P0Xixjdd6uzgdgYpicCmY+9zVUpzNdK
FLu9v5rfAmFiPwlqbp3Fp7rcClMbFkgVUxwl+qu1tgwoJ/8Hhz+f6e8GvWK3CEQ1+CMS9H3h7PRl
3R+a/zXS4znUpYXNHkb89KEnc5IAwLgkAt6NIStuHP1uIT8crMKG3QkVNkiFsVtmei1zacaOfpCS
zrJ9USA8aaUj2VEiRCp8iNRTJFpKKc52KSidPtlePFRdtSQ6sPBHIezCocDlw/apuPw7ymrc00PN
ZXLwwpkhWVHT0lWCPMoDJ71aft4FM0ztFgdXAxRYjZXWOvTyycd/uBAV/lOmH1yXZzNknm3KFv0Y
sfEV63cPa9GLEh2HlDKIv6RnMuzd6JNtqL5DkXEDvYHcf+Gmf4Z2MA1F+X9UhYIO1jTPQI4Rkocd
C7Mn46FkOsQrOyB+1jXfmCoVLWyDBqeDLMTTSnJk5BOYZA3yVcpqdKNXyvzwVSBibQLCTQMlqMaQ
Tjd7/G4gTnh491ImHzQemI4ewpfxggd8Khk2vw90SBgl9/xchha4b5zJrovbQ2jhfMPRDpfBb05C
2AkMAsZaOMV2/HinCVn1UfwsPnBKpwGWnhA0FsFowPGAr8uqTQ73NW1lxJqbI503JdPhM92PGS/o
u6qefXOadnVveXkvGX6tGZ3yJP/MDz3o3bB8kB4l6EBQVppbI82CZC+/szHVkLqFfjblfcNUgMGr
KFUQeS1zGRoBD8FZ51ifDGdhriSj9sGwiXW48yuno3R7aSTOPHW2CR1xPrZxjaSKI65hjnL4HRiN
xu1xe7Z6YK/AdqY84uKO4si0qoaY/zpDnImPhNIh6/HmOqxi5EhFbQhlb+KQqNVGWftRNLgoOIcy
vHth5wMq9I4dkmVebjwfI0FnGTcUSeJEG/rpXX108EJAPmGtZQXTzarCS0s8IkgG1fEG9Nh5pP/6
f9XSHsan5yhlfTCVDbRT9eIN8gwsw5tncEIWxrZTebvwmUmxNv5i1u91Nsj1HiQR/GhQdJH13PdY
VXZ7nPtcD9uA8VaMQ6P3jLX2jqigG+hoZyS6s2+AWwOz6miE+IZOG79kKr+5p/ov7URt3Uu64Frv
UkRF56ahf8T806FGJUhXDtz3eLuc910T2gFK2fD6kkdjrIAkChUwGLm6E/pQgycDJaoY5BuEGAIq
yq4azKQoJz/qce4RUmsxLhBxXFJo8C1CxOQxcWrOgrpJ6N+rQWwe3ms7sbYXWQlN2/xLfVzRcdhu
EbR7CitOoQL7lKX7oJi76tupZq3XRYHMqqOSnOGBmdcsNpu8BrvMaQZOvoni/rxl7AoYlaUZ28gF
+YFfEXYJzwAxNrNKHLBqbHhKv/T0y7BVvLroJTGbzlV5E6YfeMSwdUxmbk341qUipDdE7HB+GZdE
144sOJoMCufw8xspKpCT98eP9an4dkxmDDsFrdPPDCvtnXKhmS8ghNm/cGphmRpS7hbCVOM7WLfY
sPox45MXeqI2BjnrKC7tH9uyoj+2OrDiZkcma4qMjEv1j3gBHhxgoJh+BvXCKd9Mrgl6ijGv2GfD
MXuLQMnBfPbHKvDpY5DtHzUyFrcIGQiSmHQ3zxOspLECfYWAwyRSnmih/eiWJy0lR9NaI6oXEb8I
XZtZFXvY5EVO29ewF/37i5wu12ets4PckBOhnNA+6mds67ZYIfCARKiA/KmS77LvA0D4qA+Nx8YP
ZM9pbAppfMjSHoTkIZR6lg+TjmD6EDa2fiHlqa8qQ8ca85CJeUzUrkDrbw45ItzOm1ItcU4TOy8V
WfW7xzeC1oaS0UBY48YF1rDUdw97OgxmVIhUYX4DcNt/Lve2ysnQlhOCXc1rv3+FgSfggHpqxmxP
5fh85Bz8ULsc8DmoidziPVRIL8XFEjGL4KHxMje/s+yvEq5arMQqlhSHfYX9woV329r1YGSTdtDs
dAaZ25LCF0kasOEE1vvjqTZW2h0lk7HTJAmiMpsblxDf6a4If3hi+PKJb8vgFXajve2ym6Gh7zYW
gaaUbPvukQ717DkmECiob78CVDOgF7YA1vvxIVbHGwSyC6k8v32ElqsD7OXwDUwKr+rBZPHcFy2r
LI8GgYBsDtlm74tJed23u/aTqTFcJOkX9Rx0ZatCPfCicrnh5p00LeNhiuO4pdPx7YEhBxG/vFDh
Q6ykprcN0BcceKC+v0AXQ63XQOhVrHhmwIBQrQq9CfKHIrzv8Jc8k1c+yw8NZLJXMXQfQ+4ISE/M
fOaI/9ZC2hovUVeXm8DvQWuI2x8ZNGizAXtZeX8ku2Ymhkr3nqDuv7lE5gZDTHhXcW0j6KwGSh6M
EYZVB4VWhs8R0Wdl3pk2GAg3h7uBqXTCDXXW4vkkyalUAh0+oKgaCV61MRW4QsWfAE+GHdREO+xJ
+sDkY5P0df/Xq33LHz5hmkm5zlcPWEPWsANFrsFuVzFxd3+v05ARu6Jost3Xozeq7XnmyNGn1Yxe
bugayOb00AcHIgXX8QBP4uF5HrkdvzeeFlg7FNwUshy6Jwe7IBBsI/Vq0/n4FIYbmpTyp+HCg/rH
Esjohxy8bdAR4+Mcnv84ZTOMI+0rWU9WZ/eMXtGh4WXqJtjL4/jMu0Gd3AmDtIQOIEq5+v0xto3Q
1wXPFXmytVpPcv40U4j1hdjatvOU0gAfndvZc221knrDmpSPIkZNhMFI3exH5Lxs3o417B9JvgVm
+1+HS5uu9xlH0poMhGo3/mi0NoxIyLs95GKp65o9pqXqKusN560B/lGUbT1m/S3o4HNB+9YtRrnU
yrX4sL2qJh4VQi1VurDG+zCtPmYCPLUymwPIdISYL+wbfUXXsA8wFFM81c3Om6BTV4G/KgSUCswL
R+koigtAc0KYtFmbQuHZjn0cuxdAIMz2yC3RDueJqNlmenJB/3QnA8wzkok2PQpJWjjf/kuM1WuG
E2YuHm0zfVoagWLAbXNOGrWefoJ7ZOKyqfvgRzcNYMUesy3GmT0iTVda+a4CP6g1mEUnH3xKcArT
3qELQ2IvqJOk1UpGyLcaFjQSwpwJYD/qno6s9Dl7XWfdKh1KKQyrG6jEg6sXoyLXK3kIYu0bCaUY
hItu8QkCviA6kkgW/lBx5Vp1GBsxpYpiA8OXZ3WZQcisuutDO5/1v4tqBcKjWdGwLbI6u4E7RsS/
xEZgSI4uW9meSepjDtBgDMUeHXmMV4kzN98mz/QaOx65u5xFzFE/a/blBlP8rjhFGI/B1E51e/nq
2umCbdl9e0V9VJCN34NhZSK9UYtTiQbQuAO54hAvuqxHNRRYPNkJmaxdeAuKyCiLka+prnqaOY5B
CrHhWfwojclEUKBcmt1WnhExwflf5nBrxoIzNMXKpYmDF5x24NUUrTHSnmS0+BKfxUI1Q1WXEM9P
YIrHDmTqhQgJP4IIozpGrIMgPMqnr6qEvXa2ghZJWmjEDE2cgXm2kGy4E8nBhP469T7MiKmjNPme
ezoV7mUUddNe0PpjmozpSuneF13ORsSJneTYlq8pkbho9dWTOp/CVLG8ZVyt4u3xA6LNS9B0RXqy
3CAj+yW4zQThwTe6i+mMiDOisWaodCEbkICVzdUk8PYqBAWOCF6qRP3/JwDHK1DCKxTU/rlf1U5c
Coawlh6p1Pb2j/V67yOMr/+nvOM1a+RE1eHEvxDSg9gs53h14FlQLN5gbuOIkho8B1xmn1dVvJw6
hFQkjH6ICWk8tHTGEwEtBjT0a9UfkDXvAqxzh22YGzZT4N6OPT1oJOGUyVRLDpCX9DtH8bqXeSTq
d0iWb3J/px1WrBjA80CE8ryWhWwaY3jKAab75aSH3/EXHIMAlocs/nA+lczS/jAZA1VmWgAhs8Nt
jRuLoStVskmhT6WLANPmxl+76b95HabG5IN57FUTKuFRr9gsLHaJFgu9vasovM6pam/B0OrSFFg7
HvJTFvXR+I38E1BUjvOH8JhQa1wcAhmPmjnxUm7J4oQ9CzOgm1sr1xKY6pybVSxBPE+CMlNcTuhk
/R0nLcLW/PXsdMsQccOyklFoV01CwkkzPVPXNqxeR14b13vToru0zXcsPTUah2esM0f5GHlYDRzp
3aKC5rgEABpMZnaTSJzl6fG8NcnB7CjqFHW+DiIcDNJXV0aWFkqA0H1lW9SHECy4yjxQrYjsD+ZB
B+GAQPwAimj1mYgIY/MgqbW18JMaGSVMcayJkhK/UbGR6COgOQk86LpyUwT2TU7P/p+HZw+iaS1I
Gh6SCAGxYZq/FoY1da4iTByjak+2cGDF2nDgolM7IfyM/+WP1MuAyBFqvnFQHtTU8FP16SMw6/XH
AWlu/lcefJZvvczm18GilVC6eFoygvrVTx0NiPCjB347qnbm6YPlLRnIuePKOsXk7+sirDikyp/j
/ze5Xg84jpIQmExpsTu4h3lxgq2SzrecUUeKmr/2xl6mD6FRCs1CzuqtURnbs/JZzVjQYZgIEmjk
AxfTpWoLmAYN2DIvl3zf54BLFZPMyQ6KwNag72TPhPZh3koImCW4Otu3IW3RTyeBK1+Ecw7FRho5
L/xFyloAsiZer0Aas3UzIinIZ9uhJVwGDSkyACTJVqDiAZD2JZLVSrhNrQMRofmECYFhQ4XTbTWj
LQVvqcJ4mCySaG1DUnFYf+pt9M1COqQauKfPYwnGuhSzwO1yBOgq1zgPKs1R+9rXO2JAvNJEG03e
JBv1QO4OiQ4/2i/3dYk85GnVxljs0pSIJprp6pmFALYkfhSddAYMxgxdpQt3GT3+5Hu2mXwdFbLK
O6iuguoDN0SDOVA3+gzZHjt91BDzu3BQuYmyiL7mjm4Mt7ASrO/PQrQIBjD3PQ/BCYtDuA6ie3jr
96vPmjL4vIMXaXjIxY+svGkb0NoOnloz5mXPJmonAzCMOWess9CeC1m5q0YncJc7a509vohdwnJt
FWxpq9E8FzbAW3OMbUvIOVmvIiCwJvvFJnmNGPb82bCuXYZzpzyNwO3SKUNwgeoCk+0HGLw4gm4p
HdjoyrA2LazK3BFQ8Zzvff7wgXnPGY2Hrl5lKJqp+/vYHksg4CVk8YxFUVMnS7BivEEOfq14IaaJ
XG3sKciqSzkX+Koclf4CI2VjE+b2m674zqw/ZhmQxLNSzT9AMAo5eqx229JufjlbOVw9XfTk4ZZn
Ik3KQnow9TYk7d2H6BFR/+agqmWKs9j/pYwQqXtErzNO3fxtYD4vSdNzt8sVXgSJSiqHmAgceeH9
gTjlBfbhY582h7nRSIzE4s9ktCKnAgbJnlFVWQgmoO5v4gwrGZfSNebwTqWPZDrzCE8Mh+R6fhU6
gWIWQUHWMtdYSqRgzupkfAPJO9gwB0xW+j9CrFop0FzMu9Zk5pLqD48Z0EKzSIWj+nPxD5o1sfkM
JbGoHk+gAtkes4saATxaza98WriJQHxmOsn29yD8R1xya2p32s1WTj1Oqd0H0RmAbEXRMVWXIIir
g+zzGBhmAWIpfrkm2x1cETMktQ0AlAAkFaWN0e4tXKW3c89+FE8RKoLZGFg/9pmo/Xceb6EmUiQn
7pthPrLeL34jFLGeCVp6crWqyf7fybnwCZ+qx1GOFXpMFYqDwMaJoCXa9MQR6jbwIE+w7t0WW90X
BXOY0bEkRaMSLeTqbqmNahxzP0kVa+C1YU+PAl3iWEe1U2QESpEMhmxSBcyAB9UVnJuIhFqlVYyA
D7afcn8SxGvX38yb3HdUzzrcuqJr0g+wEpI6twST+kqA25TqNAEtBZ5lVGUVFtpGG4CjeP8vU0WG
aJ5EQSqV1UEobwIBF54XDsOj1LcIrT+bk+DKuVY0np1pO7TnCeFoNp44qFyCbJ09OXOE9HcTf6ZS
51aKTwsq6+0tj1gcK33ylHF06A6LpWIeqZhaO98MlihEDb9R+cxzTu5wKObQM74FclfUUq2eGeSv
5bq8dUfu6OhPBr0oM1/BawUytBICT99SdESKTjCmZspzoHit6gcbjy00rlYV82K+nfi+Vrt6zW0n
H1FfOE/hCj2EyNOZZKDePH+BafA210EJl6BwtvpfQnKUXPqTxtVY2R4ps0HlNuGRNUTxl+3FhgpK
kPz4fhw6bjQcYUm6BIwuioq1C5emJqUK4NodZ523L9+cVak4vX4Z+GsZAJRHVnMytYlxC/PKsNf5
6PKaKrDhjoBb2jzNpfTjqcGcRlfWFMfmPPz6ShH24fpUATsTtpbh05FDTM7LwTpwsJehJnbSuhek
IYiAXjKVpParifRCGzt1qjZj7ILy4thJwJXQuW9q7AiryoGmu8FzglqkIWQOLz/YjW8NxsI4LKyv
fr1091IwXgP+uy6LkIOKxsbggIyWiZkpnEyYRuPEzje+hQ1ax/W/9HqHRyquca5n1A+jUdIMmOvS
n5hz6Hw2IAWh6xD9KOih7j9XdZDJGxIs2KDpBaVRczwUhY4gmCgWyENC6Kk/TLohwshal0pFplaR
Gm1xZu+IXMDqq2aHJp8dvxCVNlIuUqSPdLwTSSUdkKeZ+JjVnxjopkAh1+I0gJpT/oM8/8kutzqq
WcVMWkGYV/KCJl9YpHq6Iv+FFjeLvTh0Lc9PZx0J598l5Dz0+RjrAFsxqjTNPrplog4YgZBb53r1
9Un9T4yLdwDw4pnDPLp+Y6YHnx1hgl7ebr3kpCldnWtftzTMVxc/1qzuTSdSr8w70isi8I2B5dYG
DEK/nPUvaAoWnM+kT4ryXYZSQ6ogK5cgxQX/j9ZeaGJOxtaPo1ahbEvdszn8s6PxQZjMT9MvGeVk
vY8eLXhvmOMBA49O+9jN+5ZHbeoW+ZofsEJMTBr4zey77pfDcxNNab37KjrFCegb0xixUgjeZSNr
vJsDh9sXVnzfuwzgRFw8mEeppwleIbvT0EGaRub6X5yC2FsIOxw1HzV/Mmn1afRvR7WQEsluKS49
ok1lJ7qgKnU4A5tvLL0Fh12TiPVJx6XsSvAhGV0kZtfc7zI2WeBmlDU5NAtA7cSjXG0tKx4Mn8do
y3Tcm+SxajWgN0K6CIL7Nq75FUu1kB3Xss5u09s+tNMWAZo6giZMOIOTx7cDaEhM5zrJ7Lh0pIrL
nKOZIBYoTFeMSotP3BlapiWdhv6kzkMArpItGglgXBDX++OIaiOCTU/HAOorcSJA2mtHHN7hRbyW
X8FfihwecLfYK9/Gr82mz7RGo4XB9KswTsh4iuSn0j9iG8ffRinBH28Vzq1RdowWZG1DPIiPJmUf
5s7PVXOsjniVljw/v1YQeg905QcL7swURH38AspgFdZbg1WJ3RIv9tTIPlqaB6fGLi0UEqHJAguP
itsoE1v+h4ULJCahXQsEcq+HI76A9vOEM5Fe/yKUbZmFn2LpaRFWkuFbaHWwCVLLIf7xBggVjjI0
b6Q8lORzvq9QEHfXAvuH+aEYwxvJtv/lc8HzTWO44HinFe4xBOYP7/crbJas4NxDYEh8Fam8gevg
gbuoQMhZpgSd+9h9a61QARENtK6WEwW6LZekjg9gHcAtyfR966lDodMytkT66RE8/NnQEWkmlRUp
ncxWObbh2nZS1ehU3Z8Ulb794ZMdcXUtZdQVNgn/5d4q9/NO5V9jiLF0LJYpDD59cUQaS+wGFOud
Dtr2ePmc2mfg7Fng2aYhASzsG/4hO3qEzY6VmMhhJQFTzqAHfOzNRblfHJY09NbrocmZ7nYPYv7X
Zt2lw1ZHvZ3g7qBGS8FXVIvy8y43MkGgNrE6XJBlTPsZSluiXl8rBGqFg4ocPxANUE5Qwr7U6yFs
qB+qJzlX4lxNokKx7PzascCXMTYwzSKlgCexXv95n3MzB6j5r4MBBwSDYDKQL4lvDD95SessII7B
LnPDIKQ1wAoK02g8poLUo+/hlCJaq3cGXX+3ypaVEQYBkLgJP6JOtA375KIS4jlv27KwDCR6zIyb
5pB5osnks8B40zZqWiku3VtmhcJuykoKl97OgyxndYCm9JbGuOG2M1OfJpRR7A+b2pMXikEpMxth
XfezCfZ7hJqjLHfCgxjpA1FegEXGT7e3qqnIQ53/5lILDyOpLO4r9c46URc8HuNNJ/ZZcLk1JaCc
Bn7B1lx+GMJNW90IbMZU1u4NJh7WGMsZQp8mQ6bUD90ZwMAIgKg8Hj2JZcxfctUXznEqEVOoS/h4
pIBmj4QKlWXUZw4bo+2TlTblzVeZgOBgXE+HZJ2pXD1PyAbVtTG7uX+GTEJYp6jip2kGAD/VQgrf
QRY8NtbyX3AxLaQCgWAGE+30i4WYS3dk4rA7/GkXwjKWzuGixoa/K+bFRs7i5RE6QqQ0o2cvMzW3
kk6ILA3dvgH+AZDUglwCyNNwb0T1Hokl1EB8bAbwEMpEqTp3hz43YD8FDnzXJFyd86hOlxzqkzB3
EGHYPG81d5DkVnEssM5Z9XFfD2uuBusR0Y9r2G+fc/p+L4U5dIdNDug8Pw1d0HHY/AnTb/bteSCN
ueRH8iVhCpa2eTKLy3pkwcHkIHWRlvbC/dSQPUfbJHJOsIXvkbvHJ/2Mpms6Aynj9ESNbNijBHYk
R0QeiKTrdCvkYTTLfXqzUY6SGnkqQsSu1zenBljCcSpcm4/JtIV0AqGO/ru79yGAdYpZ3wG+35qQ
+Og4CmVPQBXVJsrWhsanyE8NICHx8HDDfc0Xf7qE3jaWYBPiqshCp7DskOKlBNymfNU4U699lZsI
EAX0Ds4r3eUrAIC2ns6Q0U6xDRJBYzu6LwyNzG0f9wJnB6/u8zN15+TJ7dK91Fis0xHKiLs9EvDI
qohhNFoch7d5tnYhv7JfpUxMV3rPjmWXnmCSabwbaGA5ymBfPJ+kPs+u/9Ka64Ht/PFdc2gyVe0y
vV4GNArPr22ef1R3aMUJvgdmH6Ynm6dwZu2hedUARpynO3B8pXhZ1yr9eq75WALM6K/A6LpOkG8/
P47xw8gQEXKoud1SUY+2ayyYXHR6qyRBMtSYMKE8sFpmavZX+IX6PQOBSSCMo2HX7erqVtG26dwd
lRaxiVr3xgIiyNjEbCIlZbdlWq2n3MAcsrNxObinxJJIAxiUvb3+YVH5ITXdPVSnDniQRcKmDea1
U6HMJHfi4j56EshgkfMa33YmeX3ftV9XSkjKtSZQRD+3QbNMWqOsuQhOf8De5uDlwm8yDRSKYXIM
mzij8EPMAYyvW5a5hWLAcc859NFVBXFGHm+KsKVg3hNcWJHfzOpow9BlxDIcWvAu6ABzwS3zpDv4
KXSSoQMNrxOzNK0kqytwmapGou6eFCqfV/GvASj/IBSumyrNbaDu8hWvd05sOl9n64lyj8UhoZJ4
WDQismNGK15+/cftQEV7n8EOZoco0yl7f73Kx8HNhdQYSxL6x5APxFqXNalmvlywSFXedQGgUPWk
B3oWFRbYZfqCygDQPPPuys/JrSLm1kY2i1NYHJA4/B72VXpCUuLQ3nfQtU3bFhGtccAxzDIAlvrn
SxMWMl1GIQRo9lSOEH/dhoMZcEJegUd1cKjIdV9Ndhn16HblqVw6345A5Y2nenGu36zT/XYnvY0S
8naZXBZEbKFhzPVb2nw8YhdcVTAFQ2B9HMq7b7PDEJIrTA6T5p2LSZn0kfynMG8YjdMCThrrEj3s
jL+z3amv7Ii3BH4/SZ6l4Rdz2n8PnISSfgCiGzKZcTi6kSksn73vx8wHm8e7d2rRvq2Jt62hb2Z3
NkHI6xZDD2SJYUrPgE9GkNJa+IVQboVWFCWITtV0MrG+p9xfou+NldGLMVuESt6fAG6P1f8FXBn8
E0epq3kO4U16Yxr+HGxD/oIVlH2x8k3NT9iZS5gYKC2Wp8ikFwbtfOwWvefYy3NxuIeWdPqxSGIA
GJteOYifXZtanLYUv8CabduOImzCbj/i9HpjC58BrjTTaGBVe1GqTa68uzKJYmRrg/nm4YflFrZr
EMFXlKXMP89IEkErppE5NMPtRzlLSbkEXeLzB46Mmk6i4dBNtmR85FfTAE2l4zlE67IUJ40raz+B
fEj4Buwz5Ggbegimo3Q7T4wRJqPTAGBtFRZjUZs/bO5cs4ANF+QKDfR5lh3ouS46MRiTrl6oUsRI
AYLADQZhcdTpNy5A78g9RgJfzXNQcxMxEpbVHVcbJmx6yd3r1+lJ1XE4liAby1Vu90/y4ETrGNdV
+33aNVtgWcfLAfnmClUG1mkhjOiuAIqetbIrUcLMlINGH3H2tnLkfOwAt1i1EPpboCxBMw/y/VnW
lZZjoHbqczj/oTKgLCeja1DIYB3xWc/HcJiNRXKxDaf/kC5mTXYVhIPskTSbwy4OxQqHAmmba5Jv
zzBisT3BRdI8I6KeDCCrCo/bdz2WroT525eKdQN+r7sGUPP+HO/2QtQRaDWXnyaLSe72wTilh97T
dzrC7OuABVVtzxSraqaAJV+yq6H8rP6m9FuDjC2Us/svckhw6yGkYXb8bXAiL3wh/vL22cHRtcV1
TqJbZYRb5LykPeaLmXnrEv3jpgAvD4z44Kc2foIW5sDOeC/HVfmk8MOg8IeFlohxvpF5SOJIZFMO
j/Or/q/HRu7Uk5xRR/J3TUcAGYeLzhky5ySVLt59TSUwKiBPIBLWIxcw7I7ovZS9w9tIlTQKAJIq
IlKoz9/BYAMinzlsX3hW8bYF+/2RLNFvlqeS4bEcF8i52bOsqBkRUBwDNEOYfnQsDoGozWqLNK1S
ZfTtJ47fhoB+WMrnKJI/7ZzwlNukV+ZTgbU4FMF5FgY03SyIDTLnTD7j9CrBql/gN6u7l3jjVhek
vWrD/cSd4ZqEU4cP8+/W/bgSbkqbdDQcH2nqFTChlHamPSGRT3wKs2QWnisnqutLucR7QziziHO+
UcnsOkJ7af6KeuJwFsRLXAdKRYlukFns6xx/jPq4IbPmUXo6oKsGaFqYpuZaubVUSO4xFma7rv+A
PYmKs08rnSTBw9vC7NBUYemICf5NGCgFw5j2vLhGmqo1hqj35nvdeZs+lvk94kE+UIgN3R8DreAO
e9BNPBjnF49kGkFz2dhy5AU5AoDeVxVyO7i94Bc4sMlQ32dO7B3e5i+nqA7f54JCMsNrgusG+8Xk
YkE2Pj/UCQFdhcoeti39E4DtE2nV/KWT/CAS7rgYtKQzC6tvqQVHdydVHTYb4l8lJCjUITmY7HMX
oB0qakTMKme3RhZZczG3UqCJVarQQD17u/qHBY2+EfVGOf4djQ9zUi5mF1Ws2S9UFmzRELvj2D0w
G1A+r6yJjkYaTfvxSwYVVWu8R2E5REEQ/lBjwMm0ly1jIuwHCJfGpl38QNmEn96XAjisnnFSlE89
/kgpn3EoIRHjhuW3vz5OZrDaUNBzpROMeGSR0HNqp93VMSJvo5PJxyd+SqLK3SC74RPQz1gif59C
nmd9ZtmG0LALwXarEjtYGEtlRPGAL53mQ/RvVn8BNddggkKr3MQ2bSybRcu5wxdrwe7P0/18Dve9
d71ZCqBllzb6Vb8byRKiyQHkGZdcb5//Xuv0DKpGs6nUZLGWCR+3UWqL6M4r+epmAFXRDQZLufN/
zsL84HmyT8oLboHbaJcsNyewsNg2mYq5IqXza46iFIq3LieQfpDegNg8fOQeRo00RMRLFSIymJnp
9IrZx694WHmeJXY3ijAYX6wUk8rQW1wj0X3Ij26XtsejeqgrdRT/7Dz5FmuSsB1KZ97w7QbjjZ/E
HQC9ORFDjp/T76xOk4cwrHlsnIo6kpmp03kDi9iQaBch5jip7OYYpxAJE25hQSbx4MJG99rGJ1hK
BJSunbD/kXA+m6zKZ57xnWH9Q5eO/Mkhlds5w+EzmjYUZ7L1ORL0jokVz9BYw0RJx/ylnNYr+DIj
tzjw0yokF3pE4ZWARh6xqSJP2wg3Uzct9h9/dLyp7gjV2jJcRTExc0fQAKKMKegdtKjZ1vjTpTUX
2TUsI/4Bik63ngK1BM48J0wbAe7B0uItK71trtiYCZvDt4L2OF+BiMDoQ8sMZa+vrCMFio1mqPuJ
+2mKzC+ABENSm8YdsIcBN/tauuAaXvScTkDwzt6PNsAlz2C5VZ5R2gskgNmdLQpVvkbwcYashG/X
awqv3yWNYbpCas24rpp1zPXd8wj2uA1l5PjX9RtMTf6g/wX3/QTuXGV3Yrw4b8+QseXWxDOKkAxf
zocU4gj+EJcjhQIfVF/83dnhaPNb+JRKTBvzj3z7wX9ZxctmqdMkevHi62m8v7k+XHJMGttqk7h8
u7Tf3F9naekjWhJR3gH+ClMQncoIqnyAzS3DswJMnDy6oPpcMnj1y3TAUp5vUQQNZ1/Bb0rSi57X
ui0Li6mr+BgsTiUjh9Yh4/UzIxurnV45TCyEvZ7umoDzpwQwRL+EkKhZqut9se2zyixg9ZSn3C+n
Fu8LzreZMpDbtkO6UOp/5MbjJgo2eHspywvLVpyOcEgGMytGlPNFTPWB47vjFpJ2N4JNoc615u1f
UJuwzKdNB24XKpIRN5mHVJ9vcyZtpHFqen+5diSTErnVTkhe0VM2fff3QmAk36oC4EAT5mW32uqb
2TQBuVqiV8QcC1u/D9NpRpRufhYcJVZrVC1DNCgfJ361kXxrRhdRv9zEjhFM0JFrRbDASkaZsqOK
0x4NKecvFxggGvdUoRUAWa6i86LyFRdOK3y803RVTMBXeTP8OugNIyWfxM4M5rofPiNEifqKrBRT
BuRSvB+kaZ2dKc8IMiSFJyubOOypRiCyQ6Vvx721AtloojLhqgfJ6ml7GjwK8UBsCIhZl6QZ3ya9
1pT6K2rWnLjLK83PI1870UuxBG03IGU48mQtdmVG915uugkJ+3pqiICKo1L3U2PMS6285yoxJJPf
XZ8ktSk/DrLGJbV8G7h3KyzngeXPflZWdKsk2ibRnHwVG001ZwwMXXteJVC2MFkTlQDy6yCskANq
0PPJ1aqOwXm97o8TF+YA7AbHyLH0IkUM5MvNkLWwJ9VCon7iZOhWLrkScxOsT0NGu4TzdxtjXtak
Tbu27yRyE8jtDKoXW9V7ZbKTz5bww/VqIxUxM8tndp/xtzgr54ptQG4fLycHMhMasW9jUQxVJFSv
mVsZN1GluYgtbuuOXRRqOZ0gaXSFDuc/7sdY09QYedNp7mKVGf7i2BhltFcXl4VQ8UYZWWb8c3AO
j34OBV4qaX6jlfO0fDsnAA6LbwGotgGidsALh+DsQvoXzvMipXe8Djtwa4TlkAV9ktBl3/3rq4NN
KwrWKCdzvJPSLLx1PumQs5INs2rkLt0ZXWenPaClGu2DWQQhAf0Dj5DH2Vu1ftXUT5TYrLECer/M
+rzd6b7jLSLn96zwOKfUsqO0Mcaa/LOeoJTbAyQN7f/Vh+FShSBFjG+KYUD2GnlzxFVmFWhvh36r
F1qqM+FFGbzr/4fluc2/5591pCo12ZwhnFRvh9KuTmt6MupdAIV5HsrcseTWLBhW/Oj3lUSNT+Sv
cwhlxfdBA9SNIXewzGA8u3VcE8jC2c958drfPnitg6JFJltvDDMMherJjDKh6XClKIhz23XzUwwf
09bIMyHf1ftYXufQR53X7pWjx+hJqSwfFCsb2wrj8q6S1VM5CT6V7yyMuHnr6fj+97mQZCgOb2Wi
QgLtF75JMufEzvJK4YlcNnIpeS7lwo28oOVZ8UC/DFpyyCWe4RmbqW4oEtOMmsxMzS7szh/W4AzB
KyH9WHJEJeMjWcyvuny+d26IoygdcBku97wo9W9Z46lubbvLkTKw7JmyVRaP/40eF+5KTV/or+KW
P0wm3wiF0ajcEJPpTJealdaTAJQ/JjdjsvMbfvT47wvwvEVPKWJNZMq15xT2p/Xt5ZWlfcJxA8hz
0gK2pKwhvpWo3JyCqznAb5HDEJJLIZ9BADE3THPZ1WTJG7gzH7xcLB1jfHKwQtGX39Cyu7XOkn//
kk0GUH39hLRthT51izLCEDARS81eh/tqJXBiUrywEiCzCRmelx555dnRBJjWS2m+binLienF3ZPZ
oq0j7WHo7dN+AzfW0hpUlsKA6fvfjAVMUtFUTix1i1ClTK3fEsKmzUuHdfPWPhyK3R21MD+xYhXy
RTCgdx0Atv8SgaET2RLGVKXZ6TlGVUrRh7k5Jtif2dbwbbWLlJHmoKwTrk2bwuIRofG6AmoniVmy
d+fdwSyHQVY0QA+Gt9Qua2/9+YMhLAUaWgD+lTIO7T3IZ8XUQtZWAIx7RgHTg+VlstgtBZ2QMF75
w3bIVkGNAlCP/zlmCENDlMS9AIfrcsm5j++xu2+hLDQXXRc1jYJdI+2Q3P1mR4/9zsNUZJu09adj
J5szgSf5w+pmP5Tno1ziz1M8LUyLnkFXedk8duTjYXCrnklNsAPY/AVe8eLpnYiyKZQGfwSchjue
tFQc0VfqO6qRhNlF/lOyUlQ9vCmUC83P/0+0TIILKPbREiis6M+ZQP+LbcpRjnXV7DKBEiMvjX7Z
jZ/j2nPJBCVC7S67MTsU10DxULFAIMK5vYC5kfAv9MJGrUrEIK+5CEcJcxEhuULpB6m/EKw9VDh4
OybmIV62ih0HQ1YKu2r2otC8grFYhe+mmICMA3+9s5Y8S975AhcNf0W2RLDNAUfOjwlX0/4pbI6r
b3U/hE1MGCNAik5r/7gb6Qmgqf33uFXidSfljljqf1IWNIr59rN6kauJdaGCexmBUUM0619nMItc
wPnGdSord5LZwwfuv9HQtKUS9gL069EQT97SdqeacKcCYnZ6xqAESzUC51bv6VG3SwcWjP91JDXD
ciwqAWkJOMhD+TIdfp+GVZ+uaE/yAr3ya0H0NV1cRx/sdEC8N5aKj5KlDzseDHKNRO+/GXsmYpSm
aIksEKATMM+ssc0P07l8CmKdM+dvaks0Ydph1IC6mC7+GU92QccGR8Tu1g6Q2TAbuzFtSqxG9Fhh
8g6e5G/u42YLvaCmHN9i6aWgtEbCIU5vdIJP3IcJk4aCo2M41Sb0T5cLiWnOGOK6CCLfapqAZtmN
FGGfXHReQt+Mew411GomUxwjnLWtWeXyyJp0rM9hn6zJAACQFQUdUhooHLYrRC1OyQM+5POfN0Rd
F2QhXpswrPyklXZ7mq0sXMhNClsz263o5rTp4wSOmD2DhXjJY4yiQYdkTcRGDXAOFXwqCIYGNPbt
iM7F+in0Z6XRxnxBx7EXAtHciDYN73CiqtbNuZ7HlQK9KJVVsGwIzI8YTPmOPkc7vGwVYMniGFTD
6wm0SUHYvPe27mOTY1ZF7p+jRy3+CHxJfbSYS5YXjQf3n1wxcCOjzLwNQUu1pghUUDS7pFtbuslU
LIo1gDunK0HmSJql8juaJN7kYBv1FSvRg+Ex8BzdmJWdxZxxxbwi35irxKqvvDCX2J9zY4t9eROB
JU3fI8Kg2F7tyB/E/s88xu6K2LXDxgrb7AHrST/oC7/CgPThag+IVt6zGAC5cWt3M5JQ5GqdZ0BZ
cHUZKvkjq7Vx/25WXz9TThXjn/DayVKQPyWG7z4f47NA2oBTi+MPR8WaDJkDpVzHHo9YtALAYllj
xxHOcCaudXcDN+hQva+wDWAHWpl4d0hjPKzt57XYCRruQ6CLGvgDzTrUSBdr/+4XIfC8n3ux3p0b
tX/kC2VfAJloVSqopjjZktnFcVjhj7h5TEBaN/b/Pqlu2J0h15m0FZU/39T8Q37dR9ktoI2KMNYW
EIsUx1OZGLR2dyxHpH+Fm49WXruVgDNHdCTd2UK305uI4m+BMkfdaDB1egj4nbAX3xokWgwKwcqi
7v2MaWP4kOnjudi61Oqu85pvosp12MQP5SidRADhEEsPjvuSdmR8Nb2bZQONMYQhZfqaYbt0MMVl
/G6onR8EYK1Zyy4cyATn/+AGcX3YYrdOebeIz0sriv89+psT2YR6t18Vovs4JNAoasLyG+T4n0yc
oRGfRKTaDFmN6ranYll9TxTLL0QvRAQ5RoWxPcZMrnD1IOiAihEz5Ne8yHepIAFpz24b5ineELwJ
QXM+y6AYkP+zlNqgH3mbvOcHs8UXP31W75OgJyX90U109Pb2NwaZna/TLvUJX/ssHNk45l3eRp9y
FeqgiN22g4feMS3UPqc6eBN6UyUb1PAetTwOnHx/Gt1FWwDOPN7IgIvlcSVcWkMVn6M3935tQEWL
SCiOb+Ql8lkWEmK7zg/C/YpXWv8TQ47xpruDFahb+lWkw3dCZoTOzj4LyLYLRsuIFe3ANCdUjrO3
rWXPjOc2W/vM5mKyy72M6XZRHI9cZ3271kR3iFdQxbTP5TVDI/lEYR6M4mmShZPBtcElhwDU31Dd
0xvNjFyOtqUvFGMooUoKit2/WVMXIAZm507ss1LlZTJF+7FKfy0pnJKkYJKjr/PAB+V6TftYzLnU
ri3OzkeEnjeGQn5Cel/QZHVoJkSyv2Ot8zyBy5K6plxItBNlasAMic+QpHlUmZaoHv00Sk2t/VER
MULWYy0kI9l+krv21LGHb7UUpd7V0xvSSqJyhiIL9bfHXtwuWnjLKcCmZpwwv2xmABaGfeWwZTSG
wA5clPpYNJdPZvlW6RVEq0ocb9dNwfRsGHD74836h1B5xSVQFBKpCQbm35djrYiD/q84njhgweS1
3RgwV1JNOa7u9meVytKNKpnWjO+p0aFF4gm+lZ79sgd6H15PfMsKAv0lMpSKoYHzG+yVanM8+ADe
FAGBYBVJiktL51ot30dSexCxjurjYvQVnIXG9Nfo5Kl1ZEq374Jo2NOABJdguw8Kf3Zq2SFxPpkg
lo/tzuWi/vWVVlMrtVfLG4DQvOlw8jz+oaK8t0vdjKIQvSKQEBKagrYoyosoOI0yMSjIBPlqAfSu
Eiuas09r58G+SKHAMWM6HHRS5HPcA3lNGOWJMnP1uT9drMLjf9aSGnH/ThJgOg8TfmpDA3opj2dQ
aqt2Y/Pm7uqm0n5ufJ2qoms8YM4RvEi8RATMX5bFsnbJURH77dR883kTzpcERCCIClZaOJ9NKEsv
k1NqjZsu0AxEhflSMumv6b5eXkttWDSZizPgLwOeQEGWYCIZVDAdBaKJ4REZg5m0g7xjjLR+rIgg
4kpF/lqi9ByOCszbn/0/4gIt+w2Pl8Vo1GU2GynBgU5yB9QXcB/SkqY9glLr+5nTSQ2vS5I5kF5k
u5Ls5LgyVElmXJiXeEqaUh6Dkq1oUw+ry+quBzyP0iARvhmdjgSjHbwz0j23GsmVDKY4vtI0BbzO
3paWGIPZ8hd9h9eP4803Z9tnRLuBGHK6dXIqCzHyZrqi/YOHAW+zc+dPpyWRBuRfM5BMmDplYi5U
1svZ7YAqgPJvLUdZ/F1/FQUFDWfFWvQUlbWv1d99TJJrepBC5t3HMpYXUegc88nAyi82xa02ytwN
cHKWOIYqhacvHcMr3N2Naq/IuVBkKFjUQq3Qlr68TXdU2FMdyWkTnx5CGsnvOuDl92tY3PidxUWt
VtYoJg/juGI7wSpw5HMnhLU80/XUXej4W6OD8TJK8JW+YitdJj5T7sSBxmAG0K9PYEtdjAEad0ma
n2jiPC19ceFIJtA/FeFMKI975t2ChTNkvpm3ItA1DEVtoly5boRABxny/rKUKEzrHqZKSgfHK9bU
6y0wYokD3xyaCtLI2E/9qtM76hx5FVwLj1rSt8WRof0QWi++mb1bAEOgz7fe9q1LO+T4A+4vcsyN
YLNaHGI3N1ez0vPFaWmH7MMax8eUETqh5aJMwXWZJ1rbVXmOMeH3u/VePfP5xNkbRYvll2itsz+y
45UTRADmkOp4efSDD+aPLqv3lMcaJ2XTwlJds3ZQbIhAe2a8uUw/tDs9Cjt8aLkoBN1UT4uJJ4pu
Ndfo5cEVjDnElyiUeFQk9vZjQScDfO4pvoJE1o6+irKftbsj67mllrq4zI6jasmpDo9KBjF0R9If
cKXcbuZ1udQZh9JtWceE0zChwgrLMjCbMSrMwW3W2WNKoBR6izubG+AxYEYlvcxPzEokUuRjMHnf
Zh/+Htwo3hJ7fsx6znlilLO2qij8T+XovO0zJyd45SxtW3eDYvA7wBLnOEplm1XHadxkm7mE2LEr
7fCM8zdZfixmgXQ5S8c3sBoDa59b4CneAtcDeYiCe49ij68g+O94wU1FFXwjPyJakhs5CP+BUrCx
wV3XG5jn447u0TDaZTDDcRtud9SU/zsIBsz3khUBvoN6hR8ve1xObvhnCW4BdJI2dXnAJdZ5kgmB
DZZtVQJbhybB8diFw8zy65bttYs3ATe/5YNsgjp7RUtreXCuJC6ECJa8/Ymnf7EFne8cVPStWCYI
jnfEINAyHOOvo5VxGxHnXBiCVpvLfy6aIn3Hr5R//H6tOL3MByiQmTPPEDqOZ9owz/70mJtpU7Z1
4Qjn58NBsfOeamCgC6ZFQPu1MeGs2KQwOC3KZ8JVzcws8YS1HksoVv8kHrYDCRdF9XyYctA+iOpO
77ReaZIJQvYrZIANuwHG0O2D9yQtaZkTZKD7nccY4jlnwC86za7J4V7VoBDkxbb81TAw/941oQpq
BmU7DIkT5iioJO4R7cgK4RlVqLWFNmzJ0lNeODxJYxpu2vjn+/KXT05FJIGtaeaE9IT3nRxMeIx8
9+bhehKsX17LnUnTketaRsqJ4/Zf3WEvX8Vk1F37kAiF7huSEPvbW4Arb0wr28IFAEhQA1Jd7vkZ
BjaT50zvALLbhOIzDykCmPCYfjhRKEhYBSVY7MpvED8Nix++Qp7tgKDH+Zb6g65NRH5DjGdNX4LU
mlBGii7q8QA2Ck2GFgutiC7WGDGpOY4LGsA27HcboKD5YS8TevUa21BLuh3KluukCVZj9m2wLr5G
xfvEq7NbM3rwCBirc0+wUmrfssil1NA554IvkL8WrMa/TQMjf/g/yCw8TAP4yVMJ3+onc2hdemZd
Vp1IH+1NLApNNwfCBgNH2FU0pGlB9iYtxw3uLn5Dq4PHU6nH1bhMImblbjj9rQ1QZG4+y1RZHcgD
tKFTNAKgnNI5B/4TQI9uJlCA0HloVqe1yDAR8VtuDkQyynI8zJwrBlqnST94VT5b9JTZdjqUG4PS
Rw4koiHi0nu6XfEgeVzsCL1plKjCMNBa3VVtmLU7dkZYSH+cgmGGOYCtH1D4suqPWLaz9qmIkwQh
He04e5IDVovLKARMkxbwKAnjZwrn/cg3aKXERMnb2iwhg+hB+S5HE60LpcWmWn/Yj2JeYLTW+w4k
2qfWEkdP/EUexNRO1S2c1NFpm2SRHTYr4k1FNVuzqHmMm5qPv4rU0eKLyOltvMFvOTASBTgdIoqb
LlykEvI08/WwFaO6qoSsvXarZ4we2ssQ8dg4530P1w70g5uldgh8aLyAM7BIeGcxRIhj11f/iZ2n
tcSf1wfcYdMXuygBHza7zJnrHGX/CWZQGZJ2jXWWOPSzhbB+kcl5X8ntrarJAgbA37LkAn9H0vlM
/lGVHF47xvnopdhrBxaqcBZ6dqJ8TMcaPo67sv1dRqBmSFdKehR0B63BP+q3qwNnMb8iXkatEnRs
1yiUkNhpa5FzbUZ3FblpRmwmAenDbnRYBc2ET1WdcDNzX6ctlJvQavwbRm3aug5UZGUma92F/qER
4CRjaccGSQFm7yHjQZ5CiI78j8b+hnGOwU4sGYKVH3Tglm3AuPMYXb/Lvr7mIAhVYLANUBvfHpv2
IFk4zYothIMUb/Pu3HVXtB8smKSu28qAWRH5oNWMJJNE5pum8XUOxwix9xiMEYoELn26ppaXDG+V
8Tu67hiyj51/aaakS9Qli7bhsr2un6Rdyezsf2stNuPFOHXVsl1tyd2RLKFOLn4Ca1tQlx7ss+19
4EcM09uBeoUgzCye1/V8/BYoZziF6pTTwk/+U9Odcgrmmx/EH5dr2ZxxINhQ8ku4X9jJTh881upb
THFAsCa8qTiIK+/NaBGriSF3c2/wNKoWybk4qYRtQZjxKYsogZWsJKZifVgFzzcA8M9xtrqnief4
I46MaKp17XWyUw4BjdgPkRFEO/STf2gGCtKYUc09kGQb8CixA0tfnGCbGhu0wN9vhI7NMKc4beth
h9JrW9DUfezn8dbfOprwCP9Qu/mBKIpMG6SotP78qqA9cyB+tA8DmZEXV5QnB2HkaeBWgpOZ1Xqs
Ds4p4HnXrJK7bsY0qxoXuYUxCFGW37aT6ti+zsnsjvqZk0rJejZ8U//pscYR8wwgAzPsjQ14KUHR
fldnZLegGzvIq2eRPNUIP0jKGfa5k1L5LXje7JOWZ/EyVVmCB5CNUujLvK1pHDKMscJRgO2Z6VaZ
c0zRhlKwmVE4CaRQttYLeKWf80AJLhvxywNQw3vb63mxiB2TSMYjHdCtnFQWF6Dzr25n/eopwCov
ovZXYheUhN5AvIiLSire+gAG5RU2HtOCRKjtkec6ZboOZSqTidEHvgmLemxbKxxuOabXq+cw1WcQ
2LVIyoE6Q1GsK1w3xgZOvVgSDvXOXDu81m8w7XykQEUNCehN/bK2POiOjIyr+HqFyd1cmN+VGi8j
SXqURFHXpX3ypAdwUpTWuA+e4a5E+DeCo5zYRIzWUOYwwk8Dv8mYw8MRz63tb5NWXZwAE684tgEd
8W4V7fipCxXzkDl4hEuf+C64rAeQxyY+ghrS5kEwAm9IYngwZ6jtnQ1Zw8Yz4vFgNIircR3PolWw
UYD6NPDyFsftK0McbExMV6+jHzGj7gF1Gy6chTfvrPMlAI9N4cgTF/L4m5oQWrtvCkXxTv5XKdT/
apG6gJoVKlSvg3Mr6Rl/SRhOFaj3QI9wgur4HlCodbKiYUbAZp/xE35Jfb13qWFXdLoF0FNveQ3M
NHa6eC5d1JG6YkaxTAeda6qdkJBAiquPsHu1/EcM3WtCvQkmaoJTijvZoaLB0fkql7vHsYE6ASya
3r0LN/9TX5tvt8WfGWwEIABAKrbeD92+eU4IL3luKaaoibC990YmIPjQeCcVEM5icG8s//DIb31O
fOY1XJHo/iLQnZA1g5s8dc5z3V94i4tmfcUWf1fiMuRSOxUsTcg1ixuMyQUbIfQ9t+CjSqzvupCl
KoaY+LZfag6yTorV5j4i9ak5eWR09WEaRf0H/OIOWAN5ckTPDYnWKpqJp798vh8ceOnldFv7ISoh
ZuRmBNAtgvGXXoHt7BL0b359U9aGRsv5hESbo/4FAJMVnkRrVpGq+ZaOsXA1OQL2dMFl5GJaAt69
Wlx7FQrEn+XOey2q7cq1oueTInQY33CK1HjYg4iZLTDuMEbO8LlY8HSUo/vOsXnujXhsKIKdUeTQ
h7HMxIqjM/9ckuS38ghyj+88WbK8vtDvitgtQe+wrHYVIcsMAcP7lPEhpEb4CwLL7QUjoiPC7+0d
oCAoNMK2YaPXUI8DJHF3A0Zy1w/fX2fr03XR1nFCSOf/qXBIqMg5ntAV4E/ci/ptX5LJuI/h25rA
14yuCSWUfZSN350rjpe8rTM3DM8XD0MHM/18dsfgN/XrCLDOsF/he+VX7UqBJkG8/eFHBmyul6PE
Rq+aDFvMTk0VURrKlyw5yliyzgmkAKonrtsRYQCqVZXbrb4W362qUqvEVBagbFrMDiNK/bhKA7/I
6iCQNKlKz3jHmoDTpwwb10iCm4zvnznE9tIBe5fRI1wFeNpaRoua3PGMexuk9Wbj8WJn02toB/BE
OeptpmXwFb+3FpBbOb0TSLV/dzjlv+N2zdEloeGDKMep3XkO8SFK12HBv92KeoU2ft4mIIXPXVK6
fJDBUc5UI+fSZPvtCS02+dXxX+O3JlXx9frJ+rJZEqHq1ZeSYF6Eax5+ZXfHC5PN3a9FXv9BerHA
DObYvN64c24D9RTyhVB0jvgkJ/msnAtDidpK4fU2zbTyCGFNgsEfZXYtsuNeobrTI0p6UXUMGoOT
FHLWbbBTWbemGjzoJuGvmuf5Es1r9PHKorW0WywRQu6s9UopM29Z099Pf8t3SR9Dh2yW7EYlmSgh
57LENnb0jK976DOtYdQ7pU0XEHvidQkpSBdvLDuvbt8im6pcW5WTI2DvUakA5IWBmB1CrRh2tNkD
08fx9+ssBMn7mHrSkMvYYvYq+gygEo62E+KULJ7e+oJGolYfqodtITV+TKImdzksPF1LDTq7896A
pfrpWm5b8xC1O/tLCil3a1TAJ25G/Pe8pcZ5ULRcq5eWQeLLbXq1WB+Xt8j0Wo97bSd+5Jgpb4Pa
/tbe7ufruoD3d7+RUyAMif67YeAYFsJOc1hWYH6V9pEvkumld9xbzZLpA4NflVJ6k2PD/ZRsS7D4
MzIacig3Bhr6IpN30OCxKFJj0tn8RRHKeZ/PYxFS1YiwjgMk/efQA5IN0UGnJB6D+ABefhH1IzQ+
NfkclAzFnt2cOIJO3ohUvSQT1OikYlmPwffxD938pc9IL5bwEl0rMYlhb/ChrcxsFPrWRnn5HHqj
/OsZN4MZEZyqMmAVLTGlQuAWaqbuIUyPtUWC7bOyaEKbypQGMg2k1nD32zFBlucLzKf8tyEFhfNj
btp+g95sHN2UWVLcyH4SIIRXv7tEeOCEKsS+Ek7tVAx8m8HpprWNjzoX/wy9z02U1kuidvEamalg
/fsDzPHYaCqP+i02yBg4Shb/CKiHXZ4S+DKaKcdSwx3a6Ax6H1WiTHBjwlEuI/KN5gfsj86OEMxN
4hx4qWJXDhoN1oojhAH4VDALjx+Q9Ws7omaX2LnjfvymdGUPmCIAgkWp5rMaIP1KVyiT8naa4+re
taaDWn3thWuEne8o0g1KJjB3IfiYJ0HtHy+GdG6KX634SRZlMzIpCSiKsF2r0oaqaJrApHY+jxrG
sDFfugsT32kgIEyGZ9QQclR8gjcgUveeO+M/CGT+nnAOygHgz4dXsv7GC7K81bJkHnEnV2BqpI0T
CzuhR7l0NIn1bg7z+M7fZxdw50edYpwXab68YGOESJdleogN577SGSwUeLZfseCN+D4yQgTFLzBg
Diqh4Ylf4Xw8HEwxqtVSVEVOoVolKyFPlsVqGIkMN4dWqGwwGLvSd9NEE3w0sKyRLKzsLDX//8g6
2eiJddsrSEs0ZolJpjEuiHg2cJVtU6GC3TDxSZphRd9VXAdDd/0ObVwB1lOfrGoVPB2YFdM+b2vK
C/l6SOaHZXwcmqlD3ukhp8/+qXXVAMSup+kaY1yXtCl+GANeI3rSVK8FuKXoIj6AnkuxdDL0urNE
N55CB35Hcw7zuRljkUVTPF4u3DtNyALaWbaXiNyg4zzv8rtojoOjzAmoD/aVKjaftivoPdgO3OxQ
rTP47yz6PVSaBkVUaEoXEJfd3lRlhXBZcQENnx1y1frAwF5AYAl80B1MDJYVxODNvsPew/w77sgd
rJoPflunQ/K/D7GVrlBxIJrCaPDv0oPsM6+EoD0jPae+xdQeFboFBTSTY8KmAVaFWKuyQ6pkbwo9
NykwoTffT8UOP4PuV4s5Qu51EyO96zoK4FMPIZKEySzkCHXlo1scDr1CdLeEABPJ0WSOS9enMiqP
v5Y3X122JGuvtBacuxH+yT4UP5iWO6NX8IcZA7w7nzgKkiFpghs0amlLLE62DnjnWogq67rFo5h3
PEajn4UV5wDjOxJDZ90mq7QVFdI6GsiOlzTvElsUoYjIyN9LOec39dqehuhusluxLSJDM7txmEgG
XgjLyWZbW9mponzeN47idUXWHCBsnyMDox/4/QLU9a9z35reaY0wZ6JmvhbA4JKTq3+YGF8Zvq/Y
o/grSy0ZUbVOcmvbiwrLYYJ7kAEF9sVkaPXNVnTKylWbPHYMo9uPjhR8uDJA+F09Cr8IZIm+hzlq
VF3yrZab0HPFZ6KCQKLnLis7NBBuVXZlDZIEWQMNah+8fayfIhAWUL58sS3YBrzNipRu9NAO+6At
YCsW/HKOKHK5s/e2zwwx0JAK85nN+Bjr6D+nDO8rA40MCm4eW91044pvljqTN3sK46Y7lsQgilfD
y7MbBAMC7fXg1ppzl/q/Gj6qlJunrVkLmdO0YoesECu7wMwLIL75CZLVqeK7eIjPU4/Pv9uiz1ZW
jLoLsnQyCEm4Z9BlGeUdgoxbfur9/ivpa/zOCCoMfjxAGO/+sj8pQ5UDbxfmJ4SIWJitF/s/mBC2
cCG8fJMuyzQRnKJb4jGmtL3E0OBBnXHtxHif+7+vUpcrb1hVjcrlEzoQCj791p/mIHwJZPmWYJtN
h/3j6a81Dl5tPuPMc29Wm6ZZjssALvE2boYGb1w8UBFCYo8rFFbS1fbWt1N5yG+TEy97ULAnqPwS
y3MPijFdBMva/ylJTvjEy3Ups9ij4Gl0Y9L84R5plqeTLFcaoAqmhVIL8HTYFzrIPegZRtl2S0Zv
mXbio/v8B3dx1kCfKq+Ua8RSw8MLugNGxQTUDBmSPeW588sFgS25TvptJNfz4Bj0VPQZDic/dY+0
bH1Q5sRJYvqs7Ryzh1pEf63PbzvVAS6/BZsFl0kEZrmWiQ7SrDd3d2FyRhK4kTDuvBuIX7Nw0Gl7
Eq3OPGzGc8jx7sgRGUDIGB41ABAF/T8L/J98N6c5N0QNuzYyhNUfGiqva9tDqoD3EhQXTNBugaD3
iqzMiv53ov50yOtoiAn2KHUKg8z7NeIn5m+ugWINC/O2E8Qua8Cipuy5MZ5ob4tHDF2noG98qWOw
Xu3ptsNQ/wAVBV5gkvjJgOa8QHH8mp9Zjgrjk5O7T4pkbE+JMexdlPuxOMrJaQIvyOHVVFHXhLAW
S136eaJ/VHtSd8oUhA32Jt7KJO5YZMj4O+OllAKHntTE3C7D7MygiyDN+SAGnnK6akYgsDMWgtGO
Pdz79UjY5InlaFuHI/XNkVeuCgVe0ubxwh7FGa8kKfBtkWRBgI354+i0oZkfYlrlsYV9EZbEJbq5
63JIFs1xI8fXdWa+SMpT2JnbOyzDY7V41FLyT62XNiRksU/cDOczfMjeC+tHUZJ+57Cv2i/saQgJ
qh528xhhauM8V98Bh/g15QFk4MIBxLEn0HDAC4BhCzgZAX6NHN3QGgcZbhhh537D6kpTNgmuXv48
VxKwI8hMtP2o6A9lLrkAAxkAM+a84sbXdekiZSVJ7fgKLW+348N/AZ/Io74g2rIhIF5UubJci/p1
tpnTm4XBMcx4fp+wsWPG+0ONHLybrKmJusnhsgm2u1DCUGAgfStb9Zc1ssWvBcovyD8qLbQm5OW8
mWMM7Vvr59iyBKgu3LmvF2Qwo2NItWGVRNfWKH4W1EjY7Gc0qlgk6Yt5kGBvYy2Lr/fsblznNIHx
b5e1yzkgSUKRIHvIfeO/tpQPdgVyCdCudYJSZGV3LeEIVNzjT2zamAX8EzImGfH+xKbNtgmhnczD
001FwZouWUc4vamJ+3/9l0yupY3ukfsXN3jlkvtfykvl3XqGVhJPkrkfOk7r16xXw2kv9kJzthqK
Ej7wASyCT1LtATD+eojMp7THuSPPp7fL6NaPyrF6+DRDg5WYaY7q7HQnfJUdUemAXEoNSLpzJehS
jMDqbWulTFB8P4aHYHDPuf9OdB7Doz+JFVpeAdLKzS/6WQOqRXqJ8nksvhSLZa0LzFCUoOE2JZKP
DM1vGeqNoKTW7dPJK8EsPWgDoOUt4AFKEql0ydp8PnHX5RgxKpGOO2juGqQOk6UyTjlmBbwEHOgZ
cJ4rDBMlGHaIcL9oohW+GoEDDVQ6nyzzOADCHhYliUg9K3jyjTV0x+U466SG8VzamZFHdLfpbyy8
cPK2I2Kx1HHr/yb3cQuTkNFKI/T+l79U52dlv4KKSLma9caLtdm+gqOZAyjpXwKqNGupsr6E62S6
q6tlHDatExzcfBNiGULRpx9Tzaqm7FgAuzgwWdvCNbutjskqeWa3CnfV04NsD5CpXZzFAgZCTDMy
XQhDOKNfTh+xLek4dYbn+PX/DuslVopf1czqjv/FyvCjwjN6OmfKo1nPqT+IDZMCuwonanfQr81i
F4FaoqAyBdLNioRI4doEk+Z6O1ml/iYhKPaXY4WLp7HjmbXB8z+y6vkuqKlGCOPaVzRyCNBjIbxq
QrbO67cApPb0lnlsysXsOiELh13bFZBgzBCA2Tt4FPPRGWUYNdZfFkX5zjkBiWgfDWv6OHqnhw0z
lqVILCAsLi6rnpFQsL0Mc8LYK0FRlPQZ3vmc/7K3NYw632PeFu0hZfaRLc/hnnogsS5cABfrDIxc
adAKPIUZuQw34JNOo+G/J8D7ZiI24k2mnUTrfJ+plbyqyE+H8F6OrqffKyrStB5NUE25UFxb42sA
yl65TVGb8LZnOeqHiwgn3kIfC4zzo0NKzhtNMT+f4xFP6ZTsyJR3Wlzk40nVdsuuOTltphUavn3Z
oKZQQj8X6rcYdgbGh7rMB+KT/5npgIwMwESRYDp2oRwi1x4bG7TjIwxFDH/P3k9kvKQhEgDwyVPb
tv+Yl5ye86i23mx0MZ1iFXsqU1veIYjLHoL0esFqef0rW3d74KXJIcRgyVk7PdTf/25r2OfU04au
9y521R5cd7pZo3KmdWNoeOCjldAoEOqbs0oaRfdvI4SYv1r2mTLIDqf/it29WAE6yj9VFzT455Br
LD0UilCz9Vs/hm94KcTkx/Y9iUoU3rFYR7vJP18dmvHZVG9fzTi9PaUEYenq0FcgiEA1L5TvumJ7
CtLhx0gDez5YVBSzuDIZzQDsO8X9Ygz68VK4uOWFwrtT3QeaNj+E40hJF2JExV6d7D+yDfp4S9K1
7L6FTXbFvJvqf/LE16FvCPvLQDSwq+lZJDaO1O76bD8ZU0GyCAkt/y/NAlgIcoIIYOe5RmYgdCIH
CtHo0hcO1bTNF3O176zpjrfKElEvgL/0QnKmvz8iT8HvbpEfbQjmViM7+dXvLw85SetlOKq6YF0z
J4p1P1mlctFM+BVl2YYF+saj0RpMmqLpGpLDA2iWRxhJ56tORoOeO9dCMyl7pcUSvKbt4F26nmCr
LcbwX2QUHOBqrixkecwl9ghE3Cf0ocoHmBXh4jtvYYUFLxGr2gBxCqwoAQUGv3qUYzIUvTDVeCa3
FSHOFm8cMgxYinU1vveaeWc44sG1GUC/HEXDA6FQKGBR3OWTgr/mtwZaspBifnra6S0GojBHauC+
XuprUo2ylaE4OX2V8u6wDjsJo7Kxxkk26FSywLzZ0MVXwQiQMH6yJzVlXJKyVRxeFZoWdHm30wsX
oArfLNC/o6Opequz5EFq9pLIYleMsI/ajVd8R2LuZVmmH1kiJmlQP9B7ceqt0UuF0KnTL/Na9wP2
2H8XTSMLiZyp3czH47344Oo3gjYYpslbn3N3ybJnVUYZ2iCQYUYE70AtElqCkNHnTE8Pu0u6JMhR
Sd7t6D9by2lJUTHr1SZ01xYdDeVFgaPKorHsXn6OVGGK/SGD8xljEMfuEyUs2xqOQU+L8a2dmhim
+v6VyI0aFG/kkqjgCRVf0wbtxXOh0SmUMjCNdMPjYvjWqYmT/C8wfHChhvHe0xnCt85dofJxqpgn
SBsofaHIEAt1M1ZhcEFnuN41vmkaWsW2xJVu/94c5s0MpdjtP6Vncs74L4qY48VEKPzK/7T4p6c4
QJT+Yxofubqyi1s+WKldVABpj4Dm6DRMNgoCp7L4NFz8QUf1vLr/jfzOcOEXLJELlkC7pvT3A7UY
fZVE2aDIDrGn+JmR3+/ZSmyyQqgG7GzZsgT3WWOqs//gF3gepUlcqU+WtYLLKORaXXK0KN2NNs4/
TH3/Ki17ufWIWodNLiZRvsRA+H7DHll1iGKliB2F4jFOwnzQCd9Qc3bfVFswQSojLnPFgR+fCR37
tM06KAlL+UOZK9ROJLJFutUtZ4wrPkIRVV/XfXYNkAywy8o73XjultZ1u2t587ToAH8jpWCHu4ye
ZTdoejtw332zIj9l7Tcq7+jwM2qD287/j2ri2yQJ0alXkdkOKiAgZwH6DZBfe13q0/f2ic8IjYqs
wtkuCxnj4EWFb/z3Q47xPS2st5FBen3WY18/utczg/cNddZCi2BgHsJAVyKKKf4ZLnRhbSGaV5iD
hiBQ+HxnKem4/eott+C73fQG6bTGGyLzhR/eT6zCfysW6NN6AJsow99RBij9mPPy6RC4/YfE5EYT
CduYKUD+8KLjlcIVsOhdHY2LgK8+7M+KWkGpT1SpaCII8oV9neFWZMFK5qlZv3t+jsEI66fM89Ej
Lbq4pjBnExc6ZQEGl2gBCTrP0qL63bPR67SuNN4TCv6S+n8LQSEXsmGe/lhQrljZE2qd6jvgCMe7
JH9vWzZGoVOwR3K4kdpQ1pucp2aq7DZzMuyseztxezx4UCiL2dP52dXjn3cCjn50zUAdpXMnmlVf
yLyRFAsebiuVub8IwJnGsWbiAA03UptTXe7LY1HbsWViexjf9BTgL5cOWzHNYE+I+fODgVflx4TI
y8StZuY8rnkpDkVSV3WxxgUsDnJGVqHK7LwKTIlFND5IQ0L9iQa5Vqg4noB+2I7H/Y+F0do5Df+y
rbmv8BhuRFqe/rG6NM1jDQismWpglETF6nC89NKa4pq0h1RhlxPuWCpsGNwDKoWBgXZfGGsojM6L
1HbFxjQlxrnWXYpwT/cvCqzA94j9yDYV133oAHVc/zJvF9cDiWduuemB3L/KlUPERFeOShbpZ9sb
fZlgcN0NyxTgBdyHaVdzWMufBUwPVJbit9Sf9U2iKJldtBF3nU92943zn1816iVNZxi3/bmgPjUX
tfuqbjeNLBvqhoSglUc+2xEutUYTI813QPvBu/WZEfZKdgtpZiitpLM2Rj/Juar3IHXlzLAW7iAM
7Q7dEH3tDZ00m4OU5SqVtIHPhyKl21mWdqPCBnZnnE3y/9rc9iV2JSSNk4DTbOBvs2BuKn6eXl4E
9ZkpUf+aQyD5WzYvYTKkF6OzAMs8yXVzPcDxpThzQ/OXTykTF2Dompe38sNvP0/iQm2jBrMmJtkv
iav8Ke/qlMZ+jUwEcS20K8tCEYcaJYPKUf5uqKsSZyUGtRl9AQKTFJDWchT4MV7DulMcg3Dh8fNc
MN0Y8NoC9QdR+w7t9eMjWJH7zhVpTb5hzm10AeQk5YbdYgN4JBSFoKfqiAegG3fMytCh9ar41Pz3
qYBlDRhza0LJLZeowrylH3cG9AL6SdqOSum5ACxJDVwYimVcMyTMqw2+UW0SWwNP5iVUBrISAfWr
UN8+x/hgsJW3qrWfB0Hc6eOpzHgdwZbsKyCu2aop6Mf409BZb6Cbn8Tn4IMb62QIJO8eKT9MYdUj
PJSbXhOnGo2t50v/5oEaaTGfG2d1fvqzxqKrn0w9UVSTDk30K9Tu8+5foAOBfryFb2g/AV8FCBBY
1MWXAWhXdbgb9zFA0AKRqNwMes0DwoBtzK1GY6L3KsQmTwjxUym+CO/MVnrPbvOM53WKeeBsYrlW
wlb6pKlkBqbsbKavLKJE6av4eJh3nIVMuMzbnI6MIqSbtvbYSi0SP4h+jVbDPMfAzbAplAoJGdu7
QTIdt9En6zxWE1Qi4JTpYOduApAVf5T+/MR7/56bRrh09nYC9H/FAB87kpwUHbOQCgbDJf8GuPyK
hvHrrB7UwNY71BN8hFvXflvM+iRDloCYru26YyjKwfFB9OQQJL9ZoJlH83psX1SgtR/rMoQOK/pb
hZ2w24t/WPhO9JokKeFB8NvSo+7U1Y70gPOyITf0+TQV3CziuTGQyOEvb3ed6bONQp1t6iAIZZWM
K4Yuu9LHsUq2GqKcIDhWkLVW5jWMQP5imkgK1RxoPYrcAM6BS3zxKq7/KeSJB6UM0CKbswoK9Izu
rbiBqgAyAOnmvum7YhyNx46DKgN5jjPs0mbUeSeFetQs5K6raIAxJnK0kcYkA0LegRqmh7I/MreX
+A/06bDjIsEgRMeD8SUdjNSBBZNfRFwSAZLtYY79hBHGLLq37GLAyBNlzZVSmC6weFJMPX1RNl3V
hg/2cNDHqBA/r3aVa1RY/ewmAfbRPYVQSVbNNIXdst90GL9ZbBmhnfCsVZCIyrATxQEOYVy8obmc
TF0oHxckMhdQP0nbmdaBTTRr+K9h8u0NmQdTgLkSJlwifBk6xl0VJGhDAB5LIesfK1NnFJqh2AYj
RioSFjRwQsBSndnUOzXmGFEBar2J3AbQx+ZejhW15vkGsRXduKQLoMAr6e6Nki1Dv+J/aoHAQbQl
Smug+Piez2IXqh9wLMiRoSMXsfXnncXBTSkBNgWKUDg/9bK50AKRjK82E0I9XJo/bVZv4/KRc+FX
LwiiUhdONYYwwo6Va73dHZTUra40rwuYpzfekr6CdCeB/eJ63aBIozEiCaZExrcGDp/Sh4jW5qry
LuIWfnE2lx5K2C5qARsyilVeGKL/drtDWkiB3kDv8nEuY9MOl1QNlO+FmywiINNtQmtWWWIPaZJh
ifvvHhuHDDg7WSeyrBgNrTXtxsDCWuTQUnQiQkaIXruouHFwO5/HzTtoMQYocheIgHvwag8qdny2
c7+SxRbM9sCfjm3WbJELJsGtRPEoUlgilW6Ju48diyGSNCguUWnI0eCfff6hbe6z5wmWKo/CNY6K
wfVK+R96Q1eVPV1IFfJn94/rcBzn5u77ikGctW5BtG/HjnpHRw6bPYFdIY2w/lvtwytExY0tpDc+
HnddWjdj94F+QWRhEkX4YO5sxqECjoKdSYItR3W0O62FKRNTnhSTa+cqM9pZSRzVUEQvbWxe8mwq
KE5AFUhvftoNXM8O6M7OZFec6GeZMuKOyDfJ7jzVWBG/A728d5o2zm4vBrsw+mCyTOV7Eqc+9sqd
gI1TZ4GXWwM4qWLVqMoY3HFf/7zqKtSgSsh7r+Uw1QOE1lWmu7F0hmccGLVMNRFB3gzQyVfYryC7
MwlIh6edFtFjAk7dQDflgi/+Z/tyBA4p8b1ZsGY2qCP5nVPZTxiqkF0p/UIIjHRoIP4orNcSyF1N
RLqgT8gxoxnbcOHBb/w+gKIDd8Vh5E9hcNgsWdD0Eowfwrdjyg2EiTabNkEQXBI+8nf8YNSW7f0Z
5w3VjYnkGZRNGTMy3IUkFZwyNyjcdIk3oyAp/pXcJQJ7qBydGaKeb90Vnnm704aGDagZoiLRw1Dq
b9Cs7wXcU/aSp7bR4EkhJTwJzLEJq51e1ac96X7xLnR5/31430HbjA6ZTVF2ebD5CaAxmS5D/CC5
45fePCJ1WpsCPpuAoKv3i8KkCV7jaBV9wCfInPCnApXicEWTjM1jddqGVdXadXdsHOfG0RX8kgdX
lxN8r2+XBB3RyWP2zCe7cqEyPlXgH6MwpKQeH8Wvi9kQaodZjrPHgCh0MtDi+9MGSPEvbViPVku1
vcAPZjA2iQd+EGcnE8q29KMnfAKCESMdlpw4kvNWHoDzt8a3syhKGZj8aQRYvJhAGrpuW8zR+SLc
SdK+54mXQq37wRivSPLC0hhCEa98FDL9Wl95O+kaCepV27VqAPfazsxGY7JoE8WsMt3NOo+5bAxM
ftWyhp/i98NFKHGblpjISuxk/GKPPAmPO+De+KfEafYPVMhB6Ylry3bg05EK3nYx/IvwcpHUEImC
PqptTZN9IFo24QqpGH42i1R+YeYTb3LtuzKJ2HyRgoApMqf4MhdbcFJQa5hmTjuy3G5Kke/HWGdQ
fX58WB6vCBitCRfjxkdX9VM+VXyfFT0Ha/KOuszVcse7tq4blIf9bi2H5VDykRqfxAa8XMgnkqEL
fVJr+R5BlnI6YkHlFeLhGyRi0TRylUHWeQ8hidrAckQkkvVNiIRPXkoVo4FMmsTjD+WbLuyJBl9W
SG+RFulBc8XEcS1DN9YbuUVS3Bfub80LWB5lnRUNKK6OHTqvGpfrzlJHeIW0v/a3SiVnHFYEJeUn
+PDu61FajOjShLmGyuq9XyOOcA/OEc1DdQ2KR2QoVY3ppBCzsEpKrkScZSpZxFT5Ds4qgQc3nglo
rMZs1nMEPcDM73pr8p60WpEe2UpZ7nxzfnitN0stsmSdauwQrD6E5pcGaTzi1bRLSBEA1XYe4qnI
N9zH9v8DGWFtyy6MSznUlnY/z5pVpAHoaH96hp2saNRA2j1xIP3gfGdRm4llGFhaVbvPTny05ATO
hTzbmdIdRT/iPn209tZZ96KUA8O8tSnndw6ZZD3+jxHrs66LxR7xMY/UizKJ+Zjogk0xzI06VP5O
jP2mdPO1g13mYqsMWmAeT6zKZrkx6S20UAWeSm7C9A02uatQS0zuryeVdrrdPAKDlZmBg2Q6NSZj
+mHuFAbVujvwp/B6TZ+pBV3nUVEF2e5wuqhRVkr952g3rvm1YkNt7eAwAcl0RauCiTRSOGJjeAOw
bbfT7/KIgZ5apl9/5I0Ddsg/SD13CjPvaekWNpG1ZdnA9qXC6I8DYSfOrwfct7wlDdllPFJtPmDi
ilDDiF0cqOqyB+171o0fNy2yHodPQSZvkO4/+OYRYFhQhIkzxpiUZEMOAfjiZNPpwkUkRcbHXicF
XDPn3E/r72GtckkZrDoiDs11f9Zrnswjo+4jfUWFOcerM2eAo5flzDnucE8/717AS5dgxbCJpEzs
YZ5zpHp+re4YDZAH8eUGtGWsdIBIMmSBiyCkHqjak5rhC5Q0mK9RnXXqihXvp4O9rttZrOLoBkcy
HauyKMzHGeyhO8i2shhGa30+1AwaXFDh/LC4W1UEaDjcRlOD9gSczwIo/CBW/1WV4iNQ4nDTK0kY
tG78xnXajYSG88Jti3mcd5Y4QptF3v2esrCxTqg3y5JAYOD98y2I8uyL9ZUTN4Jb7nuseV8kYgKJ
V27ioRBiZtWApvxbO1H0PaGr+kG+i5xhgdxcelIwDhJ9KjLt9QvgpTy0lykxhkD49/2svtd4yfrQ
qzmnShYC1Z8P8af1GqQ0z6gkfC8erler82oX2Zm5Tch0UKLLdOGc1oznRZmkJ2r67FlHnFQjxGYp
Gjha/Fz+kGvMRtwUboTbCInEL4BvGS0PULaxj1mYZ3euIF0KF6E8Y9P52W0FPX+6mqOJWvclUR8j
VyyPhfs7xAEgWBGRF3rI0EiM9ud4L+ATOvzoWM76Z7yHRnM5LjoxRJU2bs/VsdrmhcDiRM9QjkG8
EIS2gLNcbeU3wtA0wiiTCGdMiV/hJ5lDsAZtyOAurkjo8ysGftiWLTZBbxOaZm8hNGlGgV0Wja+N
7HmgXijFHLRluSD5l6KFKC2QuDbOX67II4HBP8gpke3EokYevqOwFn0RLtG/4AeDXl8ZrQU+AtJf
4nI1ZewYxeO/GmL4hrkjxWnyySpcaHvSgAlUdyxKO7L+MYQMRmu3ET/PawkTlcjV5plWqfbcC/t6
zPzw7LziDNHLT2mIpJKGwDeVCXuG/z+bRy8pCfJaTwTRcdR0S8cLDd7YIwi0cpM9A6L00LO2q3AA
A9efyAFUkVFojXqVR8S9VIqF+J/7hSsgb7gnak5KEmMuO4JIkkywpV409eVv7z9f8FougqkCOZHo
2u6RHiKQbZmYzZ62QvIdl4GtDDsnowEBmOELQsuA80P12zHBIUHzry2mlql4cI1DjVQ1Tnfp67gE
vsRptrwA+ShA4hWu3jf+e/PhA2LDL1bUkHdHJu/OJfj20WaCBFRKybFhdJN8SfZlS5pcmg6S6blZ
XU9K30mIOE1Vnwi+HkEm2rBPjnVTYHgfL05rY9dWKYfIhIA3mYDsSMS6YN/z5HahgH0hZEIcjBrc
7S0tCrGm35ToIG3lgyumsduhAV8/EZaKx8c53ki9ntB4D/VKVGGzBSqqy2qjsAyF9NRJ2I80sUVv
gar9sS6yKmQmrGA7YHie/C0QwfKo4557i2bybiPD05erIeGqf1OVQPZ92GmOO6ZZBknZdC5r1/1R
mk6tV+cJak+B1t2MBxgk2OFpcp/Tv/yizPWa8xZHsjAkXsON9Fak8X7B8weAXQWAne+e7M6S+/G7
FP+0BRgBsmAEcFee7FXDxlRBg3I4Yi+TYCY8qUz9l9bXDRFL2IBpWpMakM4ajdHRzn7zLWrJitul
Cv+/asIpdIurQ4afaYPRJ/4LveKacKNgNgcCroiS/3zFftBToz8UObz2mbb+gW0AO54d86esHO32
A3KkVmmEO8/nECDWHh8Wfn574Bq1Q3sIXikp9rEVDRgeON/pcLUOabolhz4VDCpoLrrnrwy62JXg
y9e7Mwjo7e/icVy813YZvuNgNOwBLMle/16gTK6LwEeUFN0j0U0vo8o25NN3G9mudyWyWspYSq/U
o/TZsinjEb/+SGEo18R9EAUB/7KiB8qzHVcx0nhQprZNgMLBwoLM8J/IKq7lA2pPWDIvqxbeyrff
PF/ze4evBe1RAAZKWhQyrlyYY2K1U05tZE32gvQO9MTwu3F6XTGK/hDuj6tCVaM6kNdeYmMpuGXB
ofzwc+NKaJWeivL34B5RGO7j4pO4+vVE8+vfr1he1THw1UB2CMF4YNFwAkU4hZPRsdSb4ZkSTWCa
668sdL22nMO5EmtN7/wAm2Q+oMbN+ROQoDTyAAs7Ez51+07Al3ZxCll6pQLuuJWH7hPC8neVcjAu
ANwe8cJJ35izo/+EVRhH82EVvX6P5hmtuhRPOjOCwq18ZMn9ug3kx5KJNn6nUZUVfVnAI3TMgRNp
tfWYbgLAoxZd/1uN1hXQLEXorFacvtvx4LbomhOCOayhfsxmCg9u7BuljIkZpAO9pOFsbwan3dBh
d5RM/cw1DvCwglfrmFqfKJdzg1Wb4/0ZI+SxLzqf8+iIXyuJNBOOGhiaOKg9+2eRm2iam2H/4/9O
yTOm31CNOrVcXGi0BZovVHQDtD4o+mRJDb/cFL+dRkK9/4eG5uND8vgZlXNdqvJ/H52Nx0ECbvhQ
O1TC9kTJJcc0lwJHj6cFRda5y4n7eq6QyhUK0X+zQXyi64bCJa52AAJV9f/AMW+UJQ7n/sBmYkgD
6yTFyA0Y2YUuMFT2RhjQu/M1pUUK1hhSA+MD5xDRgFpGcAZMlZ/pDuGKx1Nhe+i5SvQZvp5fzxE3
jq5sy6Hmy3AxrG0WSBfjcD/GABloZZFv/bt8Ua+Re3ry+oQo7TrUdPAdU31/CRmK4ybVMRxArFM5
9Y8zsJNgD/1J
`protect end_protected
