`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lItBesBFYZIcBDyrjs4Y1yLA7faTX4UHsDgohDI48/3yfGYVgP6EP3Q8FRADU/6hetTSOYBg84DHEAUv0mxU6w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W7aGWCItim0nLw8oEH7seZIKy6wDBHhH/xIAwk3Bry/HhtRVnCif3Sm8uRsDqFh8n/OgohYkhM1ov+JYqWgp5iPFNDnJg37zJW7W/NqQgVfrQQvn4/VdV2Cs7aycP3vN6Gt2vsluRG66HfWRhDOy4SWTMREjXbHswaHQmDsbzKo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oIYwpqcWJZLEXidd+XVjYutx59GPBVYohrW3qu4Lnvg/dVQuaxTWfOO2oZnjvpJgL1ZnDH9iLjnfkKfw5rK3DPalJZUrer+LvnXl3nRpvo7Wcly1/WyEQYspMtQPQRG0Sqn4l7XyLX2+DLSRMYqKViLbvSx9cGijaUWAN8C9ZRQJAOBLpjHDHq/Ik26Fb7GRxxQJu45hJwuswIQ8xlqJS60QaMleLgKh5p14LrPbMA73Fc8zgOdYxHHbmRC2sDKoRH6XSkra74QoGrYiRoiDxmW0coTjyjQCzSswM3VtbW9YOtrpxS+7dbbJruXYbkTjRX32FKAIYOIqNDH5rQ46Zg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PfP3Dk2hyavkCQamkTg1STYWataViuiMQ9YOr2aGUfmTfDcGKlPvhuNE83TkjyAnVg4poMG/HOlGVvAoiJLmccrxIgu+y7PLl+8m+TQk+0LZvxtMkxvLIPIYHxuGc+fAT2XYMaS90OWHYy255lmg7RPmBDVs6K4uvpSHM22lQhY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TneRXGWJpTszCfuBgHsInnrljikrgZEF6mzL0wTH4wNmQxIqaSt+Q1MwEycnpb9O5OnZm6dOIjBALF0bOII/xwOffYewr1xkOguH6fLl0ICL9pNYv4Pz+YNWXW8gweLBHklWBJtqtnvQ6XHQ7/DPpW8+PLuM6/VsbseMVoMv5fVnL5b+QxjXvm6ak+gxrNIZo+yANC8p4s/cJB9lrHpEIsv8V1mptqafzcqWC7WrnG9OHDzl5X9W0gYcKRL7HnNa6PVK7pBBqOs5Zr/ztdBaoyVyrhmMLcv2blMY4eS9kK4Eu/nk3z8dBUzO1lpXjOQe+ABuP/de6SG1gb06InvHQg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4235)
`protect data_block
3AG4z3wAYOJEfeLw4SxghZcvBZJHp0qnkyEuyirBt+k1ooTZ1GOqX8Kedw/9nUbi6eHdTKK0J5TR
T3/UD0WoVBk8IalsxkSfRmcNNazawz/SHRDhGc1s8Hb7u40/OA3i/HrIbuCvDfOQZHSAFKvWdFTz
EbDAdc2L9TiiXJJGBA04b3EBhm6CxL0DaKIWrgJqPRklNbE8rbRy2GRmgapkckOcn+3E4YTUOaV7
JXSZXzea2kXu6LUjgvAjU3BcawCJIScHrS8hi78LTFfNpPsAFqIdBc0DSd3vrv1D8MLUvQLJaebw
KVb1F55FyrVCS1UNrU5cUZ+UqfWUZFpsvcVIcOtFkqsbGuQBMg74KqcA7zshUuYg+Nc3bPIDj5n+
KL3RxqKNoj145AXIkvqcGVIBO/Im/QAfy3j05iXSjXLiwpJUfuo2CPKYk78ac5FP2jgKxZtL0mVu
PpfHeiCgtd34m2+00vIQMQAb8HC0P5CBTemSxSMCI/ILwCxOO8hpy1wr4EZW3lD9AiUNgbzMdSMK
MERBII8NpZVVOs5RBXUvZ9xHsI4QJsXDv5D0OJrfj4F83vTfUw3SC3yCbCnOopkZ/ltixuJzVwIf
NzyLIT0V38VwN+4/y/NbVD1325/C5SnUPb02Fof+w0e0MJ7mAelWqSkEYWl71N5xUv32whUXnU7R
AwX5RIKPymMBkNRCVaYlicAH5YKgLjicqeK9JkQ/3t6TwIKZZy/p0UKZwgDEkh4DdDNJ3kFIPdYJ
lHw9cK4nKX/BmAgJPi95SZ/klIQyhKTvgPChuXuQHuvT0K3EYaMXGCcHKPHbFQst7X95LNLr1Z3T
ImoZMf4hYoYuS+xxu1xdya3fo374zSZ7BAQTZc5/4m52Yig9LIbL59hr56J3WOlnWRkG7B5E2yJb
pKklo7N3uqbd6eK1HI+fnLxcTjl/s2H+6g7atkoqALQ+46/4odrKoT/vr36Q5VysLK5IAbnSUNvh
Xt3CEI+SxJv8FMOXE0AibFWumca+P5YgHQPnae9BOyYjHF9aWu+WHh5yO6FZ2QT2yiUJ8rwnFdfl
v6qr97N1a0AfSZ6FJvX56Q5qec0wNGdECq/AUIAq3x5jbamDNiJjM0zsGInnwYYtfirGwjxh3PIY
/bR4P9zQtcqUsC7tPauHOV+Ia7PsfPRE0PXggnMhX4AKT/8d+BqKEJUnwXXVKIjAvX7ceKdaP9nq
UVdqpIIQbeMaU+iHB+OWZt5jNaiGqmeDEQjXo6EEKDgcNJbRi5H0maKLYA+OmbrI85DXSh363UAs
1YZaSAeePH8Nw8Wx2VrDhUruB+DcZl7zkITUJbtKZi6ZXIC3XloJ8+br5PpdJA/Wcn9zKIGAQqnL
Oo+mPre/xwlrTtefNw6KsNkEXiS00V+agnms64VbwUSEAFWHDxx9E1gOY7MbJBMxVbRGTKWPirPi
SoWTAdjDlJE+j1CBnGnFw7RWc261AOvbKpR+F2HC0NCVsidwMXSuMcwKGCOOzA1OKtbM4mODniIZ
qvWCtjA4jkZJ9N6nuW7cebH6aWxCUKGJr7xbJFxk2Eu9CuXvZ1zPAeBZhDQWecx7cRV+oMf6Gor3
jPdYb9bF+mIpKNPEuXhBNhVc1nJ0+MeuY9Pj4rUHu4fBw1G3yzEDWoassMxCa6RFrAJnfHg71Idh
iQHHUs174dv7ZyaTrgugQ88XP60iOS/mbCH8TvvjCee5GXR29dlbtMVhdrEoGxeYiLAOjg8QBA6q
XtJNZ+IIa5G7DoWO+hYkWEFolPsBSM6/eRKRSn32elOC2/aLpi3jf6XRiLcPWEC6hy/b5nEIa22Z
TAxD7KnCOJtmVJqD4OxML0eMGIqAT5nX6DkcVJw96IyPn4vfqklj7BwWGMmY/07NQWAeeGxEvXDi
LX6N2PnKM5DNtfnuwJgMJ4ARegSF4rvJHV6auDXzyz332jBXRWnyMOo35knFMuahyB53DuQUOITm
xH65XtQl2T3Zk/hy6M24njrdavM+hvXyzZw7xXr807ZjzjBQfF2sV1FuVsz01V1RFKXniHNyC9MV
r0as4VASnGxIsDxWyG8hejHYzOSoIyHPhWbTxi1XwRjPbrAT/S2JXlWFBpzIh1naNjWL8qL2uFpt
jd1kCqjJueffrc5A8veqdq/GegGsQSQKzc0DRbDb5MaulDRBQLxr3jxtO0CVftDlHFNtytS6s+nv
pOlFdfKYfwyyRo4gu78Y/JhVIclLGGHQzVNVytNLyauGgwSzyi9IwN8BV26LpaVWrEx/qdBUt8rZ
Xc0/kJ2s9l5YlPhEcW60Rs+u3PFDBBae65gBXr4Gu3vC7bwuYM467FSSnwPDAl3r7mThMIVsC1VW
2h3ZIeaVrJUqR2SsW68uv+qiQYNSlaDV7UNJ3GYTmvkylbQJKuliizvPrrKKIaeyH3LNzrJYKSI5
wc0F8ltBx5CFiQSK8Sr7iRAjCXqnkskqGU5ACIG3PQq0HqpKmqtLLoKxFAmGDn4RiGi6h06QwcKN
Izk18PYKXT4cOk3L13ZtuheR68r9q70H/ovynWFULZVbykXLzxBl90x7Y5L0n7rCaQ0vF+rUq/nt
xDE2KnB7Kg5WQr23xhhkjdbBw8i2cmTDqsOfyuPRrM/9WP3BzsC2QihhBALMMD4m3plaqNiyaSH8
7arn9JNnfl2555N4Mk1dNZlodG/ns6Rg0+7mbE+7zAEt1Qf+X/MBQjujSegTFFH6JJxVUptdr0lc
GpsslHj/mZaJho0vicNe4DQBRHzatLI6797CYXzesQLc2tkbDw6qlGO9BsE9o82OUBcpp9RKKURG
zoDdd9iWhpgzpfpCYhMgCJdGds5S58Z3XlGdTYkkXUl0qA/lujSVgo9vzf0hLToFUoEQHfORn099
UmNntsR9kWAICuejoQ1HqwBkssE6NAWjiR+ijOwhSvldBflNAlInbh68Dn3K430cqZsOTyi9s18X
/cs644SGGogUHN88htnX6H/6JHF+m3y4KM13d7Sg32FNBkNbI8Fq42+icg8jZxfzBzc6XfjOsXh9
iCfaOb3TzjoyM3L1UTkggb6ZVOw0t4heytTYWDteZEseQGbfYTfv/PPagFfjlvjIqdDENQcc72XZ
dKWZMp/OOqaRYEqnB60TZLbpNK59qgtGfvUR1eqRx6RuZYAk+x3frcdxpo0OjPja9iUR05t3Aso+
KNP7BeVjP/H1sB2f8LUqM8u2YyJkd82EUj/eLvZBgWlPSQl2ZahNemvqoADb8iwYtyzeANceK7dA
QU7BlD3wU2nIc3HvX7cDy2ejt4SyMVJJKj5mQ6cXPUid3IU4lQxckfluU6sZyyjVgTPbz+nepG77
XCAsknmsj0dGA5mQryXelFEGAPk+akacvoMO1n0wZyrCgMHGIiCAlb7M3/D+WPN1XxkQ570A4/tV
i4Oryfv76+oySOSRmGcj8Y2NQE7LULzE08voKBcsH5h6FMRhv+Fc8XJvhjF15qTlOVDyXnFalza2
yTb2h473mu4fhf+A0lNmpL4R0V1TTakCPf1bxAU0ppbtG4fjeiIGwnnpzqMSVvu/RKcc7oyoYIWu
zoxl+9aIxJ8Sdt8YxHNEB3kdu7tw5UeNBeaTRHatnZ/Pv+CTXYeybnH9muSytBmaPmJJoUFQBPV+
lTqhMXnBzujHk7na6ytng/GhyLUnXi914VOwAWuY342Gm9LKwdQubwdRM1glFxO6NdtCpQK3Fl2h
SLdm3xGlz3XuU/q01Et32QH4a4UnayPkA/FHa36eownGqsWzUk0DWc57GVwXIqgGv2LjlmXQ6CVH
aKXEToASd+ac0MpvKlpO954lU/+6r5qZpMSp6LqpomdDC34KOSGoKh6jO3oTyHo4JyWU12iXXXNV
T5aqIELHVSY04VCMtMVm6zUqcbDcQmqSNHvH9wIPls3H6GS8x9Q8Auu269Xt5fQ86vHgySwEppVB
DWL8KVGqd9/ZYsA1tpC8y+BZTzADdP5YOUjAPi+UJhcp8gXe7UD8i2U5ND5tkuLXaKQLo45WsUIe
zpwCnuJoUF3BuFhPmVwy/oI4CYFFGs9QJnbbGNwDlpanPAHBHcHlkG2Ty9QR4Ti5e7A8QAAyS3j4
a8jMdZQQiyLY5QcyHBuDj5xYGqTz9CM0hzM7ikR13+ZtRcAYf0noLjRz/u7hqxH9MvqPNW0UuiFo
/+Rw1OriXY1a9n5f13vSapd0dgLPEiwQtgtEdJri70oSskVGV8w1ojHoqDUrITPNjwyDiS+QMzcZ
hfLHdclyxs3h+1qQd493QtlpaAe4VL3TxYRq2rNBx8+jPPiIoHysz4957TQbllIYJ9yUscBCcJHF
6Tm4TOS69UAu2Ss/oOGNoEdcwMtOpnXIStJzMeu2KPxMYxusz1EVo8FJ/tHHz2qvXQczwgrD/OsU
nAnqKKJXmpr6FGY4qKO7wrOT5h9/g52xttnxkM8TNUWmvkNs47BAmAhBgGb/3Df7efosh1fqagfe
CR6FyK0JUmLRd2SgP9LoDS79GTQwThjLXz+msHx1pLpoToPILeGPQL3+UIfubdUSva1KKdzGSFZU
XIU6t4kxIoxDiYwCtSp6EqsTGGiDpNr+KNS2VptUs8zo4bMuYRBBRyWvskVAVvO83TXIZntFyyBX
2I1WvtGko7X6sUJvFzGuMeesSeQMNNA4YNkJPOtyD6oSDnWVvFE3mfadUYq/GM4Q9TN41AeyhjtK
Ppx9I6CqKCC0+91VQOW/TUmgU8qHUhMyrTTMLjyENTBnTrPGqkl4shOxi/ItBrxU09bpCoA4FXYd
fNkSkUSBrT5thSIJCzJA0azHg/s8936VH2oRt3W0fkv/oFyj5NQ2W5Bb5bMORhhN6Nwzo7z2NDOx
kEwp+4EHZDNw/JnlCWZf25Av4eETMIFtEM32KHk8wqUtmcxFx5PpKCv0Nh4+YwGK2yogvsjjKWec
8QrzIHEkgUHV7DxueY1YXKoHqxpongUDOEOiB3iV3fMUg1TgYDCGNGK16pycctdHpwMKKgg9QTF5
EC0rHE5R05e6NNIUXz71i3vhM8/rf4ersqy/q6r7QBYwbFwarKri4N69aUntAK6+jXosIYajNZLZ
xhQPe8saUwPcoR+ftWfCndmwgrPWFjXFxtGMo/UEjWPvrzyJ12HqVlVWyuZr6e4fBemP3swoUwt1
2fjTwUnMxpl3LqOODPppqF8gcCd09ibLtxkIMPxeI41yNTwc6RnstGqtg4q3zfnowPSAP6RUV3aX
blPB6Yeume0ks5aYM21RsXZ+KFR1ushjXCxTmvbym6peAdQwoEw5kaMoGeJ52Z4sy4apOEihEEj7
fr9FwYutCB7uWGy/ttreX1K//Es1V55o+N7Sa1h3gFpXeyN6jw2G2ZriR9UOvGg8LjoOEIaqO1/0
2BcErgmsvNqe6QVP+Xyq71a+PvuM+L0ie81TeqPtoLPsXVGYbPFQFQcD2NaKzVRiC+Mzt5VWcj57
SnDTzCnAI2GCAmE0eS/JgEuP1kfce4Zkvv4NPI2zT0YK6PRWBqEvLshph6aAMSzKHoFROh7S+w8u
Uk/iLrI+15sOQvqGGDCNICEs95ZKxSN18tuog6FXfBM5wpWEi4h5sk+eZ3KgLaQSquG6BELZdDRE
DXYcRY3jxZ2Mr+mpUYirgRKNHtV4nzmk+AfwanffmB9XzgtPEFw=
`protect end_protected
