`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fD2wpqTd8Rj85PHcI1OZzVwKo6nRDN3kzD1Q1jwdO4toID1uEbeXi0OlC/Abj314uvPs2v6xjd30U6kBBxWeRg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MwYFBfBdBUELaPAGh2AaPKXoAQGXpjg3DluQm/d7vbCLK38tzBgmFlURCJKDqgWheMpq8qcm/Yce8+MtXoqHGZ1uSiCk8bkz50c5p99qQtI1aA2XNsnFnwlio0hzJYsd/hZuBmg6ZvWJ8VmL9+deKg706GTnDNyUMeoBM1DBSVM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ww9NY677+QIWPFVblmPC8a0YywO6cQ1Mn3r6TbFtvloZ1flMhACCEIc5VPvYQ1HPZhjijp9NeQy21/EE1Td+x2kFeSlr3QxtV/OgNyYcazh7xvrww17M/xk+BiGjyTO6P+rsQAao7zuGa3qWtEPA9sM663Rq1LBRN/fMczs7PLdkXAQfbV9N3zB4kAd80f44ItvdtRHzyfj8RG8liGWQ2IBJow9LMyf+5u4WQSXGtqixbZC2Z50+0An9qjrb3xn8Ym5kGLLw1ljKfJgT/TWG0CJKr/ZPxP7sRZ8Ny4BNP40jVQ1DYkf+Xr/8Rx20BvpJsYE6Tvdtcjhg8Ri+6yHKAw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3Nn7057NakmeNaAw1COQdxYpJ+vtA7xczvonrRFuRF2Ub850YR7NVz4XR2lBHqPM8EMQ/gwrNttmCkUjypYth6UcDGiyRdrdCgm4QDtPrdXpSJPtq2MNPZlQm5CiW1iUtrNGzSwkVA2+08ekK46PIQ8/qSTcTicep0JWI402iMc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WEQNlfUEg8XSx76SXZuxZMljo/EfVRQihJIvJXG7cK9mHDHZ4mD187f8iT85tVYDvNUXmjY4rNkpn65NHDswH70rODjEmHJ2vJyRrESfcdTzvv81yvkkHGJFzpj/0JL6mO7w7b4sxVm3iSkvwzNJtVzvCS87yo/gmcQekWGw4vWwRW+mkZwmbzpI+dh7IqTtj8TyxytlrMo6d4sq015R5IhhiCNZCjgZK/CGCAup9xDo9Uc0tUzlmnWfrj9N8nyh0Jy8YNfbryFtoeASWQvMzmSWvKWbnXV7dKMC45hwGTsErGKsSI28xVLj2WZ2Ast/eIg5Btr4laGhfzWFgUmcVg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8296)
`protect data_block
Kg31LVsUE0jPIE7cJZVTPPLbS01pr444+ovpPA8jsdcRBx5ivIvH0ZE+JOacOLdrb+o2lZd1dcTd
j3At1OKS80LfQ02utcKXi/fomWIfnbhLfyG/eHTAZOXkgkevuuBFdjHt6c1SFjJifrOOTErXJOkJ
2YLUQcNhN20EjK3eNewlQ2IQcThyQfO3D1ivowVZT5CRaqmJTj0PDLjTSyBUGLRxs/MSYqKCd8U0
xiW03kLvP47a0zuVR/RuUP7aYq0RCRjpQxItLLOAretTim7FKG8QELVdEuyP5LjHYrT4rTEoT+VS
IGT7ZE2wVfZpKwuRLl+ln0akIj7hCHULJOu3dqFt7hiniX74J+vy4JfkvljWi1HttqakLwKyP2+T
jIrfJXzvHPViemT7OER4DrV3ijck4LabjGPyHFHnNrONaCjaeTgzP/91wlrLp8sFxBk0jdoIdEmS
fYLIoOgFmhrHsNdSyML1jzQwwZK0VTphiZWx6IX+4miBfH7sZRPl4chiZdCPllsI+PMvn2NhZAtf
E7R0wJ4tDf0wvW1lNWMWP6RI185xVZ3j68BHvzNby+LLHOzyJOZKPToft3pZtVPyzIZT3xWEreUY
sHorfSDWLF8baRPUyBSlQgWa4yQ5IuQpoHLNQcDu+O6VEBAwJ7hfi934AaPYV2RJshR5CrFjtNd8
jDiyq5dd5FhmL2WmNGioE8NoFW38Q81Fzar8dljosbB1Axjz0jcn+9ZS/iMrK9/3kRNjvDhvJiZJ
KggYo4YZmcto7j3XCx+nBIQyM1I/ZknMZxXjnl4FXD3LKIjDpH3skYTeMINcRfOrAGT17w9P6ZVq
PyovQhVRIFURGXdE2A3CCZQvRCwSU+XsxKXM8i5KaiuFgE3tSMkDfeZlkWKmrVgYfG9FA+kEO0mT
Xlj/loiMpVsCbAQwAj5h/p4NdYBaC6lAjFOeO8URUgfuIduTrxGZcK0fWl0UWwZBf6uhxnY+1mO5
T1PMJ5qz0CjdahKU+k5fl9E3/aMyL9daeX8bswrmWrLEJHY6Zzx5jk7Ah7jbQl3/721FXMrfDKbW
lCFCJx7+O5aFSg24LU1ObDT3AhTCKoMAY2e+YDOtkCANdmB0dhgj9wANtaKm5OzK1Dr9zrbsxAbF
4moSaD/NJFH/UBkh00dUnlHb5hFlCIPbGFNIMLJLISn8eDljig2Ny8CfWnd3hE7UsX2yxFDt013a
4Bifnk5T5sZd2Y0cXfeZpa1J0boqySCFlMl41H9GsB0RFQy4YmireHkfHG9VcjvHZafOsOXNYVCR
ihhzOGQw/XB1yDQXaoWaq5N7kX/9yWjMrhe/F3/nmQ/ckfMPmfvjl//x4Ko6vvxbvi8pisXTLvU8
wZrPqkrL09PIBHvJ27DjywA/j4FqEMfhiEuiV62UpT1Jg3OO1OUC6lB2PIg2B87r81/G1GxqkfoE
Hzp0xwWXJwys5KL3PwhfERLrz43NsS3AGZ2p0pRutegq0GCERHZX1ajCyWPP5mpRR4L1ShFXPvPR
+xHs7gNY98Yx+kk5pLkwXJvkeoC8mrxBpkmSB5hkLgEgfDypyL2nbpXq+aRYicoLGVtfI2FvWYOS
DickuNyd5vxjHKCrWTKcIejyZn3z0pzOowFNuqFQO5/+q3cCRFgX+I8vUHVA4Ycr27nEdOAJqnEn
zAi1Jpr7N8y/N/MquaAEiAx8kkr/SaMkhogP70qdKv15SMwSRUciqape0709g2XUrqz+L2sBp56R
dmuLRX5ZtVWAyEop7wQgZnQVBn8W2u22vbeOFxPUVZXiQTQA1cn6RPQ6HhMAp4eT25OIsEiZi/ja
FmuohTn2Ik180IEKRFYrMRqmsO8nCnmucXqbeZqBChm6WoXYfnGEkQUksUj0kcDZDJ/FbRtfYQdh
UzHXiNEajEa0FrzoeE0zjhCdeVQqrjXSNKCv1CTI0lq92PgeLp9uYYJQtAZKaSc/B1RbhcbKkZXn
cwM5nMRXJYUGATQ4M87pqmCFxUV0qou4waia0EtfkgevPCAwE6FhZw3tgmUSMRr02RAsnQW7zYUk
+aUdheBfADhC9SXVBVTParRYAfMm3+Obe6VH9Z/8MzYTubPidK1IpvH3Ug7+VWYN13JVYc357wls
IGEsZkvQSSGqWn7lKOXkLbxFaPv17I62pquMb+FEyyZG+nF1f/Hv3M0jnUI0qokSiKlTtourNEV9
ZD+RMM7ADagJBCOcWCL02upivVnTuxBIo0KzUKqthZkqq1MzF2//Y9j1ErW5t2SeDcCnMYSe1zJ2
BlyTAQ/KLDmevhtyIYJYsBvDfwjhGtR9pj2h/tl4LLNoFJQP5ebtBZWb+kCaj3frrZBM7G72TtnS
cjCsORdZdLa+BTK1QlNbb61QBt5yH9bJmhKs2AplIiFpnX7TFjk6ov3JX9G2pfOXt1YagKUT9uTR
rxG/fYn6Ui0ISs0meYPB7dJ32d8P9aBIHlAZytW0fJY/FymkvSMDR1oQiwvJFjq/gTKt7nv0/BUA
4UsC5TqUisBcOVOGN91v5rkLxDFBsz8PCRG9i8+8MMxsLlkF467L5POAEPXqrCqe/J+WRRCyiMkP
joIZIFPKvCodYE5r8q5UeSw/x7l/tTHkTxy1rgUlDlgx0RKfk6hdPTn4dVijtOJMeUa0peENlShK
bxcvWzbYuIivhpIWUNlSt67+frh/kcLA38t15IwUExIoP60Dm75pLY3ofep/dhqLvk99I+BP8e6J
KliqNK+2iLZWNBV+jB60dsFkG+thJCE/asGEzP5rxIt9PJwpCPEc1cYPDBczFd9Q6VzMRuj3ut16
5rTVRRw0SBlHD6tnoXkJ6zbLatwfYBB10AHjnFzw4zl1pq9wzRSIUE2lndqWuwXD8o17M4qF6lfP
P5GtCXgLXrH/C06bwzmcrI9lTEu1XW2UxC09aSgEhrX4KX2Krv1hArwgo09U/K0JylM+slkXkvHo
bf3FDC/EbSYyUyKsPgEOtuyRveDGNOXacHSm3nd2VbbxDkHPqTH84gG6QE5jtuTVUI7DuTp2r11h
tVMAD0dMCe0wSf7bZfsU1mUqGoFEQzL24FzfWSN98E49lKpZfv0EupLFw0uCKfEXY9s1cdUyVKxQ
08F2ADUJ2f+ltxzxixbtry6l3kvPLUgTx85wE69ak6BpqndPlZURLRriwZNu1iO0Kk/sXI+y94SM
oFGm1LI+fu5gdYWmn0Whv9qqnT41Bwy4T8Rxbl4n+pD+rN5LVT1FiavRczceOSeKVFypk2Pwmlr3
nr/7DdiX6Jzp5KqBr1TzbYAMcS5xHrXLuZXw9KPoOSx+T6BYswUNDCt624rl0an3G2KaKINaC6KB
iA3VpTDw+aT04L6hN6u1GwH0dyXk5ykB2RCWsygwUAQ211TLaGZdTdlsoVKxoXaGC03CTJoLz6QU
aGpQ8WIx/DtxCRSY/UCTaC7hWP+fmsJm1sbvnDW1uJS+dGbfwcssaASCpD+1Msb3ibzZA20uwo/7
42Q5wzYGdX2HLMuMi2mr6xk+OWVfGVz/axvwAn0dXotxpkFsUnMYBx3sRnqBEI1sXqw2Pheep+0d
dt5kXxKLVbc8c3ajDrHfrHUMACuuoFf4VfHpPHGxxSAwjGZFyXeiI9jfWjCHipA5P3L1ojxQ5eYi
dugMu7LJvCti3HbQMDZbZH1cFxOIDbsUEXwfhVLHDlNUg0cM8QivcO+92qoIlNB1MzYqnA4AcTGL
YVvK2SYMs4B+1hzwQmxPvSOX9P/fM+c4f47eb2Hczk3CKIHqx+9TMBTgNITSHRrwP8v1+9sWH2Wi
rMUExS1uEn+tnXRpScy1B9Ld+UT6/Wkf88jtdkrPjV34FK3zs50n6QQzUGXkaTm0yQjM+6ur9UGJ
Od3vaCGbYcL9zEhpg/2UN8yLfDTecaGr4uOG3M5+LwiGyQbkK7sowrw6owhy7scBVnyNuQdMCX4k
7NfabOmebFR6WbFT9bCg5+4RlIY9bwGdWxmxoTd1LAb/sn7q1UXrQGi0ayv14WZlC8+fbyKLU3Nw
H5NxiRXImBAepH86dUrBQgGxPNI79We3oYtV8R1Gss1E4fC8Gv5U3stxwJZX/BHhJQvPDHPglMvV
rohWiTrRTk/smOoM0ZZ7D1V5ZGxH+0UqsDOK38XhZohlOcyfxpQ/DKxq+WdApbTICXZ22s+jTuEP
wDCZzdIxVQb2OnwKydlTUSWolh60iHdlVR7kCNdS42OTr1k4EfcOSo9TPMxa6KGh8wPTlilPYe1n
ES5M+weHFNZClxqRoDlkv095mPY+onhTTeMqIHdYWLRDeR9b8QsNiKgk5G/2aqqizBK5kcuj5yL7
i4k61gcbovCqF/NKLjqh+euaQkcTksb2HSn4RZPEJ2YCn9sZjJeFthec92pC0WAQy/kG6i6tQOkG
8oRcz3Jm1fSy1fsapulRn1AFWYzKdusR5wMD12I7DXidvV4hmFw1FEAy5eLu/3wC2Z0zTOj0O/2T
ePcMgo46b7jBtGUUmRkxZLqOVWUBe0nHoAiRy5LY+T/BpU/6oiDOPGVdqP3YzYU/DtYSbU5L6ncf
3e8waAFSzAhX2BsfKC/8htUCZeW1xDLywUOrxj/zfjwj5GRFzNczlkj5jqKz8QIYR5/JvmyKuXiy
tgG/qGrjZ/DRxv4VyJH72bexw3xhXl0N/0nFjNjUu7t1o0c0ZrGdqd4mQhtDitRDM/5wKTaC1f7X
wWKwzuHNnMY5pxkcgDUFLha6MXmQ6jgLW+zt7uLxRd03k0SrM+8Ritou2JDM2BeEG++ByxyfO07R
ajpiJcVL6nKypHJe+m/y8M5zAQtPxHPZj0fq5MrHfcDvJ5jG7FuNwnWQtIACkJL4vBkcNWL03BOr
AEZN0ewKFk6TOInNKmjFOaWLNohN8Eb1VITJe0/9ysxSdNAlMHOSfvxkmL5xDbUeZjoyClC4kRFH
Jc9Qnz1sBJrrXIOHur1b2NTy/RvyficwNRRG3P6D98NOxNGDxd0SrdFqxvn9feIr/RNoBwr7Twho
kQ9Ok6Rwuljf8DkcOdMCfBmWbRoeA5eQUWykaL8zVqAqA7NMRKJBCOZgigoZ4bBG69/PAx3Mlnph
FuSV+ClxbKXGYBo2b1gWetIn+4aTzQhYORJ1R9k9eBlL+cATBWf1ku4DTCFVeq+pYh5c3UByHvSE
y5TIg5rYpALFiRk+5JDe0W2Yv+/nQ3t8HqhjHeWTWQzKbiG8/zd1WGX4dMUuVttlaTDJ3hcE8BTZ
zD8wPZ6+rcNLT3UGl5RMoUgBpgrMqMsVhSVICkoA6Jq6Gdl9wRU8VeIO6YaGBujCEBj9GEHnFah4
+ufE3m1TfsjL6wEROC3NzFbGkoIjLTRbTQL6f+O8NOv86z4kH0lAQE+TaOPWFihWHUWb5H6LMpiE
ye86i0RbS3KPsr10+FXQM6pIsHKcFlYdrLtopLi24F5d00un0mAIa/5z08Mp8tx8BlouWG/QtO/g
YleZocIM7wHvuD63qzAfP0fqepaGdG1H/YvcelBZHnra56O8RbA2lryyLIclkHngDVICu/KAdODU
eUH33Zf/5PbLw6EWi3zpaQtoXpQmWZ0pTVISIeNDTDeSRSUTixvS/GiUvk2iZVb731LaXAL/XaJV
uHHjBbpzbYZdeNpbsO++hszDEXrCTBBIOx8s0byWEe3+7kBa6jsbohJEOPLA9nY2GxYxsJlJ+U97
vR6x2kXsjpdcPXh54bbnFqiHyje7DAZs97kopcu1lcoCOdBdvAQRjBSzV8e4ae0nRpMhGkIAMrya
vJbg4GkKZwVYu220j0K3ROKNKcWtOnX7uHvsI8BpabPeuTI74j3MhNjy11emM5OP70i+oW/l79ep
8LbSeDefCm9R79pJ0eORCZXh6lUmCxvNApZ9g/slqTXTTDzUbiJMkLWAaQZfAmmfEB2M3RJD+ueN
ZLcOjAieXk0hF7YtNIRM4nTa4PCPXKC7bx9LOx3XDZ53WIeYxQNyeErh0QllvjuI/+wrJbOuqY9r
BIK7vvCfKrY77bkvGObuUlv0e4W9GFWecc9APw5QMYNH3hRZpBiBGvO6G2Zfgk4URegHvO2vfHIC
UitIvbo9/KL+Ig/lmEjycs1nzhamWM4QPr60y4hvObeSzMd20pkHaACAIr7EI9c6LhLMJO8Pb5m9
pkaCc7IjbgXwWQdI5o8RbYFcWfpoDtgeEdAESE37M0OK9NoOLC8WOQSTzTaMnV9Y2gmAJ0ywR68k
XFHtDL2cKuwJakyiAquJfsbb2ag/dS7567aiDxLiNavFOcSru9RJW0MDIyua+g36QiKJ2l5qlFuU
u2Zd8HfW4zJPO1HfkscVD4lEEQOzmbWVDJT6FLOrQcHQ/S/t6bgpNy1V4fAUH4SwP42d2kHJRRZt
GnoFuHcRCY/Jo0ri0WR81/ZIgieSIzbWH6hedRMfuy57KUqdW9pFl+gLreWhnctsmLLpytxCvQ31
wtJyZ+2Q6UCx/EtMnrWYwsZNYXv0GxQQI95npstn1gBznx6MhrOP+SUllaCsU75xk3SI7CeqTeS8
BeC6Jjeg7SbaMLaa2Hu6LWHAWBGhlE1+E7ZBQwYawXuloKAm+XtQegy27oPrEUaeyYybnwVXqi0R
ggO3iamHLvUhzadpTptaK2AMcBk3z2+liNxq9Ett7xnIW+7tPsMxI0GhZnLlyMzC8BpWQnh9jhxc
D+ul9xMK5IszpM1Lw52LoUp8r3/vQdEfGivSEyZglkyAZ1j2X3s4B/sWZH114flGKLftuDlG6g/F
zH8gtTheqOzaQFVCGm6PgyRXACzhZ/W16iBe5xND/4VcR6yFd4i0UwOWiLBh6mB5yMg4XP/kzZQp
VP9ry3HjgMt9d/44G3Dqb+1JQlh7M3qmpY4o42P5Y9bP9vCVENKzabZYaSVaGr3otBziVMePIiPz
ho9x4kPtMAmj5MvvAp5pmQIA/JI2OprFx/hfqhY3K5uKRIfmY8mGY98BHf7XPD00bWjWwKj+y/Bw
cwpyNAzSXo/TT2FF4SULq47V9kktWCS4ylf4jNTLqNnYumY52mAXPbCXYly3Od6P4Nq+NuQBA2sq
KNmKnFDjZCVtn0WwMcMQHnco+IvPXXAlOFG2lPhjRTOndKwBQKSLDXHML9X8INafMxcoCpmvPJ2g
uVDQo+eVZSNItZBVH7XySm76Z9lqJyeMk0z4AFVGgtPEPEMd54V3uvTK9UsjGo9WZbyDvS6xD5iR
ay1oRR2JYcHG8Ck1kEIK+t7/X7j0GY4rXx/53Y8sj/ciMuZj2i9IsbYztfP69mT6JBPQ+ck2pta1
los77+Ph03U1jOBXXm/jDSBfF1nUHMZMj3iVGZv5Cbi52PT1hnBwWRb7JhrfCPDPFcb6dG/y1TVf
MI+VXXTjZ2fQIv7e93dIzA/fE5kRAU8XOipBVVuaXo4t2V85wCkEzg11QeFzQsEipYjzrEy2ZR+7
zjPxLlDG3PWJ6pKAYE3nvgPEam5/HJYvRG88JEgK9KeFwDo5JZ1DuxXqMdYOMvxqzIQIbVgGsRdG
yXab8cun9PmRa62i1PK0Z4/8UgNhtd5mNteV+ldsr5QvcFwjROAkmr3ca3k2pHRKlsxs1p6UO2ji
9C1n9wH6eOyT4RT22KEMN3/Ef7/scoFwtC8fLAcVVkyDkHYcxL8kszdqSoh3acmPXuF7/Vb9DAf0
UdJrLgd6h9FvADS2VAGnhXVwfrOSeW3D4kfhcunR3Tk6ieLCSK6f3YZQj1U6UvilArINy8QIjzvR
Q75WiJ1WXrz8Qao++cProbZ/J9uO4LW5iVim6kLABhldpyXp2JUhfKatuqgbXyd9Poo0kM4U9jtL
EL6uEluezh7+uxOYLaD60pKEtzySnBntf0+4OB1p0ptXjwg/EPkd4WtMq5mGsIJWhf87OntHeRvm
Md2t6MhbjhiQWZe3HGn+l8U1sjb7YzhyRijfJlYYGFLbyVXw1IzstrYbADapjYRG4NzMK+gsLYkX
H1n/Sv2ILYHeVMlcaw1CKTbHQwqzSGmh/4JbdBUXqxGcGlD94G5IMaNh0LSf3DWvmqrAvkk/I5iI
LW5fG0GRkVQWboVxhqwhpB7jgLZBrK70Q9gOQ2A4bEh57FUEXE4M8yi2QBnMbyJfTy1Ad8JDxwvH
tCdGxB9FZF51iVecRJ2BjMjVR4oMdxZNgJaALTKtwjPxL2lJ8O7Ln9KLj8fIl58IUTSdTcEWB5PR
NYQ9m8GH1vE0HErsIT6/qx4fL3xaZNMAY1xDOUNirwAe4pHzWF1DB8whtzAErXebusLNquBcNwHq
SIdBKOczssKeJGwRszUiocX4ummmooJqqQjLtRNVBg6ixjYnmsV1kZf0NuQn8IoEimbh5VcbXYtD
+xLINelO8Si0ZCN64Y5rhAk8QUmvK0XgiLrVdg6k+YLa21aHfwZY14gmzWOx/avzQZECZLuqgrHF
6gb/nB2Vjx31w2J/aiwKMj4cFL4W53aSsWqbhyg7/erkd68a2hJJ5fM8PQX103NBcgxcuA8Mbz8n
qxDbLvGUvvSdvw4gTCZLEag9Q0qUT5Ab8Ma85kvZ23xR7tPOoqXPpj6CV3Ql2PhMxuZLa8oO2pMc
hKBJxyXGo1T0uF0zkJDqnUGhVR5MCcUxiDAG9RFZm/UbDpDNvx/m2atzDgmcenz/Cmw4BxNmWJAn
vfK1K15h65jR1SrXeyZPeJFIi7PyqetA1ff25o3kg9LJlFLReVbh6HXpprfACZFuNwelXN/jf+oi
7ZKuZgwtq+8yc37xSXW79BtlKhyOkdLhG65dkG5cXpxhDZUunFCCItdDX3cX5DNa9vU3lSp//L9M
0oh5NB/EvgL7FxVRojvhvLiPTMcvTuwUg3fZIDf351ClKR7Lnk7UzBRY+KPGz6LyTlouxG/tYq2v
e5aLmXzS0OdNaC1514CfW/IPCeRz6Vsx0MUo1/tqy9QGmjxanr7qe5tkVTCaoBc1jH/5RE+qfsXS
0s/3LKkAhMbpJSCcHVtt5OEDUbIcvHiXGUFr88g+7VPq+UzweUKKllVP4BhYCv1VZyeRE55Msa41
gclmZ6iUeGtxsaoiEBJf73+m+bI5wCxReBLEEP9Gdb9/YmLcihi+z6Xxz+fhoifrrWddFVSRlHtc
DIHrNCPtH9YsQqMBD3P6Pgwfy2yyIDqw2SI9TOAyvpQyhGdzEA5+M7JI8UqlkNCRngt7dbGx0wKe
NJIA4BYN8dFDZ7JVGuwZgkvpQYKk1c6Ye3OnhfdFw0NzNcMls25t10snyVW/wSXu2U6oExnFS3HF
505lbWsR5BR8qcYi2dW+sZbohta/YXmZIe4QqvMLO/YR6RZWSQYmEf9yliRMmX/0WXGY/PxDMf5Z
/fKpmu1fvKRRltJbQUNuYyNWcQRpb8DcZRSqBoerpY2yCOVI5ViAw0ivZxC39F9iyBenyGk3yVMd
Lf4A4KMTqnQ1WQxeunj+vambadBjxUXykN8Xh2E3AawUNJWU/mSWRxw5dTdE2yWhrP8j0B+Mje+a
doQa8ha9heM1k6j9Fgg/4t5QvcFrXOwhDic3Np9smM9Al8bZAzu2sTZW6/Rm1LcQGlAbAhadnLhV
3lAWHr4iF3S5zJgMZBRv1egsrVSG8nf/D/nPebvDyh9ZrwO/koIuD2vttB6N6ugaxMpfWSqE+qrr
ii2J7slQwuBhKQ8EYWHhPnpojjV6hgWHnk4oXeXfSG2ZcgIAfFVMyPrrF6GMr+YjnIfg12Joyjrw
mrSp5A/XatEaJOwt2sZEcfBAfdM+d4aJwCtNjeDAuw5tSqw0VAvLT3bYGggjuW2JuS7uRPXdNld2
ZjcDzMDF36/5zqQiHt2ngM79PdeGCaig39DuATM5sD6Q2GhB3R0dx2oCwWfadZ8YGmyz4/WwnYcY
gKuFLTD2s/ISCC8frao15F3iNIAOvEvKEMXy/dVn5crzmrEiAXxZSUS4tiXLwsvEoKLjfgyxpmHB
hMWFMKZfI4AFEm8vlfwj9RaS6s8lQStfpCrG0B88DN4OsC58RQ7aXxC6A6RwgAS7Ttv7Lgb2LTxT
+D0d91o57ORC3cVFELE8eT+nlsB61tgaiWknwyMso0ucEGWLt0SWSW5YfvGKUV0wLbl4C4Be4JgZ
aMGPCCmgNz7Wbi7257zBHF4EsZ49YWJ28ly1xkhk3picv8e8BouVhHXxPfnZzYiv45PQl7mDfWud
Z57KLVdutSQ9JT+TnKdwofJlEkAyBK1Y0DW+oxh73ceEuudMP2vgf3Zc75K3kMOvZhYgxi8B8Qvy
ibO240TVbHIX2PZW/Io8iX35I7cXIpGq39gpz9YYxEUVr8NDn2uk+42EKT6JJxmEjVLOULErbnOJ
NaRtDhT5E7W/NN0t3eAecOjt0zrCeHRqqv7WR8rREI1py5RvtLHu8Ym3mNUyzSBmJr4QULUDXgjx
+xIwbgR2ymCUZkZS3tNv66SgNg45t6L+X5KbpptkKw5g4CVElpD3V5CoMf0EW/PNEu0zezeryVdv
LxggBmDNFpZl8ePrZxJwCWzTC+oQvNjn8CTl5b8vhzXbPj7GNrGIQrwmSfbKDy1xRJMfy9sm+ftJ
IuBS3jN0q4BevcAXTclBmodPFJbV4LnZUZAIHVHczNOqiWDuvIE3kUzioNXzqfpjiwTFL6sBLEjJ
yVy8zNx+id8nqh7qAjVbToNccb0EEN8uniqNlUip4ufCCLcRRYMgBUus9MYBpxqkGHlLfsvYCYT9
JMiQO7FZM+w9dle4gSi3UTAzdk805V7HcHEGpiIH89Ep2+CNBiQMhxcM7+RijcEDkJGvEAvk3J6Q
nduejox9ANYAixVUmehsMek+fv7fttvtjEWlZCIHiBQEiDTylHbAc45EA5XPrY6vUvz2ACIX262k
8uQDdTFVuwv9v+V9NeMrTFxHCRw0PhqY90x+h55Az17aORLkyix+BxzRVZc9A61wfQ+MyQEmOr5E
xyZ82X4SOiPgZdeyy7NmxFqx3sKxVcj6DKhOFgAnmMRPr2MOLR0ppN/PFGUqBMz5G89j8zfGnD9E
GCwT9U9/s0rHdR3w8gBeYrdNaIZ1cRUg3n17rwBJqNnHmxestycNQCPMDmtLf0gB
Z6D6VVlTNA==
`protect end_protected
