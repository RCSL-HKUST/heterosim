`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WGdAYId1gWrvV8rZuLJwI3jfs5VVYnbSuaa1R8irDJRr1wMwRIy4KJGHRMPX4rlJdfwTGL0LY6qnuwDoEhuBoA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H9C60+dosOXRRqlk185P7CWWrru6rci9n++AA8nrNC1Ks0K6Z6oa+WUGyMCxmM4oCfkTvtkqx3GAd5yLX4CRRZIeD7iK4wwjd8OZhiHGjQBBEJgF6WmAG7QbTmURIanLmP5W9vPuFNlzBuFcBjGhbioc1HEpEBexMknBZ2ZXdZ4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XFGjbElBezqW8PQJLk2t8PtWqAlPIXA1CGVtoHBBrlFtjRYi8gVzN4fRcR9Sxb/b7QExufqfl+g90fjJkr/VX+MzmeKWQN443v+kf56BFuJoRQo6hRg2c2fI2xud6INThWhHcWialdQw+dToo/SrJbXsQ3/KrAR3Y5gocJpG9HE/EyukWPL2BsHRQNHvwSUyacO7190PSHQgApFwtgCL4zctj9SN1Cc4ac367n6v4xbjCz99MuuoChc58Dw3B/eihkjh79ASZ8xPmGRKNDCPtP5TIeORoqjLtQ4jn5vSQZBziX/y6yv7HNlasn2o32fljvvtamJXG3ht9hbSs/aPnA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gDT63fPiZGOFux8QsbHX22f/5P+bQJkVZu60itL9R92otSrDjw3k1shurx0lf5NA/dLKEINUjAmEyeb4+44Sa6r5Lmry0F7Z2wOh4uxK++z8YTntr2nSzc3fdAlayxV+rdDQqzt4CRq8BL7SRjbzQngvazbn3UB3R37hVgzMibw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TeBnNRoAqdflRLY7vG7V1MiG2BUjg4thjjsxMtt9SSaqk6fNEd+MEjeZysD5kAw8lUF5rK2bfu3Af+loakGY4lNcwWfErLCU9ZQRcQ6xVVXQ91T+C74GRabJ0hBAyE2eE1V/IQ1rqpCRWJEQAoU7d1ay44gAo/SAx91HR/jus6KQ6AZUTxFzyi2rd0V+wcMEy8G8nsBDGAzTzo4Ypd/4lzGSd2+91rcTg/mPJvPwgeGC7ixF9MwDzyCiB6Uh3Zt1dJlY48xIp7mYdpFrl9NuZozk5xXMkO0ywoMAHYWRWipyHHVWZ2mU/NyNGByVUP9XmegPMROu3uvkg6zkXxRMqg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4230)
`protect data_block
dW21+OeBEsjR5rRmtfqiGYvN1jXWqaCI8g6EQTgVo2MO37Wjx228l0691d+J5lF15ChQilj5+3jh
VEaBUpLcohLLG1DKc8ASTgX7BSk7L80shkbtd6EDZjQ9gplnJHttUy0xPakfL0ivZkDwE5paOVVH
EA2NqXC7v/Gdir8I7RuvBy9jXmlUlNxpOj4rdybyY7/sJfndreHsJElU8KWozHw6/oaxtfCzKBtk
un58L/7HLBtViaoPl+KAYqooZbUOal87dSUzZhU3AA9+1nMdxRMWVkx6He9Hl6/X0bdK+ZkvsNgX
2n+X1dBB+ulWyV/Wnp1B9dXadVlP9Lmo2kQfUTfBXGcCdMJj/vL0A9OsyorFcwnTTFsWvr35nmsH
Sro9YBJMa9vKCrPpfDMYNK1AFYM7IxSMezSnyuILuAqVDz80mcXcBtLkYuqnQmokYrvRSn/27IWM
uE5fdSkBtYi/uXypMbuX78wr54hDSCFTlOURc4ekyj8dRb2g2LSqWVvz7IsJBJdegmLRmWg6g8pf
vlQSIWkyay3E1VSekaMSKIz59iLa3aztksTr36wiFXR1134z5gFtXey+MkxYO1eud8tevP6sAfPu
wlmOk3VerYNWlSbTqoI4wXPJWQXZEhqiofAPo0YeiZaFPHkGE2N4wUnEpwbIdHYrJmKAezmZpAoe
RrtbWeqcnIwnIXFFuQhT925NyUmdtsL0wiprgbmG4VJRkz1du1wLYtTP0wf08fuw3p++w0fRecaY
2RKJjD66PCqL47Y+d9yxL6TKrqg6QGcuSYcUUltFrYzDLXJsewaGXIDv7PHsXb6KPn5DLl0eKwi0
gknT0gQFSg3V92PMIx8ZxXWzPFiF3iKuG8IsvTYIWqAuJbsYrchWi6uwu2+rtRMhNrsuW1oxQoGf
Dt77Vnsp+Bh0Kz4kz1pa4lSgzORhWrMCDsxcZIAZz6xHsU/IFzYin88eh2eLxG3QNznXIF4p+dIH
PwVmVGKyECAtoNL7vuVRvrSRmDaAPMQFk5Yv5NMzZUNzHRwBwRDulEfojgsy42lPZQwvpcS1B9yo
3Tt/2ulA6EhNImBOTEGxQFZy7BSdOSZkjZQW3YbtKvBzZs2Kl61rGZJmpHg/eLtE3YvKo7VLP5pZ
el3i96fgH+bSjUPDjapomw79MZX8d+xLWLtZNuiViHNp400gYOkX/tw6+Fv1qUKNsQCK/94PARDz
dIXHc9ftqNX/wcKpjimu9Owt/wZ/r4RbYsLidTAuORWDyoOaO35llhsJ4HJxJnz9WVKftx4BGxm9
KUiiROW5IxOr3kN8x3NwpYAk18o3nHR/8AGmboeWDpGUz/740019PfcMhvfff0tAbOXzPFWOxAJ/
a81k1cgJWY2Zcz/ON8ZpzTSDWrTOrLHnkJIgkb5wpFf8arXuZU6mqjQAFy3MeL7/Zg26v5mib880
J4BfgYz+p4Bu18UZ50fprPpVXnz1sutbWmAA6qweMtlmiOVpX+NJX2fQbebe0QwHVaTgITmwu6YE
rWAlAECuAYsHXpJ/9lJXaJ0n7N8AGS0SW5qmQnD2wR288cqoECruRPUvTr9sqllpH5XX4d/9KZ8r
iTRMbJaUneXiCCayoZtPPCv8sneB6QWe0VGOKvVnhUCWpxhXuz4lt5ZaC1ogqB0SurMoZNTeVpG1
Nel648jUHfaTkOEgtlVXUkI5fnHRffhzsUU7SLZooqevtrnFgmMn5BOhkNNP8Io+6Kw/IMQQTE+D
Ybm4qIsUTKXmJSktW4I8rTwRXwm39k8ZfP+ktoX7d56rNVJFZ6SdDailP36ibeSYAFeSjFcIgxzP
RVCjGmzKbsFhboVd4SRNiTNzzC7ZjlJqDUiusqbENb2gLbrLsLSPpK6Om7LRJtxCOlfps+zdBsK4
o0kPjVAZRHqZ2KkeDtjxdUlIZdJ7PAR3J5r/RZ48oFtIDvP4P1fs4lZ7HROoWN3XJbro6+DsfjcO
bz5FNmUDRJdkKNSxAt5/TIZRS77lc2vfKauHydhRJhpCAcKl5c5VqJurYxAhMczaHI5M4TomAm/c
9QwPtbPjIR61+vXsM829p2J0GGg1l2CVRuiLYnx9okoDUy41RJzObDDnfh6txl0gavoWaRCoToPO
SeUVL5P6t15Lpoa/+otN/lzfV7lqY0PZLN7es9j4E8DUKcGqDzBOOwLXNzb1ByYXYgBDF8ZXyjfj
VkDu4HZjCImZwt/+q0OEiKSwLA+wDWNNH3P/4eTpe07v5S/4nBYQhtdQsXcyn/4H9Hx7moI6L8OW
ueY4T7OIRedUcp+9pHP02VEZnp4zJ4d6rjJ9gANYjEHjyHMlYGGVZQPTJcsm8mYmjVD6Mf6mYLtU
7a6l0GXEd069acZXyAEQrZhU//lI0rOQuob2kbeazPjhHiaElLwUE8GBNe3BPtomFr3aV/HK+yYu
VutydlOwxdMpBH5xm4IuwhjogxPsqexIYBQJob+5ogwaQS3fXX1Il0YqI7nNKOpM41GNcNps+2MM
u5OxiDr844cHgPmcmoza/5GR5gy5Z4b5Z1p8B4LNcGbo0/rW5YuoTwkuX1CrWAkxbmroMaBMMY6y
xot4qjkOGc8EpST11QtRbtJ/gH+tkIW40tPlZVfPtZLos/brpPkpCKHwcH4mI5bskxXUHhlalQzx
xnsTzq4lfD46hxXqeXdoqVpRkFUmZJa3FIz9gxh0V2hNyNrxcmVGnvhr8cDQ4Mr1q5EDf8ALfC8O
A19OgWTPa52INbVPtDBKF8B5EiajLhcueWDTdlvyZu3Q+36k0miZFRFsYgTyHN8Zp2Wo1n7RFJbo
BFRrMsOLAshnncNquxbbJ/SNwomJgzloUJgr5K5A6FVBx+jP5AFyFJrFmbIKNr2XWKsKfvBly5Qs
JSdeYfLB8BtYboJRbh3C4JJ2M1DmmGSG5X4c6/2VWphEciwnL8lBlF0FwrIg78HOYKbZPdbtMQLb
5hxgwTQGOxZV1NerHpjKnvkzXtVoQozw0Yu3ce0WGtCHNI70zMaLaSjslHnQdBr0CjCPzQSYbbUv
I92h4TOsCj2WfHC8ZTUgxAh+pNzDCAO7TX5CXrWQIvRdg32olJCd3sRVNiFoM/V5nWWbPZuNcHVZ
x9Jxxp7vwXHi79gBtE88f1u1NR/HLdOeW5uaNnS1vDl+tEl1bmAcwRniaYnRh5wj2t6WbH5Q/nkO
ZbaOOKpInWoZs7YXE+qzmi3jB8NwssWwbjx9gsivqaEOc7ymeSjyYtl/Oyg4gnrucHufqtgZbKX1
AwCG3ohoNbgTSrHe6LYW4r6d5zsgFVlxRoIBHnTNhOt1zmYBwyajLhFZB+lJuPmwt2vmd3w3mq4D
X08P+XYPpqqZGs1e78u16+6T7jwF/d0F0Qr97NdqrjmiSItqQgDuRy7KCATr7IuJnnXzDuzHESi5
SyQxuaXv0hFNDPDxps34NKXdsPOc6yROcsxjxV4iPU0uG2hO4UEm1CdcY9Qh0PnAodGoqmgPs67p
Msshsdcld9XGeGPMgg96XRcDSKUiwgY61KFHGAk9F1JC0rqdhZrd1nI48Hse+8on6RJTvXIHVhqe
7aDarLscilw7/xnBC8XBZHrV5Zj4AQzNl9PzUlOuOsf1ereQ8JQ4sczExXiwbkkPSgdViqboWWZf
VCWL9MZ3GGztRsyCWW0fMxkd2s54Wzdhq+2duSRJGBUsG183mN1cNLYRnVmTGTYm+7L7nutMCOF2
k1rSuO9tvvGJ+eRCcuxPN/pCJGCksZLTzraKzWgtAKKyNh3RTq4YRitYfUFQzSpVKiniEmwkcXvu
rku7ZpZ/6iLQMd4NQtf9vZb2pVcUwq6Sl/80NV0PxFAjWq8kyD2U2FNN25LPbL8cdSR1AtSIUP2r
k61DG+Jmm/zUEic1A7vzImWEIQ5I3rY4g6kHLdoI1rw5HAbO2Zm65E1FbimWQ9OhPSxHryJycHDB
Hc69ZoOhaJHV5v2hEHmKXl0T2FWPnn3aDQ4K917QIFEhx3lIeOL1C7kV9mEmWllK3MGzW98TJZVj
WFRCYkQQh9vPKE7RCypaNBGy10E7Kv+Xp4qxCjyGTiGhKLAdwBLK54oPRNC/7cdAAD7UNJELwy6S
SdiJC+7hz4ZsGvnM0LN9UcsYdmydhx2Zsxe+/Qkd4h6nOYIYf61ZBZvsiPxu5nJX8ZhdJ+xE4EmH
bK03T58GDXfuQ3XWGGVIWYPj+0GvxH/3tE60SXaj3elzAYYjxRPtSEp6/udPR5+JSOepvSdGZ5uA
+8KJKbjJ7BuUE7xTIjFUocawN/HwwSvNCb31G4LIu442FfyqSqKdkL4CFJInx5JvdR4xNOv789rU
4aZ3cJjS5p65/5Q3/mNHGEvKgYPEnNmahdyOT8SpBykLjzuhS8UXmTB4ga7TDaOyYLYal07Cfr4T
koErMfzU8l+FlTMPgeYMFnyZAvNy2nFCRsOkKl/OPqUBLG2tDS5LJVMnKoZ3vVexjdW/FX2VIy+w
O1q88ns5Hmz1tQloVkvmliloXk/4lTgkT8fAtRZcsPRvGBXegCv+TyyQ5VtGZrYaDOZJKjw7OxUY
jWF5lRPaI6n5V1qVHMKDvwkguNu/IfQvP+21xhKst8m+35enZgdUoZcrg8h934+LINRqAEBvMp6D
/cdDGiXORAkEfHzEUXYU28B9dpZi8Jegl6evL/vmtYwLDAVFiDsG9vYEx2ChTnIhggID+8FYgqGq
4wov8W4liPFY5zTXzx1vWSaJEPvh/oBJ8BqNM43va6SR3fH+PG2/XUK0XEh4BN8J6uGgpLGfQ6lq
J9XjjZ0G5n5pNclTy5L3OJYrKsG1fp2LELVkWXkkiodhR+irsMtwjT1rCFmb++lNU9YPUvKo1L/U
v44qy63ZAC2xJfdtQnOuSALcZTpXjJ+mL3JE+jlgXO+TNUS0c+rThwpJ1qGWKNh4sJoArTxjLFWD
mukIDP9TT2FXlnKF0iGi+oDtxFrO1NtLkgfI9tuPs4dLTVKgleUsoM8Ktodl4FCe+9Q4BEeKb6sb
6ULi9u9aXY7Uudjw5JyuLXC+PBsQfHL8n6OUXXQ0nx6e+baGY7fFcfZVIgtWEhg00/f7MghIX8zz
F/sFfY95nNv5qJrt15MjWk6f0zh348tssqWDy2zNpuolsxK/vODcDpPGjkak4Cyq2VyB0jXqBOS9
BigSCKghIuDa5lkgl8QB70UvXCqb+2nqVflzehqqkpTPViGjG2Ex6i5Obf9scNLmM1NyJkgwxyTY
ThGJ/QSjEVFusisLtVOw3E8/AW7z4rJ3uW4nF9k8SZgki3rtagPlWrhWLO4DYi4e6lSA8gANFNfs
rRV6WQzlfMubldMH09nWjHxLXto5sIhZ6PIwdJGtOkXEqhpTOR19YhQH9oINdkpf9xLH0liv8xmU
pOfw3//ckp9moBXZQrnQNnOxQ9Ud1MMELFS8GF6hGRIoWjWfCj/dY5Uq1DnDXlAlTyunIT+T2h/T
yCJR3AqD3dg5vELEcXtl0arLCbhSCRJXCgjhMfCuTZd4P/pfI0WDmgQx32uIF0WIfVx5fud6jcrB
VF6hnnBZAWEnjHe5zAa+7cjZFTK13uZOD206JR7V/dx0/5EmUVHbaavmy77w97pmqG6S3em2vHwv
+//ySptjsHBLxgG8vqbdsJiYPHR6BiMyQyBvIj2eKAJ2xQnDRF4=
`protect end_protected
