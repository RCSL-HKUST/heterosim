`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
C6a+vGSrwnlC2F0A6D6DKUC9HO8QFe+t+8ngRVvsSoOvQ44WlPYSDCf7I8Ov/RQyDlq1nPps1sro3w+PGu8IKg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nt1mRgyIVqP7bPIU/XnfBJ3HFPAhcjm5dVxoKiCkwykfMNWN8dGSbcLOdWuwgAayLbD+a+DQh6Zfn/K4qOUupHogbRwmtivD7aacMo0wXMoRLIoHS1YPRkY/jBnSeoECLRkZUSeMwyfFEcGZ3emf8krDZuWu6XrXBa9v+xpwcPo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sn4vEI1apuz4LjanhkzMT4LirKE8pRcLujitJ0pi32IHFtNtSPxJMUfQgZgf2sxfw7lo+CTsP112XiGD67kUBCp+8hXnUrrNZu5K2GsRy2ugisAHdrPp9FufbHPnZ3xTCavKZfdOIR06GoF5Wk8WBYOhZEmEt+/Uczqj72DFqPzdlAxCFPuCTQgeCzQOUqsDWEzBVOdL3b0mou+//lFjrK6GfH86EtC7ciQI27X5t6T4Pu8R56mgxI/GlTSv4X5FFxWwTX+b8Tb+Thth1FGAhlGpxY9OXs+3h84Jy3mmApAVBmVpIdfu3bOtr+dIUU/MnvFIxCODuDXgB1qoYNZo3g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fVvlmkAKxaA4pKdkgVemLnwP8JbVGrr7qy3DuRTrlwgkRESsSxYoUH1+jjE5fZmEq/WNl6ZYl8FZyzScO5K3UgJ+HgybVY3JVr8mkkfkeZbAgrpcc4SM8OEQrIsUm19aPLzC0uJvVlnZ9/bTAOJU/fMz4aA5IC2J93z/GqtxXiQ=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oUwnXIrDlVirozFZU0PevVHdTfbFm6I87nLHHdi/6BEtXXp/x2cFlpyGP3TS2DjWoQ5qksGlvVugeX3IUy0LgVmk6+JKrc9w4Z20Ogcv16DAM1my+XCiwZKu3Hs1v0JF3Xncco9vUTTSuwW2ngqEd3558I3g8v5hxO8egcugOkcPVDij28Imu+9ZFoNZEzzsZLKHBcCappbTgXO6uVPQJUrGR5yNRNijs6R8AjnInLhlGX5uegC+irjdI5mB6jrnjUD1h8ioC06EKx3Tt2EFs3WHfa7lCBPy/KY/UOcjhTulO3VHS5xF5Cz5F1t/vTZiQPji2ZrS7DWcq8Xtsbvcvw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6994)
`protect data_block
ypBtE/AtzwDIgbEpA6VdtgofexQgv7TaoTLfXOBGrPU8sLDk4ZcxfLAPY+GxWIn1ZquyZs5wpZQ0
2xZlBPdg24lhbsPKYTs+XPCJUoIdwJDH8iEeq26kRGepd6Tz6WdEgd8zyO28SZ38SbBeaCdNNfLL
F49wLB+omahC6jL/siJZKCN8ncskSrA3HP7PZukqUndtU1fmMdYGNPNeG5tK7BPgwegxN0AmDk4g
0r1IqNTlwcr0/7FyRFxVyV8gxs3+Dlo7klxStNckvHtMenWJ91iuXyjaDUaXAZlmziqXp+4Zc2gW
4jH2vN++ia6bgkHfLeSibJintpXtwgmF87DSntaDEyStrGQr1U/goQzP3rRM60iKIySvOR3GF182
bIH+cCPsf+Ii3JKNsJuYNilX0GKvjhlsGhUKEgDtMAo8DiH+cp58q8wfqy8qtYbpBuCw/drYm6P7
22VGcKlPj0chMMY4qMBHbl/MhGNhROuNJsiBCygUNQm38KrraTgoFkTxv/DsG3qk9y8Npf7/u5KH
8wdGvxi04gkOTCtxG4Cd97sFs78U6z5mk7v5+SLuOMvbnLE1/JU8BLEGD6KEZcaq3qw5MrB2aM59
7pkEh9LhBR763PPKqtxENuLuTdGAcUQJFvksQJdlBxnZiy9gF/kvP2/P8v3tK18pvFNz4n35hqoW
5x42qLcI1x+9uczJlGIawO4accAjt+lGvHt/G0XivdiAsEOemoHH75Mflm7SEHGPNjvWgDRL/2KG
HRim46kkzKtWIUVAjsPJKFFMPYsBvQKeBi429Ft7TSJ9ZTBhK7Ov0JlQiV72GQjwYOrEStdVLXi3
vv2R+ZocCWc0kofMpcgZ8yCi+ikojaYZD4ZRXmtq7QV82nUHCKD85G/DgOREvlAHWGGeVBRaa0q3
FJNC3odPsVP/r/SHuD6ZxxqdvVR7mlyU1ofhbduRNnNsf/4mlLkDwj53JBKnFZEIBVV36bYRRXdO
98MgTaHt9OoXp9GAoQnBimKoyGJwThG36meCT9eM1AAL/8yS2pz3GzRz9lndi5w8NXIzqkO1zLiZ
wVFfqOiIMAW54QtmxnP471Icgd59Q7jEomrxnT4ji9abnpUa0A9wkuLueHsdRl7LwOgG32L53op0
zVg9BI1a9a7P732bkXTY17160YlZbdqZLbBnPE6LxRFE1vAmzafIC0D/OmR1GkJZoVMXDhRbw9xJ
DY8SxfDJ0RMAAAulcdCT/YxE8UVeyWtRUh6ut9wWkszbpfzQxDXhC8DSZkkO6f/ZgJsIA0aZHaEj
mHuf02+U+6M+RLoNmLvdEy29qpp6ahkjcFJ8v3g7wIoKIM9i/NIiI+ZUpb/CGAb0ctGx2ARmdGhA
1FgMgNEzYdShQEZram4AqghgiSlxxTjOb+B58n1ktZ9WZBdS6hHQJpDnsi0M0z0pxKjEikJAqDtV
NomQkF7Nc2Quf3eoay8XI56qZe1SY7yEll+oPPKBCX8+MKU2W2336tG4yU4L9xcBzXdXaF8SOsiJ
xDPW883qq9HadJnsEiafAy29VjwCIJcerEyIgIwLNS8QdSQ30rneO1Mer3xQmu3CZkrQlZcu+Fdw
JQ94Ei89a6VpCXOx9b+mka+fag9lmzvZnxTNr1HEWCburFRN+bHsEFWpbH8oE9CYp3kV20/nKLj8
bTHVR13aXU6SKT1yNrxoplGGfRVpu+VbOOl7avw7CQBp61IpywQ27ACMW5fzmRM/Eb9X2qwZX3Tw
+mhBgr06fmSQMPkLpZoKyGcUUxn7zGkKxrCL99JyNmLOih+yMy4AfupYl3jL9pRXhg4lshhMxuEN
Cpq/wGKmuD9bCru2mx4SarD2KXz/GB9dBw/Gv9rD2QtkzSlEU5cYWjRePWhPT5z34QNS3+SKAO2C
qr8nF04NnSRZ53JCT2pqawTo38QhlZ7pAfdHWAoh+RtF3Gd6DRqTKWSy235W35JxnajgtcYZUAAN
Lxy1sax1+z5cXUUuwQiz6Rl6K/e/Eo4jjAeu33S/41I7sZzAomY0BJaxjle+kf6ruzXSEj78IdFS
U7cIMUHZEl2YG6i90O3tBIdkWZBFQV3TWJumSlFl5IiSgq6q+XeHaYt1OKTOJDmxnaRL8ebZQIdq
YBMtqliY0XoylXT6zxRa53h7TTIT8HQO1SBBpieGivnDl213cq33Px1gx1quYbslO5OwS5ol5Y1T
HK04Q5pIY1Y0sHii86hd7pVIUzQUJsOPF5NtY32f5pZWGPzJjnKfV0KD8t3RdV+TEO6LHZmCjcvK
k0f0Og3X8Co4NNSzjGbY3/jlmwwjhRc2Ft8LHk4CTfMBXwVvfDsddkzOilTO0NPL2El93e/KW626
J7sdE0diBvNXqqK/oXurRv04OlXt60pO/RfaYe1K5Fhb4+1JdJmS8tl8E9odEPFd9Km3zVEBaU77
6CBwQBNRfR4EmcPEw6fpBzqLb9CBH2CgDpvPf1RoQMbQ7sj/DnXG9FmduHQnkNK4QtYL5DdfzmQC
dpIS0cWNPJoGmSroQhT3c1LVo7eWDEGnQVwD2fGTEKPRU8J50TRsARCEIqOnXbC5dZwyw2qhoM+4
rqVY9XxoPiHrBt4nLCROyXKQk5PaQPRzMXDZvw0QTvfh0sP5UBDmR1T9vKNjQmuhgLwxcoaV7V22
WbQwygCFXxH5r3fwVPumJUkLKLU3lFL7UoiLUBLZD9FnCT/zFbv8l3X1q+4ugCsu6NCRs3ykLj6F
qIutOUcRRvi/m0l72VVJ4zkgEplPWan5f9RBSWFAt+aw8ntvKW9mLkmeOlBu6FZ0j8pcFEaPllXD
RJZTr8rYRtU7vmI7l9/xC2Zc0Sl8hTamnJrxBtmdLC/mpeGyfSsxkutTT4npuqaG3Etm1UrzZyry
+lXWGkae4t8DAK09aC9gXZ2Eg5dk7fmP0Kyk38fa14h9meRHzzGqE42lJUYAKeKz+vUmn4WZPhNE
+XJ6ASd9n6gV3E0GDy/UkpL2rXT5rwHZrH1JoeR17GjuewLJlJpCF5/zwbrQOgW44LH49KPFVIeF
5Bl44f+C4lllPBitK3/+DpLdpXhTElVoqEYmeIRNxBw9IRaoX5f2ft3I86H9aVMf/PBpai8TUuV1
pcHqxNEgr8IEdwsxwf/MQBvrNxFGZH5pUPJ6AEWqZywQ8+O++gVXOhcr7hfA5Xvu9bInXTJwIMtx
ElmgJQKJqZT1A2GORJjdiv7BONz9dUXIX4rnAfRTQH0aqxe8diOcRyLgCvpq3CHE0tY0PGHXGrmc
5kmun85pIL1xtW3V60yZoV6xR9BxsPCzfdzCk4+PBFQyQnwO7JRVY1x21mUppf4yBXItArG6Z3CD
/FlpFOrbaYMaEfTrlZTOm3B68/4bleJYghFGxgkOJ6gHsb4rpX9CkBpzFgKgJ/VLuAbr1nTX5TnS
GB1nvhfdpWT1KDYx92oRnpzuufpK3x8ID4X87Y0dBUA4UF+tMTvpX+1WBU4GfL0PLtGcKCTh+uaJ
c0F/83idEwJjscw+a7uiSGZJ3sNP+CQAJryRl6sgtRIgR8h3/LYJjryY4pS3bfE9pcocwhEg5aYn
yGea2/tY5YJ+pmnqqN0Nmlm8SlohGJ/Mt7ON6bSebSOlEq0hF4Gy2Zh345buuAbvxzwXCnjG/DyM
qk63rYLnMwwSizBJBMuIi/7sMAwlGPB4ecNacNTpqU9DgeD6xYuHO8bB6duCxPyfqYnMHr7a0Rwm
oH3NkAk65JggucaKGwrM6EUT5qBRVYnHhpnxU/ih2LrZ5mnUIovzgry4kyBxTPJTBKWYUMSfHLbV
xr3J/7/ztKiVBFooCht6JNSye7s0g1T719tAzrUrCaTbjd9DKRG0bfuHr+8Qo8dyKd74p1X9hPzC
ocs0o65aFhD41U7nD5rje6Loeyu7d/KoS67zbuPmY6nPA3LzLkSWHtVjL+SPVo6X7KhrHfIUpsLa
wqIhZAv78E8B3epoO8+fO41PqwfqHJlkH951TAHBjPUg73//719EgK1U1M7ced2/KK+yJZjyl1bk
cp9YakBCi9MGNGpiJFuhgexo1SxI2UrP0SD0Z09MDah7aEgpsTP6hin5gVZjywV84wmqiC58KHXd
Lv9kkmfp2l2OOgTdhlFPt5MgoUbT5DeNfIeTyybzeN5Ywj7LIW/rTKGVWAR+L1WcsX+4Gf2cDNAt
T4vcHGf4sdF9CqF6Ro2/PlDV7KBaXmVpkbqQLeQWuLXmpsSP0Do1gt3E4gGUCyxbivpCswCPoCym
Y7cYhTxbg5kpZaPrQPAjTKMGB8G3Q969JFk1Vc8kSuCWHK/6wOR2KnYOh6Qp94JJMbyoh56CGRFN
SnlsWQb4ZQ6PrDII3jF9lhw+726uXeJscVXP6LX+cD5nXgOSWo/0mCJ8tSDcW82UHQYqWqNahOXY
4nuOW+Ug3XvPQx2xEc+ZVQFZ+j17c4O3a2duxW3rGeBGEiJA9PCr4gOnrpZeZDEzVUZi1kRq4m5R
a1m/+y5j0LHbjgH/ey3F6IHsn+PJbSSFYgk1HQXnwpRADC8KqhJt4WsTq3jYiE4numG1PM4ok6ua
x9UhDdARwOePBbkdaogaU7vyAcFHv519vng0hDvvJQtvYfVJ4g+4yTu2SnS+TbnPaVrMvOyKyfmZ
H5EYd7r9wxCiIIgMUpdg9WhIhrovjX/77ibZLQ95Rq4WsPF0DlHMGzc4RDt7uhhxilKYyVnuEaE9
0CRiTmhW+LU1R8wYLHax/12EL1KvnkMhjh6TQMMIT1C7VIpxnBAz6bsRwi0M35vGm3aRJzUloy6N
DL9bEHNrdlk24BlnvO1D6tiDPr7P6+NeKRy2Q31/gF1v4U+ejxT7p9NyZdjthzwdaGFvfADGJMNQ
uLRJR0WZrEo+jpEP2+SCEZB4aaaRXbfZKLN+uUPba8v5nOPV2RMsGorIg14durPjX0zcUqbC920F
KUyBmJIlMRzRZ8e+l9bqW1cSEj+zgZuJ4EaiRLJ+gbvhefbpEN6OU7PSz6t+6EFpjrEvvF1avtZ8
caRoigwIXfeUcfjS5ea31pC50uxqI84FXidoDRppahvGv0Y5HBmLgrDS3oMZfmONySLYYH/yJjpf
w7BB5EMSfYII7I3yf2QBDOEujUZCMllXqFsdRNXbirN8812nVKqUucqNLOOH3+CMljk7lVXdaUeS
5UvIpcSIWwboNcYzi0KY2TKDqgMJ7N8dChwF7ey6Yr3Ot16t9GzDYRkmbBUjMfpEoMgQjBtKQexE
DC18ifLbpVdDRWQc1eZW6r3n/upKzN0v3ySo6bYQk3t4xZqLNrvnuutHOsblmWYy6TbQc5Im+NPi
rY1pnCD8uQ2l9JPOdf9s0alajlWUbT2E7E9q9c3AuRHG18w+8iGlZL6jG+URphPo15gGoxKyTa0M
+8XNicGLA/SmQRdvrObwGRvnftOL0usrKlr3HsgZb0hWnlBo3Pdnvhsx5ww4Ec5bzTgfl85mN5Tw
8x6jx+zgkfT0zNQ7dyFHCIQt+jEt6Jk731cmWnUuO6UHJwQdlDgbCbghuivqlymMVJmt/cgwJcVi
GcBoDq2r3BoWxk4t7nTvuCDDSD2v0QPRe3ssQZjiy6d33DsP+MZ79IUUrilkkEIO1rY5rTF25BY9
7Ceg5dqr4EzCtT4YfZifmJWNXkm9W6rvx9+nBMkEoXFo0y+GDZBoHzmEwVG9VajWtDTzx2akP07I
IOrkq55Xb5RjNJTPzMIEP0LbQXzcYLDBRXsWCM+KREdNCluHqjEZfI0XlIufLu7iuRfgmDZVqMHA
vf4PfFh/23rUz+k9IwcFTYpY8l1SaIiXnRZW36HMGIZ0rvfihkL6PMkgXZezLxSeLE703z3KavDC
imZFAvT6xD5hyla5MnpDnov7AN15xUwWSlqc76L3ZFKOlQdciiDOcGF2wj36FsMxArfhzYST37jm
75rzN6zcdHSX3NBIzm3TVbUPP+3dwAfcbMWbj4gyfNCMTDBQLbwv7HxT8u5v/BmFkR+bphYlHjJv
nFziTMGQAcjyV0tAsz0qbhm8P1386coaT5o16QZ7TJ7e+XayXtIXZFrqoX2mXjaBlqK/a6eaxofT
7Knf3GkuePEFTNMimTrqDfrZqoPgEavUEdfmz+XqWemk65IYfPDrSN9Dqo5yjYJka61yxhsEFZh/
cvQfl2a8ZkHyRnlUVNNbt4KkQp9Sba18pd4E9lC4L/GD7Ld+bAJi4YL6FSn97XwPLDNLeg2Opui9
cq55m2HhIzDezv3BgWm2P4w4tZ3fUj6PWuPAmgPCf4z4uNUaIh7rFNfplTT4rbkkVnLeXr7fGz1F
/cz5cq2QyPRyaK3CuUJfj0oSZuAb/0cLSp5XtFUXpoCPfmabwgUHb8YTr21A01W50BjVRIc5MPUz
WsalngpUgYuRtdPjQVpTVKYNn+bqFrE24x5wG3BE1pIyl28FrWAzZSi73H9oR0x44HhPFtfNrcVN
2jHfb+PkLAJCJNtMZmeLQMKssu3tVsnfiHzLGujelikh0Gkwlepo6MhEvcCxzY0P2e2COA1CXTZl
TTciPIm2zp3BcfKYNDqpWa3fhJc/3susvawXiLx8f2MCfwxQrXnyOnNVxpUVqKJY9jg+CVrg5Ooy
rHbTsuLzB/DjOWkIOtF3J+G+CnzBlsKLL1V+QAt2VRqY+bHoX+eeEMsvirkpourT8ojeDDh4iL8M
nNZ9NEsAsqOOvR4kA6EPXz5gx2+P1vat8I52Wc0SPyMzWIj2iYu6NCulyYD4RqhzDA/2++Coke2S
tUYsNQ5f3KgFV/HVPxFVSsfanTWWZvvRnTrlcILdtLRiXYbXe1IVNI/yFouYIpwA5osmvac2wDI9
XaojdorcLASaB3JGhGqTGoMuZcIX5gscyAdQQus08dD4VlqtVSbTWSPkNhx2mOF/YPdxbv6hcH6Y
Tt9oJ8yInYHqd2w8661THdMQc/aK88fq39jg4PfB2ezAjMi8E/xwBiqPBWPmdYImypxPhyQZ+SoP
E0yO9BuLpAuD3HqPdU8kcHfH3FuohZsi95k4EN4D9Gm0Y0DxqdDvN7UdqaMBra86o9Onjxu7h5aU
NAhbjmqzFPm2cmjEReVOB2/WUk6dmSED6Dn3R1lT4z9W5ShydreLi6ZxDZZ3Hv2B6hCgZ0XZtsTz
wr7acUfZ8aqCzog8jtdqe7Tmf4NIiAHXqyFUkiSrg6GBuBoSS0f7WglasmZNQ+EKAcQjCLeybBIr
LOw5TaNlpxj8tTH/L+MPY7T2JtyuEaoaOy+7cN9yfPypnEF2I5/0Eeq1lyPMfV2fhnanw6kau+YG
AWqlsL9UlepErDgzbBjKtITVvAIi/D65gWXHDqGM0aQEQvksGHdZJ/ab+XzsA8/RFQ7PCRevJJ7w
brzNlTSBUuiccF7ThwQdvrfN0+/awWvlcUyUFaAxD/KVjb5Vetjsz9Jj724klRg4/LdE5JsMFZni
3fv0qglXjI/l3fE7V1CiYv0B79g0PNLjl/B7VJIw1qpjz8OaJvy8UoLxq0V1fe/R8DlGC2HZ5kfp
GqgzkMnbL/AD/NA5TuTALVzWtvZ8CV4hOwWx1JxOP2NY/HmAYMsRcBhvzu8+H5rRGoyl40u9VncB
7pSa33BAF/osFHTeJ0mgX/ns+5qP0kyevTsrRTY8MRTnU7qBPpiPGQyxPTovnzCvK5gmtyHUw2NE
2ZztBJ1bV9IPnB7oMM1D0SoWvhQ9j7XzB3EQX770r8EhwnuFulAIJeOjM+OF3apPS0d/HnJ7KEKV
nxps5xcP7LZUEHWHMmcZ7Wo1/bA+7EKluFC3zziHiBQ89joxXKH8Q2HxrpXxNSQeB2yPMiSA31YM
5eD6gXkmAWPvIsSesA3RlSxyFPfhNXweP78SbiNCgupyxJplvDnryPpdU87a1oLZOPLceQuIiY2k
M48qigYFDaVA9R9r9UTKp9cWGtSgKMZMA8BAHJ+/p6GbJg07RtEyXkTwjQJqkWQByXdoRqTttdw0
qf0tdZyvrKYgUUdgYTIXM07eIgNCVO8ILsTXimn6iiyn5TlPeClVi3RThab4zBa+jscTl8gdgOMK
kF8ytTyGBrWK7QdX9HaeI6c9aksn62e0uDtZ8vcR6abc/pYxng/q1dcwK9CBWk/AIAqTU6f5L4fI
w8ya6OMt6XxDF5YZh+ktbMpYcs9bDnm9Kj0LgLDXsiXcHC2UEVs9QTECSL2COg6G5EWEZm8EKGSM
qKZ99vBV43QEq56yw4gO5RCBmSkIhVO/eVVnJ/g4AS6FsslJc/62/YoOa4ZKxqFUYMI/L5vKZXXX
ewjWHwPQQxEpr6zqLSJh7MvgKd054+MDwf1x7ig8kJgA0mcEuDMZTR2MfikSXteQAvK2tP2TiQBW
EPaZYOcFp3zfb6ylESxW2jBftElCzSXLQRwuV8GNWQWmo3NugR6TSlveo/Q6Q+T7J+5jjObzOE82
vnqxqdMYgQWKCq/CfDzTqspZ2W0yxOG+IdFdmkHEYPstuf+fTsK13FBevw5QtFvXBw4zX9d6f/tB
wGrfarZ142QM+382VQIPX+ZO/667Por+jIxJEBHuVxPIrfTpQf1+XZl5KAh+WcO7LeTHdyIJYWPV
6wg2JQzdR9V/qwmLwTYhBecUkJ2hEa0rcJp/7fc5wBvKRhJVgwm2qQmk5/X5aYBXsZl3YvVvIGRb
7+K4ydF6cJlPKW/ZLoK2r0+O7qBCjr5Uu8nIEIQQlE5cFg5BtVHHgvmxHOKqMlKTopc/6reK6o6C
l+6aeyRiIH7xAN+wBCK8w4N4HtPYy7Tgkg3yGJaaIWjJTZ4IIzLz5sk4OT1I1s5eKa/a65uEpp2m
nQw1OHFZHUnskl/ZU+JH4dFtXs75TZbYnkPFId10up4YAs7xCYrCr6Fz+Oh9FZNo/EbLaDQ5EPC7
Nuwm6laTvb9/VFfsv+0qC2fJtHPqb6bOYDrCjt2BA7J+9xEbLH6YKIjsHa4+e1fNm4A889WGEvKA
4C6cAC58Ua+nULWIMT4JB8Gr1Dvu7CRAOx6Ey/5Cl9rzbvr3QNqULfCQZu645fKdMAJYz0FH5exi
h0uXXqX8ApJX3H/gQoSZVxjdGiwm3PvkI7Y6RJ8GWdCgEhZJHJqEEJeqs+BhL7Dj9QBaOtXuJBXG
SLP2CbPTDHNY6jchetBi69unbAjm8GvUpSP1iPFI+P9SiYt5AGQ8CaLUWksxLnKI863OhKerm/Gy
4DmSPXtmFhcSa34X697bAN2aDsJlNPCwh0u3h/v3pCnwZ785hBSYafkL+glp+gMrAGm863EPNucL
M+NNZxk3TDYhN1X6Na7tPfINdj18Y/nCQOlvMS4EkByaa220Gm/D0cvaV1tX90IHXKEruSh5WJBY
LcO0QM03c1+U2Hmwag==
`protect end_protected
