module our;
initial begin ("Hellow World");; end
endmodule
