`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PN1PYpNwuGpIyQaQXLk3VFwOMWW7ZaudbN4ykmPM3z0/FqDWc145HwNY7tVhunR+pz9EztXsKJgAloaEUFJFHg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
naaDCYTNlArMUsKQDkFaovX6iKuu+l02qA2W+dDPAme42JtmhdOr6/6zcdcoRzjgAPSruOIoecFxaN7R+CzSUE5WPnqqSicqJRojOF8m79oqAroiqFPZd3kTWGYlidnEwINbjLXiWztoesK3YEVjkYGUt6kbJKfmE16AH2/YHHQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e/DqmWNFG7OgqhdECQSJIxH8fSQTJ93K1vKRg5FPMmScMHCMi00oVALXTHr1LWTint6hXUdTykavcu82LntWfFrGPfV1m9OGaRj/vsBC7a2t7wifc5CbX7yIhsPIx8lnsgsqnS8XN7emvcmAxZjDO09HgXku3UZKyOs9I/YzG3YQwVCQ8rYa7kAbiFcHcT2FU6IrnfTbrkvwdk1X+KwcVt4+4u7hQjkGLtPw5D09LGoO7wYVoKZ30rXP83kUmE0TiDn+pvZx1M41mQUuMAujwuGAEbbky71ctgW9hFrtl3gsOCioShg5CAkZMp85qOOs5Kdtt3XMOPsg0p6pl+ZO2A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cEZPXBHpTbXLhc2WOo9AFP2Xfwfk+LvJpZm62D4T9OnRp+OSmE+hFWXdIRfKML+8Wb92YJmiik/DJlX3fY1VNbK4kxGxCBNm+isEPq2T8yzEIXa0RPbWsAyJ3ybFpYd4XchjVL03Skw0lGs9VrE8qh/h05i82064O9MxSbZlOLk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MN7B2cS98H5eNYWFCOAHPuAFZ6SwQY2+uq0NlECNmWbNMs5owUhQegr/Pkj75OThP0WBMPzWtdjwYOr2u9UrDQzUI8P3RBovUbptXEi5JEANQMuNHl/1FDqOKihqJ8R1B6oY1E7LGw872HRJrc/IFWIi2FE3z4qwCcpEaPvJ1/0Vjh7AKxalj8j6R8Ks4EiGINsIXeiieeV+/chuxqZ+DuUZxnd8k5nEgIjmI9yCKujld3mJCiiG6KUcYWs4462oSIoIE1RGnCzNR2HprNgkzRhg3SrZvRcskefAUghYeLNwrQtVd9HxRoAiw3w9ZfRVuOxmoClnFSZbb0NUi2v5ww==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14091)
`protect data_block
tSUIpDbJnYI8tmH5R6xjmm/dAxCkDhlU+lg5DIfmgph+MEk3PUUkDxEI8uAwwfXHwD5P5+5ICLkQ
qTSzjzyRSvXuMwA7R9wduGwUFCRAJnn5kNO8JNwG2MUNbv8GvcGGUoEtjGpug7SEfzoNP8PVk3vP
tDluR05DS+i5JEVDGhcXqaaS2bUi7O9YHmYGKaniMDbaVeI7DsOnUDl3oS8b0odSL9Ldk36yTVW3
QpAmLxyD7pwRGOh+YodOP2j8QQWMUzUoMnwuIy15IZlg/VQAd4JCFWGZ3Z0Qw+docL8RD2keKIrm
f6Q/ur9jB4gDvwVxT4nILEicYFw300dCLiD6lTrI+ca8Cv+W5pDhzY+hqIuNaQ4zvd1xsdaTWhm/
nu5EdOt2Ui7za3ZuybKdBuDnCeOW1R+Ahgmgu7TG1bo5CZn5wbtIU52YoYHIKwN683ZkMdrboTfY
eGmBgcpmisTCMR/Gj5R53mjIfcTEb5PKhFbnzEuG/PJ2a8WPAop8em6heQPdGDa7mSQ7OFeJMC9n
2FWtwQEpI1GwQt8g7j3gH8PTZWivZjHoS7yfVmWyFpKImIqzz54WwkTfCDPf8zRWTY7w7U7sOP7E
ZN42rur31A13gHsLoq1DKwrYTXgDKIYRuAjN2oDqgh1qhf0wuwWi0WCsHVzSUP3H8pbBTA2yHpm/
uZvJUtY9X/VxyZtSmzemuioM5lwSQ0ebCc0u1AAoKdGSPRREug1ECcg5KFqlhbt1RuSEulx2aJdQ
CLRFZmJruvBxm0yK5G08Le/ZU2HoZhXEJNZNMoNXjQbqz4u3/LwUupvb9W3eVVeosUCc7EJqKOyF
uAs3hxCbN5CHXsm9TG3FIdrtMCLBlBvrDLYK2/ehWQcWpIDHceE+qtd1J1Bk2ANWLdOGaAv3tgIs
TbBF7wcVjwfsIrEvwBQb4MgK4NBsgDD3Cx+w1iaBmBr84cSD0e3pHWW0nJ2cSKlM8TyM7NFLK97/
XmJfcrRsR+DtQfwWqqmNhjhyBT65BK/W5d5BwiiQZOYnsIQheaPbdqEjvpadVZiWgsDNdwS+r09V
nl9Icil5NrFQ/2BBE0/NSHrTYKsRsumzND0cvnZA9s3frXMhG44uM85dTDPPaNmwdXl3ywkufCUV
W53P5kAyzizbzMqs2l9Gf05ij9PedBOs7ojpoH9VJb3+7o+HXuMsH30AWYMLLwxy44IiaWsmPVNb
6wzHl6rb2oRMiG5c8NSkt29YVtE5jfATXI9UWqDexkr5/g8AL2sqlgCM/bhvTiNMUPsMB/QREPuG
mpcnxI6psuFVp281kmH6xfEKnuXLhMFLLBUiTLNlPLaa06l/6RTH4srgyjNLkcuEOPRtKHCp3ILc
OpovkBTa++73QmXt1V9KztlYnSsM4ulrY0yr0TeGFOvMuQT7dFDEFhW+lXX6gL8byrvtnrb3C4w1
Zu1WJ7OlsTusYoKEBN8oOm8iPpv8NjTzeLazDizWNfgiStYeJTg/u9oqWx0A8np7yOqNOwII/+qW
gdP1XOS20pO19tgCOCmPjHL8PSwqcGW3b/2tFOmHKq4Dwjifl3AcrVWAXQHj+pCnSJigtcEsIiez
kVGoFrXvk4Qe1mePqla2cAqA2dvjRlyHT6N2jiRTK3ZQiriacLScgl+HR3/Mx2SJcQYth0QXvct8
U1MlujOFZPcctPYPgmEMjysY6wpOnFCJokuq0WPIWUfitfqVuWsdzAR7DgLOB9eyqCKhP1CCvPdh
tGqVy2DSWUBnzLir5pTzVK1q0OLnU7hV32joQCtpBz+lnCB0iIxjmVnYWW40eOrwr6qarWLtECKX
4kY5eWPCIRk7n3v8M5x+iiDPNeTBaKXy3TpNcCoGFPEQIffHyoC9X+wy9f89xl7t8oc/g8e69kGZ
5jOAa0+Lx8/9oJoG5ppioOWSooS0/XyZGtqP8zIKc7v4cohlOo8ByZ6nny3cqfz0bh5NUjzNEPcR
dMT3Gq9qHBjTqCAmYcWx1wuPAGMi+oDzKjRI5w/ZOXkzw5p23hLv9+LjxM6flg9w+H5+sIKmNw7f
f0SdtsrN+/Sf8KVtB3fqQBK35aWIwNEyGrmGeT2w5eeECyNq1f6GTlK+lwTz9LRXq6oZ7JrZF9Lx
KvVtp4N+RKPVH1J9/MQxJZpbPCmoSHL7zH43XTdB79gWjLaPG9kcnQQsClDHPr8z65Tc9kEcWe4s
tHf/LUFrpl5K3VpX/ZilV6P2Uk+G4ISIOtgxuGcXQF7FobbuNiWicFfiL7WkZVoBHTKb/Qp0z3yz
DS/ALCMHb/7pSy+zW4wCw6UP66O7VILUJrLx9qVsKrjGR6NpuyADL8BUcFYCpPux6NCU25lneeNp
BMRffMgq/K7TnpnaA4+jwZNrHIxNXjftCgpSSqSA3BpqyR9YKIJQ3kBNPkZnENKhv44Ar41pscYK
UqvOgzoa8H8Uk8VviZVfINf23CvXfDpZ07NxdgAq4QP1vc80WlbzmFjJkHI4A/6m2+jfNRJFQHGo
WH4LMP+O1U5/n2zFtCvWvAZYKRQZMggdV0kKzdJS4IKFGAUMQ9SwwJNusoyFWfeObWBIjtZSXLVa
fb8UB59x9JY/0Zl2yhbRU1xm4+mh42uZlBqjNnSpYQsvQlkPhkcagXt27xLPadWZfljgZikmhfRV
3oUvuRkAOAa3lgw2LVhGJyg+tvMAEZCaZaaKk+74QwWOhLLkyGAlhV+bi+VZs/XVuu2Ecs1wrIFl
CZ2QlRkMx3cSwxJJ9HaJ7sAHYRhrdhXzsCs6xw1WOFAvn8JO/Dc1GbFhDKuw+Poc70rMtQHyfc1u
GwQ0+Usz0X4wriOHwV8Se50KMcTxm8MQX0pxaEOCk+lPeMY0TPybZRZlq9TXAgi+ElIhJWgbeD0/
XBUQTo4lvQRpelRTNl4aBDf6ARyNUDct2R6k7GxQUZj03aa3Cu9reeM6/HzVpIlDnobaiGmEa6E/
oNl5cYhYnZmKtJqbQiviAnRxvW4Occ4mGRvZlZlSSYJnvR9mvoAtaa3veMqXpnZ3+9z0gIeZvL5W
nVfU3e/mXmrx6RpO7wotkrDXDhh1grHJ9URHpLIsK6L7lvyz6SnjCKIisKxwF1YBqzdHEPC3Ulbm
nsSt1g/fZEMd1YFU7RILUjf0cI2mP47fVNKHfPjpWnOkFA+ODjOGhx8kMZCGQi3aKFhw2YAf5Y4x
B3aUEOYGjp/KHVjzXy3atJBc8LWXhgZWDeOBLzgl8YkEZth7GWEkF6aICMJfFoipw+2Ad/fNF6jT
UESqMDocDu7tYHOFjqPZz/jJwCWhIbw2upyq8Hk9POv7mDTfbCVDgxs13J6q4TNjnXR46+5zJ5wL
IpPqin3w94oNWFFKnKBBpmf+WvirG+Yq26VqwBOoF9Bo6JurAD+6Afo5I2rmkYuWUNCA9brsEVBE
BlUmdW194LU1hf0V8nK7yo+2S/acEyCkKzjaYe/Tt09dSR3Zn2QxD3wLFiDFOqfYv13YrD/yddBQ
j0mlQQH1/7+Yd5XYVoaXqFk/XWCXfSc+WD34FfHYo0eYc51bjGABjU91rBzf4yiX8gXDi6McBovY
jKfj0W9WtkvDh4VddEbveJER27C0b+tKg2e4xSk674cCjnCIRDY2vICuXDEIB0lT6OoFAl7pRzr3
BuoMZ20ZvFofcdjryWyws0ingwadOqtF7L9648FK5NMaLdi5TNhlwFNFvK3WOI7bN6/lluBA1wsB
fIKK/Tc3sKQnGt2uB51BJ48Y4TCisZ8+vYVsvlMY5/ydRYBhECtl0XmbYR5pieZvVKuSmHz3KlHX
AXfq1mHW37izN6XVeVxyHd3O/eMjVEntB7Mc4y5DQRHOeRqrnEex3ev86OrddmPEJn7/iplrnqFJ
xf29eFc8Pmqq/maIYlw7K4lilbDuGdCE7BjiaLYai9X8rM9ak/NCQJAzrP8Vnhhcy5wI/EJWtz0S
V8xxklGrb/12Gmbvh1JRf+ZzYmxqU0esSknvoUMOL0Yn79nal7WPUQbfQ10/X9g4SoQNCBWVIgcu
cCUZS8W9FZG3zxPiHflmm6JL0nM+/cvFyhnHYlWsLM4GfHXeJghyj36nnSxzoT+wmpdG5Mo+kvfl
ffFK4p0t1DBSWGlYOuf6H1e//vJk8Oqyno3EWkTgIm+7akC0LqBWnXQanooJgKJlWOzGAhisbNqk
XrjKj9HAWcxXZo86MR83IRHGrToUWT+swIPVS14u//17Chk1DYRILqGyO/dTEMPQLHBc55bFFJYG
sQpQKK9LNIQxJxgl814fgQjh3aUQlXMnxW2JzMJYIxtomvoOWTV2onZb6Ktul/rDt8ks4bAuC1g2
oplKG6bOXrdIW5cVUaQwhQqJ/lvYaUU5MZ6PBaPHV10wYl/SqnTsgj5XrmoIJFGr+ksvIVbmWht6
UbWMPHKc8i85UuF8EN5pdMjD4UZV98SpaVshV/dzQAln/VPY5RSVVwVEfYNe3UcI/hbR867jIItm
Jsmd95KLvHEEZ3yn19d14x5hbqDRvHtJqGv0RnZoS4PBt0iOxuVVyrS6+x10/0BAQR5kQbkT0/ZP
s9eJDR7gj8oRY2CYe2c4dxcKOAnIMUIkbM9tZ5VToAKa6UNGYty844hzT3pHSwEeZ17roYaoBXoN
s3M25PvWRF0xnVP7XzCKKYwIk2zwO+VoulpIyCZbBGfaQpDB81ARAuT1rf9/vDj5zsVF9A4/X36c
IDQCVRDvhoz6HlbZawWfSEtXcX2mdpP5SW9uNeY/AeoHXC0+yq1Degxzq/YeQF7dn3bVA4qNvtT5
vbLqh3g4LUqDhkIJNtrpiCLX4yvgJbvY2hyyyXXJ0DtVKTQ61v1k+BgsD9AuK58/sIV8UCdUdwIT
l80+g4QIdIYJ8K27xfLSyMAjStlvsyKFFEX5XFgKE0uEVKBdkIrY78EQnUrLxg/yzVkEzU4TOiBx
u10/CXGUc2EzrnORR9lZuVAvTRcVeWY6ra+kJgCPxKB7EfhwCQqmH3L4zZqOrxYqolvgCzyVKhKZ
Lcg/WuEq5Qxv795WT58eZYfHx2U1OvBWtE9oYYaooDJ47rc/WGzn0ipjHbcvO6W8fVtBceQPOGjC
5JmoBd83gJSybSl0TYLRdK5KbZJ02gayiW4rvgL8M39r6ZoB1OgNGi6AZYQ0hAc8EUHfaVxZHQCu
sUUqi4um3xW4WH7tg9R0r1p7r1azK/9dYFNrEodsbNh30aq+5ew+iWWdgPJx0TFVXc0ErRJ72RF4
cQGyLjKTlIzYqgidc+g8RH8Fx7HlrFje4XvxCcUD/gO9fgiruxsg1Ij8OD24/2cKQMxU1/91fPta
9OmgCR5NJMVk2/z/lcIM69ioB5dAzoSZ13MkcpbjH/n6CVBxDwFcmdXTahFtPmrH3Lj3OGQP+I1e
gxUoqHI8gJk2qYs2CTFW7MJihy4G1qUmnklLN5LhXZxBwE+jYY8m/4U8+4qa1pHGM+9RpdEeHo8Y
+YUDh2eyf4E762NY/XFhCE+VmDeuE1m2Cuz4KJNPn/BEnAF7evgtV1siQXH8xS1RM51hOUXO3AFH
QH5I0qihjE4WpDIolgUFCrrVx6mUNsPBz8SLtnam0xA6AQPvnqyjTfY290+888002KSXpi84KUvs
QriCAf54YzuOLdm6dzAjg+VAjzVWDwgQFckKFV9IbgDOm+kxYbwEqSt+xMo7KikdpF0Vjs2o+aiB
QxQx0i3k2V8Ttv7a0NyT9qDC5gaZz00tkCXJf5JR8bt6hs0fQi9plPBGgVngv1WCprN3JT+YVPRY
kVW94l2ehv0VQoyx4gAOainAqL6cZQHLHnh/MQG1oqx4EfAwKqa8HpBCdXnv2KlQ8ZfDmECkIMyg
5iQ6ultDaDt1xyI0VXKei84ImuFoBCrOeU67+NDH+TYs3aJuwNQ6fQ2xS7tQRiW6BCh5ZXdXRmsJ
dppGqO6rYffaHRtqJzwuaOeFvO1DdNG7bKwnR/NgTLczphDqLwIDmWY5SpKzymHvuioYx1OCQzg+
P8ibuasXF0AkE6TYn8FfVmuI4k5zIpyXldPNz7K4nKhW4BlSS4yVY+gj5Ev1H/fhbcXVpvC6Hu1O
J6V6ZxtgYBnH/bwQK08cfQAyVe64yBHgpJVOq4R7Bk62y1ip7CnbnP90y2uTWdWB7GAq+pFZyHrB
ZPfHXfuxZL64UxZ8cdiqsGu/aVspA/3lcKjdo2uNr5g83rhg+rFAaD8OLBer9eNNd1p+fVq3admK
xrkDcwqMvDVfE2bh32LUuPXuaI7uqlCCg1PzZzVwZIz2hzIpfQ7DbJ8cFrtuxBpDczqbNMp5JdYV
rgN5+rmSYv1qf8eMQnS0mH9ATrNGEyC8XTILvzQZMES6ZZgGW/aFyAWhYd2gSEVg9mqcsEly35PQ
0fBvPbMVYoAdNsdsxhtKwZ6pvT6QksoJvpJvTGBiPpOA1+EQdHM8zLRtTJedZP0CS7UdfUpR82DJ
xkv5FKogD2gKbOYM56h+tx79V+vTNa+eSSE52C9A6S6je5S4qAwUOna5XeZ4r/7PG5rKqFwb40+s
ECMX0Wjg7cj3GEqegmKsJqMRL9thZXAQDXNtXWnNnUbW8tD4ReiaN3NK11EAKmGXnYqCwbA3+Wwm
5YY4VK8UJciy3IeQYcJck55SzX5JlbWoaBymteh8e8/gIrRuAjvdyM3HvDbdVmLNuB9l5qwoYp7j
nW6OCT/t3ASAHXJ8zChCE0H5yWEa3bJzfvGlJegjt1asz2awQ/Gi7MIZ//gkgWGE65UtTSDOSFsb
uS+25gGyTkg72p2G+lAC2UpG83O8KEM+dTRFIX5mHl1+w+He02pX4kVTWLfJ3uBg3P9FUUCQI3CK
hgwFm3PEF422AyB3XZLnBIyJoUqb2ktEvMMP3DFgVv6jBTgSXKpBQhN20RdKpb26CIDRob9mWcaQ
INWOAaFx9AflgNiqqYp2e4NI0bQVxpbqLYhBzru+1WFv9go8quI2t04Cr16sNTzbBmCCnsalS5Qy
IZ0J5Eq1uV9b4IzvbzE9e+6gHTWW2AOXEKVNOKtCBswiVF++ymr8Afs1f/4rWv8r8Z7IB3+14ZII
aFl9cSJXh7NlGUc9Efdqz4smnhrGo+BGDbTQ580bL7dCIxH4w88V3UC567cAuls5FQNsBEq1h2wB
fq9K1Qvxxp+l3sd/Fdgk1B/3rnyLpXRaadhm1EV6yktgvXlJCGtlTnnT+svZn524Qxjx/UGY9wz5
N/cs7wflWmEaSacQhlQFuD3zgLhWEyb+cQh9O4y6WdywdGMz4hgDUbVkuvUHXp6vgw3RJcYGN0Jz
FSPZ3yMPrBZNJxdROezIyi9xpkmhMy2R1h45XIOYkCJ8CkesDqs2QBSOkVMJCAeBg9lQQlSuUm8g
BJuquK6q7nQ9W4W46/2lJ1XPG7v5yAIGC15C7uHcEXXCs7BpOWHyRM/PsUiug0P/3g6S59LCgCiA
50dnNWU1QIwImQVDp2NR4pm4cUzSJiQrzATlAtzZKhqwNGQGOa6bttAELeW9rLDyfAiXcp0+ZdSv
h7gXH90eUDZM+ZKQ1oLzNs0ewHjICb/lkIB0qmz/nIINEGKun0bp7DV/qDxDNado1DzALdZaT0/9
VE+d9Dalh2bTgootjJA0PuC9knZx5qQWkB+TWebBt1LyTY923KlpjyVzY5BS7L71qps1kYH/6VH9
0cJzJqnrWpN8QBGJGoQCF3iHJ64boDfM7QGa2CepnpMy6+MtqDRJ5GGEjbLhT5XtSKvAWkzyUHlH
JV2zaFzSzHrJC8PDg6ul8AMSAeTwYVpsHxraZMvQffJeGNl592tKA3ULJM5DOLv1NP1EwGi2BtPt
6g/aDBjhRKt7Lr5ztRpYcg+ZVUtgtXlnwgJk31PaFau+sNZfo37/N/8B0NY9KXt+Z4nJQgsX7Gkt
R5T0FdF/PFylE0II9ruT1xZp/yQENWKRO4TcXc4a1930mvrQ0HU1tb470UAKH3agCuk+dCVKoiPY
NatBwl7N0FZrB1QWaIl2feq+f+78dJIWSb+r/fVOpTgLicn7eXv40ez7u6MfpudabVMhbGD4WLF4
q3qbiAtKHh8rvXyr4/I7JOXvtHWb3yBMrl2+jBfM9dXYwegJsIWN09BKDPXLZatao3VCG98tiwKP
joeGgeC/HF6FHdOPuj4RXMmmclrGx4LcX5XYfR6snEnDLCDPwDUnlkQH8CKCAtbeXsjWqITSd0en
kfs5vpKyIubQoQUgIKIsRc4f+NcVpnONp/Tt1ThKvoAhFOBCfdhnweTXvnPq7+dNXdfusGscBx8r
vUEhZ4HzLNdMV29vfjF/AzhrIJA7/uU7DnlMZUyvo5FlENLVRlO/AuWj8Vt2nmbjzj2jCbGXPv12
ke/0abUQ+/ndQu4+EP1Ww/n/sI1eezGcJWDsi1Y5y2UswuGVKT7zpuGCvLgPOfKxVZ1CA3kZoekv
zRrkoDZftZkvHUnksGQubfM/blfFhnPV+gxbHLQoEUqQ/qwGmP3gCi9yAM2aXMwz3rveclW/yhS2
WjkD8jNhrxwwqw2cDuzYgn7bynBHegHGZVpmrhX/f9NXBHbfPJjWGlKoInwvg7GxRMYgfmTpovCM
Tleu1YEAj5Psk2W9G9d50SAQnQWlZxYgd4E0bPSSXnazW/LO75uM4nC0Sv7meTE9lmuuebXhM5Fg
IMoC/Siqhzmt5qOI4JvPTn4UDc1jSSYc5MSWYds87dUcwCCs+MPaz3JfBpJuwY9bGPO2lBWfN/Ux
p9s/i03qkl8zM6cMef8XLM7EQX/mkdRCW1BQVB9qaHrb1h8madYQAFNaX7sxugWTa+5/SlNn1HiF
c/nMODOKnncJYggvuZzi9nXDmGKiwiq2dhTptnV7hsw2znbWhxAdCGASsVp9GzbaKp5uNPUbC3M9
h0DH1kPuNhtwjxnj+2ExUEcdY4ZNHWA7u14ykzT425w7ufhxNNDnMhYfunbfzEc/V8mNNoKGKb/h
fqRb6B0HOv2Tk3Jgx7NfyAgRXEf4SFd2mlRxTXv7XHbH1iir2vCpWzFRoyRANKrntXcncRvfLX4o
BFGdnP2VO2PTvyBhS4YA5YVvs22R+uF0201+9haHDwsD6oIG4hmsg6XqdvJvHqOBV7EbLTbq67k/
p7iKygAVc6euiaA5a+IFi+NjwjrhtuKTT2W/jttjG4bKWAyzg4pJSaLkKnX6AufktOo5jlXNYDK2
B8sDy8tmupw4xR3vmE+bUOJGG2xAivETwXInf9eyE52fueMu4E9eImcmeDlt+B65JgmJ4UdFx6qC
ldtf0oWV9VUONkxX6mVhWrAgfRob4LRcwoiTgiZZa3qn2x+uvkDXMIYGms3vg639IxJM2CCL2Cwr
jlkHUpRus6hxFS8mjzp21GxRYPmG2CFhcKhhK/tEW30GrGWVipM6lqbJIwtMyAm1ogjKYRlunwYS
zsE99SV9omEhrblde86F60ITxplZyiWwmLWwHklhQuoVTIkuH8L1WkGEKfIfLOnVmZh+f1kzcu0h
E/YerW+teGl5jT2DawK9wmYo87F/4mfQtuluV5u2b2YgnVldmPyldfGwAkulCuLzrQzmmrgxPjjl
bVzSJMRGFUULNd306DN6N86Kg9ZwKlRO0YK4ffjLq1P3smCi4ehBmd6ACmTKtsdXHhOvIYgV09mv
g7HqW/2IX69fYmiLdWiYRdyOFiMhEKeoI+EM/I5hD4EV7FUHxCqnj//y3gb714JrIzFLILSZ60FG
l9x50lM4c30mREI6ZM93qmw2Sb7WkndwoyavoBmKNm/nmoSkLGyPFK1zkdtB7qY5RkBvc4ikPSsp
C+1sOo+VbvBZ7DJVVKlTw14AW8W0+Oy0fj71FYBix3aLxqXUayZkcVfZUlsqU5x8oZZzHO6NjQjt
L5baHvmaUU0R3NaoZX2B+ZJdB89Ye1WG1FP/4NTQrWS2OsBXXwIonFOh/BnNhpMeWhwqQLi7RFrL
/lbPXMCPdIgzyADiN7D3PESjl/gl6i+bke230e47UTDR4MNgUxpcsn/eSW8HwokOnFXLu9WnHFbB
1f/ZOOuXi/qBN79TlythJzombJ1JYtrgVw9jEYGb1EugRB0E2zuwrrxjc8Q0qS7lgIhKE4c9gth5
es+gVcJqIufx6EbCRyCuEQ2KhCNm4SbgjOlGanEZJ9JhZUV8mfnHU67MgE+pGKaQQZxJ3XcsPhXv
mqifJQw216r5F+Mrw/CO5Iadc0eyCRWvw8VKE081eB8JnV4o7J9Wiv5EcHiSI43wVpCf2XkDHIAq
rMQC36Nb3zEyr3gmBpAtu7Dq4OnEfzFtL4tjUd6pH9Se5x3x0IwhaiFd6RVDsfyA06Jo/nqtGYRp
f96WheT6FTyWEh6nNpU/thXInCfNpVODP94vsvPdVV+pRMXKbDvAos7zVC1u6SVkteoB6/Ob29qk
1DT9Cm+o3GUM3647s6cEtvy3CpDwZyNCCMfXrjXC5T7qTxifSVs9zYAKAOklPhh682aJzJopE5+j
tyFpjeKo6S28YJdIjIGp6gWKuVB2LII9uQMr9emvWYl1XPOHORYZ+KMMFnxtOXkFa4ZzyPBjIx23
XaLvJxwshTpHuHA6Gp5PAEV1LMqcj+u2+DCt4ADFn4+cNV8xNikAP9N+NbRljAdg5DyBofT9l9UO
1+CT7ylUOCJ6Y5jKwgshzGdaLQ/bpeRXompFWa5vzfHc4fbTaGp9CWRpIaMptgCZMmU6YVESaO3M
6XchZ6A2ve5NYGMczlVK4h0MUV0V13J0QovCfCmJ0IqeWTHlHgHVkyRTO+0xh8algqOkEaJYw++O
hmJciYOlgpaPxXz4SPdNOo609IlpjR6HreOofOtwk05YiayxvXBYc3XjK80vUMSlI9bJmvGujzAS
vaobFxl8zORQ58FoTiijZ/DabK42FFwnsUIMmDGqYZ/MXxeX+vAYKeEkF8+opNIM9jSrW6OJjUeY
VyKQjJIXpR9giDNSCZsFf6VvZ1DrxhDd7PMnU1LdqGCajilyBiOIFJ3iygWyABe/cBdWt+CkfGU2
51ZIxv/V1PwcEZnRMFRirGJOayyKrsyadgiJzDvymGD+nznZA+YymNkk8eF43NeWg9ZFfvcTcDFY
bqBX3SnfDuzfMt+rKKPDQVJMyPOMWoDCctbk2jcXFKnVvnGQ4UvKtChNUB4MELcJC6GD5OCV9EhG
MyoT3I/GbJq46wWvbpX5BRId+2ILJELnHKjIeUSu+rdEsk2HD9ekVulnRBPfXFGxr2QA5V+89H2W
WVt1PYKIoe6E01XaxVzl0R7HrzI8uNv05IDmmHGQQaXfAobu9Il2Etlvihpn5JiUWR1d4f1sf1kS
0FvznZUpuxbYQkAwYxWsSBUE6jYWkw0tcAAse95UmFtN5AKSY93IPvFhqGUz9WXUQVXqRYt5Rmg5
TbF1BAATl4AaJRGnU4oBYBcyrsr8ZsVn46epVvqsUeyYjIj5q+CNCmzX74QB4cil2esMZ3P2tybA
eA8o+wSv8moTgUwhMY0EdU3C3ngiiRkeOLLZBZkOqB2QthFqua6ZCBjXaa433d44nuV36jim0ZLP
2ntYvIZK/9hqd7ECUHBxY0gtkRHntPvpJGr08nFAlhlqS/NW/kBmKENypkYxdE7wGF1EEy7xQNNn
rFtLioul2CExRbFli4AuGYPJ9RxfT6/LVZ1q4ZouO5nRSYdELa6F4KHJJ/VmCRQnhXquzL6ZFoUz
h5MLIWR61N8s0SQljrD274OARJg6S5ZTXDDjJB1WT5NlsKcOkSvYqAI+YPWSsbu8ZO/Va2Jfk9xH
/fVkQHVDM2PqR1w+hpcbmPOwfpgaGAeHvIQicvXCax3p/ndRwopbDVpW6LBD42ERAjm0xJ/lBEx1
wxAiL/V7MSGszahI6viV9ftJg2eEATcjf2xJi/rVUvrQjRF477XSownQOJ6PCJ4q1gnV/2dsluln
CJg7H9mRgMvcBasB2yL9T20il7mt/JBmKurfYsu31ScPXKaZqKpN26ro/+m7mnYT2n6CQAcCQPN/
tf1RqZCzAuSiFY1775YyJu7jcmg2IHxVCPcBEz+2uysadt0NvcuS7HzWwt0CrFE5JQnG9tkMrEm2
V3Uus33ghSn0uD3kSfCU7BPqv8WuzDxzwrTRtB9LiqHQvuw8QLed+AkBBtIyZsNvndx6RlZRpZm9
pDwupZVmAR1VqsymszD7yc/gh22tqKyg+yamz7r8p5G8BRMyR04K7I6VvRG05llVsej+XdjngAyk
uV8UabEgtH+wS6wjkUuphovWCvDz6b4bVNhxPtpP4AuqjlxbtFhtWBnyvZH2Up98We1BG3Up6oZk
3XIgf2qbUi1MrZlKmfWY8gzpQEhxQoxgRiFYHWAheAlwznH1yjbR+GSOb+3Toi+t6xrGj3Qmxvxs
zdcc/d+808xz9Add/X7CF/G6EFJrT2SPggCK/xfWhJ8gcJgy3UW8Pi/5TMVCL+PewCOzpnclJzze
R8QzG988mLUXhNo9PRrFm90Ff8sCZNmP5BnsxUAVX/1b2OKk6aYcjd0+8P919VJO2J+g9L7T4+tG
zf8477y24MEzSSulXRP0pmF0swrIE4WUmCqaOpMlHNsRCJNTOatJBkfJJ09K/h7dERs/lbgEVIR7
fsQDYKTuG3bTmfSEgXmoyvbix2xwjXZNf70qvHlpoIJ87rV5gNT+YxI5yo9bjUFvo0MoWRKzFjvF
VJvexJTgkTGiuKrF8TeH1Wycs4fNA8PVWhmKpYlGcuN5S4U0p7aK0B5FC2XBQ5BQxL/5XVJoCy+1
vkIrwVnGJbl1q3Ksf7LN47hB4AOIWYuUl4MZwV/LQBkizg02+y2eAztzftl7ONjLh/iZSnSeuQXX
ikmtc2FofnQnhzt7M83TovW69LtkIY7IlT/SBC89ySgV6Z1FNrsbShcA/LTVa2VgUz5ZDMi5hGRk
x3Q/9buBer6TefCWL2p9xcbBLEQba0X7NZq/FDVaSOZ6okRjl2Sjc4t/A3yU4gX/2hdm4jJBSv+b
5mrT5soMv0NTbXzYFNGe95oI+1/2VBrCo/3b14OqX/GGZRdJutykwii9w0Cj5GrZe0cWlN+m1Pi1
lLaZNffKYLILI03JjbZ6BR3OaH3Uy6gIc1c1fV/ySVbrmTP/9ue8tDrN8YHms3htwa+b4NcFBbg5
+KZwP69f8L3X6tTtuFF0gZbRsKIjIxm2usnwPAq2dpb/OORV+8VtFnl8e605z3S8YgAlA2tXwAsi
RLQ1aP5ubbt9wEWbbtyHf+hX5YdqZSl/OTI4vuArJjuAeCHVxu94X+JVgkmKj/K7MJdSz6BEc8ik
1DGNDSYBGrBAQhTw5Zf+Ukv/w3swtaiHhFIZwmj1JEjEvMuuT+rS2TQ7c17M8PNEPbIKlYfD3V+e
t3vFGSJ6NsH1u61RhDNxwoOXvZGraEs1irZwpeSN1pLyCVYDPFEf/e7IUxRKnSnThDAN9hq4nkIn
mw4o+0Pb5tXP562KlZgmFcb5vupDayoKllnZj2tkfvYhOXPy7zWh4gUmFH1DmmPZaUiaz6U8EUBz
evhdKWWhDID74bNDalpqwcazAgse0nmsbFpb/l6qJXvXNhQIP62K9kJ6dIux16DeFc4qz20au0/E
3CiSe7R95hjSyl66uc79kwEnyjgNw61SqfBm8SONxUp7XfoHZlpZX6sWYiAOx4MzfzRP48b9ClvI
CLdxSWek70SmtbMCzyF8LKONoVRZyM1ynFUy/suKJZbGPKxFVSjf/VNJeqEv1wNCPMbt7RUrybbC
N5Y+Sy7DoDUMFSOVc8tqY76Esgwwzz60XxVIGUNOrvN/1KQlNCLyMygc5PjAAcgS6T6rN9oe6FX8
Oi6+bGmaHy8wne0pJQlb0+fHMh5acBIbPmbbkuK5gD+aoPEd5Z32SAvsqXhCzkk7ltFUCfCb7mpJ
Mzw/Hzs7bw7qRu0yet5EYAnRrXvpXcd9+kYLCn6PEjxA2l8QOlXnBvqPzRlqEeX9vEFCzWIyowja
DugRUdjo+jilTGckCIYEGkJmZnLEyato+8wTOS4XCiY4ZGugyMHSB9A2QjLMRpIjhDGoJd78+YY7
DnOADak4UMqa/zQhHG5lc98lNhDDuiytMnteJB3L6QiHqjClggj8LbWtDkwhXuuiTFcT7ZJMI/2R
lsbLWpdDxdxNSdrjHp7Gjs96B0tvNqCk8efYukxyFZhLHJt1UWiVj52cFeu2VM65gYqpCucH9AHi
SQe7AwzGlq7H7TFlbSDjnKDPgVeURVBZ9tRJkbMYJqmUzM0OwHR2tf2BgcCPzjSRPWOo+yAxpP5+
0N/qBcb2v9BgxDaXOsAgYYsB+tSWd3cAONYZdaGIqFTz7w8lGYo7WWm4sf+BwynBWocYQqfkGmbJ
CKQ52ywA9EvbJk+wifIp8MMCMM3PqBLL8vnJ8zYi1bX3DuMdqf1j+aOYOWEznOD6at6WomrW0S8b
JpcNAu4nqLuNkpIOCGues3NzK+BPYcyyjp4fkSSZINv7kyvt0qQWs2vPQsMyt8B9zzXo1Mz0UaJC
s4SD6u1hUhyNssTpNEKOiJlMVgYjlH+P0xaYQK4/ng2Eso1wApC7oKtC7uMnvLUCn8KubJtkkm8B
r5A3AZDCDQnF4FA/yhrGLTaUrWrjezvoG2S7cp9X8HDZPXvADiX9WmBbdG8Y2K0W09wGxX3ZbHh9
Y5iPf9iifJ4cfPQELOTvYcX+MI6Z3gtOFCLZbjzxyEpvKN8ZtLR8fCMUNRJsbJ7ibX9JLHJ1QGKt
8yagevINqTKbJPb5QohIEUQGIWeoQ/9efDC9xOFhlTVJqts6XoOlSx7C63G0upg2yJIgm9LE2lCX
c90sHgEGfZYxQui0xvMc83O0WyhyEA/H/ITKxs0VdKLWe8gSgM9BDhJUPf6L1FVpirL3HP5G6EhC
BtrJ/4IAmw8yzrkW4DK4tZoUtcBCWhMgo94uqKXRM37yIgZaHPofAnzgKFkXdxdsec5eFsDDtjmZ
EXT8vuIgevmKPzB8GnkAduyW8ukMNulUFEidUVedI/q2O2i7x8DWAvIYBTWbDUoiz4inqN6Wk/fQ
rzvQKipVc4P8YPTe7D2xMesGFQrbkd+KsRqB0PxBhfwuki3c7OkiP74EWwpQbCTpHB7qZAX1VODK
CCXCNrpfx0AAB292hjMm1l8picKe0Y8FHp63js0Ii7bDpy6afJUJ8rJiaf9lQEaBtBUH3d/+/5Dx
lv7LF9TthRUQ6MgD9tEZr88/buWb4Kkq3Mbfvany0UU9Swa32GbR7jlFlAbVElAHvi/oQiTrTNqi
D1uPOiTQSdFhtwLOH0k5jazlIBlc3M87yvGxv1LODsxMpPBjawbUq8MhmnnSiiZf2TAVYpxYXFPp
DUTcoK2x6zvAV3irhaYu9um4Uzsp7Uei7aw7YGhKrVy+nRDBdDwAAWoMsNpdn40HmmmXuRr/7beV
LoZnMXtXZVSjNbY4CioXL6F5/WZTGSmA8ACfv7aX66XrucaH3AeVuPKjQL1ikPVnrFmwX65Thrjo
TbHm+Mpb+UdCmOxhif9Q4QNNPzgk3Tj/CY3Pp6fYwlixQQn1dtf3dh1bx5uJldgcMeY1pcDr070S
UiYm8dLzrFkMHgxy2E5W8H6IDxGHawIW4iwcxXCsvhXQ+78TGkDyCjxdc45u2viPwbkLXPquEQvm
go+YopzXJUduQ3RMpImftZkNhkewA8p4vs+7inkjrb15SrmjCRCaTL695SyAvYWf+ZLzLUj7rI8D
DhJgWdnJMkb0Z9aQSYIUV/+AwOa8ocIFvoiekwb5pdaITP8vob1/15rIs00zV5tMYhZQlUJXHUzW
7yQwAJe2rbnraBuw4wPvpZHaR5TFsXydLFzR4ExZMc4EVyoJQkkxtGTGRXtDtwuV0OCLs2N+h/ye
zppmM9jf5PpCwRpBsNOEbwOMO3V5RCNXc+2gSXZLCiG2MvBNpF51Ojhz3LR8PoVW//JsGqFH64ez
Gw1Sgq28fd6Atc6q3N5FQXu0algQo8JnswwGjfDy7Z1WvRtj56v6KvFIqY2UksqN1dd5InIfPuF5
A4lZDKwfTCAh7NLuPKZeqA1cVHKQrKlQW/cOsTVNCctTXYMTa74GgXWWbzmm/QsCaWyanyRAGGeI
MHLcwTxe+KUhjv28ng630SJpDh1YQ4IMPNCah6AVV4jccbraIOkVyFortcgI5h927nddqrdyNE+5
cyKrzFPfirjsaY9jtRMSAPo2FIc6maYRQYDdiNQuTZEq2MqF3ssJE/FjhJB2yGOVhhEsoTGHvtnC
CUbqzflPeu8GKVUU4Y0BCZWu5FLOjmLpFCwoqYsAe5TQ8gNs0WJHXITItgxT3LtIe5VwpAmqTLrz
nM66NAXvHYCpnTEM8JUqXBLftygUdSAv1eY3JeQCG1+20CsEQQhADZ4AfmaIryJ8YEU1Bh0YabK8
VSaobAlN8YFe/MGMB49Pwv+1CnYeFPlu3bY0p9C4NG+OqysUG5+wzmbkOhB+fyDMh5c0vjzJ0EXS
FK/1cez7hgGXFPaKwo/f7uBUWvDhHUvptH0AZflQ/ODVsjC9T9MaW3ZeSO+uaUvfHrc/02Z1s9mZ
EqwcRNdvIfgOsE0EmOmov06DuOOAXgT44xmLNgXho2wKF0C3kFSQSA7dw/u81Uj3KrSw9lhmKalm
jjDMljZOkKOI8c2msXSd1ByrQ/AUJfIJkzBD+NO7dZEpUywiqrDqtzD+/YazUGBtZDK6Cc9xmUUs
NuZRL7r4UF+jNdzvC0bDibf/fnzwbWCIqsUUoSu6XjTzj1Pk7unYPfIToU5djwleaS3tVxgqdIzS
FGOj5JeBLoZYjg9hbYD4G9T311EWl6bHRsT7FJOTWudc8XJgxN6Zi0KDPOAzE07wPc78hGrXD53g
1vRQiUNyBzXom2vKswr3zUqKgSdRmRcAhNME3qt/I0PSFO2yA+LrRU+nw1I0aua94NAP7eBmOAxH
gK4nswm3JdC2LBBgAC8/BuCqMHfryNLnSEhEFO2S2T1bYdmduz32+/UptOqH2IgHlydh9ph4PEIY
YJoQaxfUYOzhWAKrjeKNK0sHipWqSn/qd6nvbsYtw+raa466dzepbKbf6QiRmektIDgJRgd14BzA
KwK0POh6RH8v8bKTrKhbbh4+duYxIIdX9UHrXtcHvfgCamB1GodI4eIqYgL6GLslA2B03oIejQwK
ks5kmuaMmlM3y8m9PvWQncdn2QDafrFk2Cqd2PRgR9ekKpJy2wf+oNA/puvaRKdHEt0hxgqSBb5h
HD/EyqH/i3J+CiSnQk1UoJQzQx+RLV5EddLXoafpvUhuWiM3gybU4RwxQq8K8WY0sjxM73LMoFn0
CvTlg0E5Qp1Ga1ECyCCXRzQeMiXz9xPdQ2WLJJurzcI4Dizj0TnW9b3xAQYXt64AtXdkr8QZbwWS
TUy8BOGka6cHx3YDuqQ1ZDAKP4b4gRJm//WPzziZeAiuVkfFclspu9tq7ItNawmd6UI5o5kBbcQy
s2mXMdb8aMnj33mirfwvryhQQhyufOTdbcJtepeiXH1/hdkVhpYLX7n/E03U/LZPM9CpJVfNWhdj
uhCejo1nvTziy+ZM2FRwSFkj1YKLI1z/jFhiuQb+ZC/T2Kh/vh9vUwfivGLlxuVHoDxUKpge5xip
ObGo/JNakyGm6nMmcv8JNx+U1ecpTze3MpfVYBq793wmbxrYOw2TJzl1WQulQrzSW76rQi0dBBUa
CPSh1K++kdiVxWfU2lcbMuld23PsqsP+BbL93vL1qv4Y+mqFf/U8bmfTZFter+/I4O2gjpsw56KG
I0nGkS75SaidGpIsn1d3/CEEQHFesOoSewgdaoQcDIuWuoyOXgx2c8QZ8E5mjO/1B2RjwQyLacqV
aPMUb58kxqbQxeirOzUEI10f/6p/mE47KT1nra1VuPEhhwMFg5psS+y6CH9aFEIeva4P//MLRKF0
xvd5SadWZ5NQD+o9ONY4oZfwBapY8XuxvF/X2Gn1zmZmigZJrGGqvXbtvaSrGt80ybEWMlXLOERs
HS2eWf/JhO4JlBIe80iLTjr00sUSfLH6X+l3xKlS2BUMEWgUPXA1KaZnwmQxe32KXHeLEI3JFMr7
jXhP5CFmIPR+jFwgz+7t1nK4LUnfCyPJJ4N5apoZBQtPFf+m7wxA5dnmXWZQ+8t/8lCrCVNgPVyF
CBPyb/y/yK302AhoJ09FOVc8B0sztgj1t7x0FMu7kGyNho02R6yS8KhuQ1vLvVbAbfLT0BkoGzto
C5TPNW9LjyuWb0+Ka3pcU4pbGTThUWdnMpP5QvOC+LbqCfi/9GM17iwQPZqgYlZu11/vJ+h73/8P
GzLeTpUOTzjulxwc8mCMVTgZQgxmTB4rIsozV/KYZq/h4hiVA1NdMONwBy693SkCyF//y5iPogQv
V6rrjRX24H4rDIPFHGKiXdf3AH0rmGMzJ9kQH5+h+R6DYgmH+2lseY/LWNmWMt8R9wk3pCfAs1fw
BY98wKdoyJvpGCSGOdJBuh84EbuDbfK7X8GmSxR6LGel7SvLehAUCsxFdChjrxAz8iQCCNnFw0PO
rekrtGqFSUsLHBVwJNMT9TLKJqCXivA9IfPrFNyO9PB8Wrd7ye+HIZEJK1aBifPX5esINR+F9I1l
0t2KLSFKo0JaJN2VuLoXBlXyd6JqAj08CHvjSO7LrUmma6qHAgfnhd/mqWqM5LDPx7cNZe/23iuk
vU8NBcN3d7b2c9WCf318NDG/SHVz6rjMda1PzUDXkez2Wv/dPrHEpQIqdKqIB7++wSkSqluMqVZd
FmDFdvbkWDyIbgReOE7T5eA+cbd3bPnNpZymRiSrXaR7
`protect end_protected
